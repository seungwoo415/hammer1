* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : DigitalLDOLogic                              *
* Netlisted  : Wed Jan 29 01:01:39 2025                     *
* Pegasus Version: 22.14-s007 Tue Jan 31 16:35:56 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 1 MP(pfet_01v8_hvt) hvtpfet_01v8_rec pSourceDrain(D) hvtpfet(G) pSourceDrain(s) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__dlygate4sd2_1                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__dlygate4sd2_1 1 2 3 4 5 6
** N=9 EP=6 FDC=8
M0 3 4 7 5 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=505 $Y=235 $dt=0
M1 8 7 3 5 nfet_01v8 L=1.8e-07 W=4.2e-07 $X=925 $Y=235 $dt=0
M2 3 8 9 5 nfet_01v8 L=1.8e-07 W=4.2e-07 $X=1895 $Y=235 $dt=0
M3 2 9 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2400 $Y=235 $dt=0
M4 1 4 7 6 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=505 $Y=2065 $dt=1
M5 8 7 1 6 pfet_01v8_hvt L=1.8e-07 W=4.2e-07 $X=925 $Y=2065 $dt=1
M6 1 8 9 6 pfet_01v8_hvt L=1.8e-07 W=4.2e-07 $X=1895 $Y=2065 $dt=1
M7 2 9 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2400 $Y=1485 $dt=1
.ends sky130_fd_sc_hd__dlygate4sd2_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__clkbuf_2                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__clkbuf_2 1 2 3 4 5 6
** N=7 EP=6 FDC=6
M0 3 4 7 5 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=400 $Y=235 $dt=0
M1 2 7 3 5 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=875 $Y=235 $dt=0
M2 3 7 2 5 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1295 $Y=235 $dt=0
M3 1 4 7 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=400 $Y=1485 $dt=1
M4 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=875 $Y=1485 $dt=1
M5 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1295 $Y=1485 $dt=1
.ends sky130_fd_sc_hd__clkbuf_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__clkbuf_1                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__clkbuf_1 1 2 3 4 5 6
** N=7 EP=6 FDC=4
M0 3 7 1 5 nfet_01v8 L=1.5e-07 W=5.2e-07 $X=395 $Y=235 $dt=0
M1 7 4 3 5 nfet_01v8 L=1.5e-07 W=5.2e-07 $X=835 $Y=235 $dt=0
M2 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=7.9e-07 $X=395 $Y=1695 $dt=1
M3 7 4 2 6 pfet_01v8_hvt L=1.5e-07 W=7.9e-07 $X=835 $Y=1695 $dt=1
.ends sky130_fd_sc_hd__clkbuf_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__buf_8                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__buf_8 1 2 3 4 5 6
** N=7 EP=6 FDC=22
M0 3 4 7 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=395 $Y=235 $dt=0
M1 7 4 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=815 $Y=235 $dt=0
M2 3 4 7 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1235 $Y=235 $dt=0
M3 2 7 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1655 $Y=235 $dt=0
M4 3 7 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2075 $Y=235 $dt=0
M5 2 7 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2495 $Y=235 $dt=0
M6 3 7 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2915 $Y=235 $dt=0
M7 2 7 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=3335 $Y=235 $dt=0
M8 3 7 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=3755 $Y=235 $dt=0
M9 2 7 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=4175 $Y=235 $dt=0
M10 3 7 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=4595 $Y=235 $dt=0
M11 1 4 7 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=395 $Y=1485 $dt=1
M12 7 4 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=815 $Y=1485 $dt=1
M13 1 4 7 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1235 $Y=1485 $dt=1
M14 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1655 $Y=1485 $dt=1
M15 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2075 $Y=1485 $dt=1
M16 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2495 $Y=1485 $dt=1
M17 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2915 $Y=1485 $dt=1
M18 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=3335 $Y=1485 $dt=1
M19 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=3755 $Y=1485 $dt=1
M20 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=4175 $Y=1485 $dt=1
M21 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=4595 $Y=1485 $dt=1
.ends sky130_fd_sc_hd__buf_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__dfxtp_1                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__dfxtp_1 1 2 3 4 5 6 7
** N=22 EP=7 FDC=24
M0 3 4 9 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=395 $Y=235 $dt=0
M1 8 9 3 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=815 $Y=235 $dt=0
M2 10 5 3 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1755 $Y=235 $dt=0
M3 11 9 10 6 nfet_01v8 L=1.5e-07 W=3.6e-07 $X=2315 $Y=235 $dt=0
M4 17 8 11 6 nfet_01v8 L=1.5e-07 W=3.6e-07 $X=2810 $Y=235 $dt=0
M5 3 12 17 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=3305 $Y=235 $dt=0
M6 12 11 3 6 nfet_01v8 L=1.5e-07 W=6.4e-07 $X=3900 $Y=235 $dt=0
M7 13 8 12 6 nfet_01v8 L=1.5e-07 W=3.6e-07 $X=4405 $Y=235 $dt=0
M8 18 9 13 6 nfet_01v8 L=1.5e-07 W=3.6e-07 $X=4935 $Y=235 $dt=0
M9 3 14 18 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=5410 $Y=235 $dt=0
M10 3 13 14 6 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=6355 $Y=235 $dt=0
M11 2 14 3 6 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=6775 $Y=235 $dt=0
M12 1 4 9 7 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=395 $Y=1815 $dt=1
M13 8 9 1 7 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=815 $Y=1815 $dt=1
M14 10 5 1 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=1755 $Y=2065 $dt=1
M15 11 8 10 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=2180 $Y=2065 $dt=1
M16 15 9 11 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=2655 $Y=2065 $dt=1
M17 1 12 15 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=3170 $Y=2065 $dt=1
M18 12 11 1 7 pfet_01v8_hvt L=1.5e-07 W=7.5e-07 $X=3830 $Y=1735 $dt=1
M19 13 9 12 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=4305 $Y=2065 $dt=1
M20 16 8 13 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=4725 $Y=2065 $dt=1
M21 1 14 16 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=5295 $Y=2065 $dt=1
M22 1 13 14 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=6345 $Y=1485 $dt=1
M23 2 14 1 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=6765 $Y=1485 $dt=1
.ends sky130_fd_sc_hd__dfxtp_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__a221o_1                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__a221o_1 1 2 3 4 5 6 7 8 9 10
** N=17 EP=10 FDC=12
M0 3 4 13 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=395 $Y=235 $dt=0
M1 14 5 3 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=875 $Y=235 $dt=0
M2 13 6 14 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1235 $Y=235 $dt=0
M3 15 7 13 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2175 $Y=235 $dt=0
M4 3 8 15 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2655 $Y=235 $dt=0
M5 1 13 3 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=3120 $Y=235 $dt=0
M6 11 4 13 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=395 $Y=1485 $dt=1
M7 12 5 11 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=815 $Y=1485 $dt=1
M8 11 6 12 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1235 $Y=1485 $dt=1
M9 12 7 2 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2175 $Y=1485 $dt=1
M10 2 8 12 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2655 $Y=1485 $dt=1
M11 1 13 2 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=3120 $Y=1485 $dt=1
.ends sky130_fd_sc_hd__a221o_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__a21o_1                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__a21o_1 1 2 3 4 5 6 7 8
** N=12 EP=8 FDC=8
M0 3 9 1 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=405 $Y=235 $dt=0
M1 9 4 3 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1345 $Y=235 $dt=0
M2 11 5 9 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1770 $Y=235 $dt=0
M3 3 6 11 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2200 $Y=235 $dt=0
M4 2 9 1 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=405 $Y=1485 $dt=1
M5 10 4 9 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1345 $Y=1485 $dt=1
M6 2 5 10 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1770 $Y=1485 $dt=1
M7 10 6 2 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2200 $Y=1485 $dt=1
.ends sky130_fd_sc_hd__a21o_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__or3_1                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__or3_1 1 2 3 4 5 6 7 8
** N=13 EP=8 FDC=8
M0 3 4 9 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=405 $Y=265 $dt=0
M1 9 5 3 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=825 $Y=265 $dt=0
M2 3 6 9 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1245 $Y=265 $dt=0
M3 2 9 3 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1735 $Y=235 $dt=0
M4 10 4 9 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=405 $Y=1485 $dt=1
M5 11 5 10 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=765 $Y=1485 $dt=1
M6 1 6 11 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=1245 $Y=1485 $dt=1
M7 2 9 1 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1735 $Y=1485 $dt=1
.ends sky130_fd_sc_hd__or3_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__inv_2                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__inv_2 1 2 3 4 5 6
** N=6 EP=6 FDC=4
M0 2 4 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=405 $Y=235 $dt=0
M1 3 4 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=825 $Y=235 $dt=0
M2 2 4 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=405 $Y=1485 $dt=1
M3 1 4 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=825 $Y=1485 $dt=1
.ends sky130_fd_sc_hd__inv_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__tap_1                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__tap_1 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__tap_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__tapvpwrvgnd_1                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 1 2
** N=2 EP=2 FDC=0
.ends sky130_fd_sc_hd__tapvpwrvgnd_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_6                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_6 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=1.97e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=1.97e-06 W=8.7e-07 $X=395 $Y=1615 $dt=1
.ends sky130_fd_sc_hd__decap_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_3                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_3 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=5.9e-07 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=5.9e-07 W=8.7e-07 $X=395 $Y=1615 $dt=1
.ends sky130_fd_sc_hd__decap_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_12                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_12 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=4.73e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=4.73e-06 W=8.7e-07 $X=395 $Y=1615 $dt=1
.ends sky130_fd_sc_hd__decap_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_4                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_4 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=1.05e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=1.05e-06 W=8.7e-07 $X=395 $Y=1615 $dt=1
.ends sky130_fd_sc_hd__decap_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_8                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_8 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=2.89e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=2.89e-06 W=8.7e-07 $X=395 $Y=1615 $dt=1
.ends sky130_fd_sc_hd__decap_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__fill_1                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__fill_1 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__fill_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__fill_2                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__fill_2 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__fill_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_PR                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_PR 1
** N=1 EP=1 FDC=0
.ends L1M1_PR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_PR_M                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_PR_M 1
** N=1 EP=1 FDC=0
.ends M1M2_PR_M

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_PR                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_PR 1
** N=1 EP=1 FDC=0
.ends M1M2_PR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2M3_PR                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2M3_PR 1
** N=1 EP=1 FDC=0
.ends M2M3_PR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3M4_PR                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3M4_PR 1
** N=1 EP=1 FDC=0
.ends M3M4_PR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA0                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA0 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA1                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA1 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA2                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA2 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA3                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA3 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA4                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA4 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y1 1 2
** N=2 EP=2 FDC=0
X0 1 DigitalLDOLogic_VIA3 $T=710 1000 0 0 $X=0 $Y=0
X1 1 DigitalLDOLogic_VIA3 $T=6230 1000 0 0 $X=5520 $Y=0
X2 1 DigitalLDOLogic_VIA3 $T=11750 1000 0 0 $X=11040 $Y=0
X3 1 DigitalLDOLogic_VIA3 $T=17270 1000 0 0 $X=16560 $Y=0
X4 1 DigitalLDOLogic_VIA3 $T=22790 1000 0 0 $X=22080 $Y=0
X5 1 DigitalLDOLogic_VIA3 $T=28310 1000 0 0 $X=27600 $Y=0
X6 1 DigitalLDOLogic_VIA3 $T=33830 1000 0 0 $X=33120 $Y=0
X7 1 DigitalLDOLogic_VIA3 $T=39350 1000 0 0 $X=38640 $Y=0
.ends MASCO__Y1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B19                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B19 1 2
** N=2 EP=2 FDC=4
X0 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=190 2960 1 0 $X=0 $Y=0
X1 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=190 2960 0 0 $X=0 $Y=2720
X2 1 2 2 1 sky130_fd_sc_hd__decap_12 $T=650 2960 1 0 $X=460 $Y=0
X3 1 2 2 1 sky130_fd_sc_hd__decap_12 $T=650 2960 0 0 $X=460 $Y=2720
.ends MASCO__B19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B22                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B22 1 2
** N=2 EP=2 FDC=8
X0 1 2 2 1 sky130_fd_sc_hd__decap_3 $T=2030 2960 1 0 $X=1840 $Y=0
X1 1 2 2 1 sky130_fd_sc_hd__decap_3 $T=2030 2960 0 0 $X=1840 $Y=2720
X2 1 2 2 1 sky130_fd_sc_hd__decap_4 $T=190 2960 1 0 $X=0 $Y=0
X3 1 2 2 1 sky130_fd_sc_hd__decap_4 $T=190 2960 0 0 $X=0 $Y=2720
.ends MASCO__B22

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B26                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B26 1 2
** N=2 EP=2 FDC=4
X0 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=1570 2960 1 0 $X=1380 $Y=0
X1 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=1570 2960 0 0 $X=1380 $Y=2720
X2 1 2 2 1 sky130_fd_sc_hd__decap_3 $T=190 2960 1 0 $X=0 $Y=0
X3 1 2 2 1 sky130_fd_sc_hd__decap_3 $T=190 2960 0 0 $X=0 $Y=2720
.ends MASCO__B26

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic 52 26 66 40 1 14 54 28 16 42
+ 3 68 56 30 44 18 70 58 32 6
+ 72 46 20 60 34 8 22 74 48 36
+ 62 10 50 76 24 38 64
** N=181 EP=37 FDC=3456
X0 1 2 3 4 3 1 sky130_fd_sc_hd__dlygate4sd2_1 $T=162260 18160 0 0 $X=162070 $Y=17920
X1 1 5 3 6 3 1 sky130_fd_sc_hd__clkbuf_2 $T=171460 23600 1 0 $X=171270 $Y=20640
X2 1 7 3 8 3 1 sky130_fd_sc_hd__clkbuf_2 $T=172840 18160 0 0 $X=172650 $Y=17920
X3 9 1 3 10 3 1 sky130_fd_sc_hd__clkbuf_1 $T=60140 23600 1 0 $X=59950 $Y=20640
X4 11 1 3 10 3 1 sky130_fd_sc_hd__clkbuf_1 $T=80840 23600 0 180 $X=79270 $Y=20640
X5 12 1 3 10 3 1 sky130_fd_sc_hd__clkbuf_1 $T=134660 23600 0 180 $X=133090 $Y=20640
X6 13 1 3 10 3 1 sky130_fd_sc_hd__clkbuf_1 $T=171460 23600 0 180 $X=169890 $Y=20640
X7 1 14 3 15 3 1 sky130_fd_sc_hd__buf_8 $T=19200 12720 0 0 $X=19010 $Y=12480
X8 1 16 3 17 3 1 sky130_fd_sc_hd__buf_8 $T=19200 18160 1 0 $X=19010 $Y=15200
X9 1 18 3 19 3 1 sky130_fd_sc_hd__buf_8 $T=21040 23600 0 0 $X=20850 $Y=23360
X10 1 20 3 21 3 1 sky130_fd_sc_hd__buf_8 $T=29780 12720 1 0 $X=29590 $Y=9760
X11 1 22 3 23 3 1 sky130_fd_sc_hd__buf_8 $T=29780 18160 1 0 $X=29590 $Y=15200
X12 1 24 3 25 3 1 sky130_fd_sc_hd__buf_8 $T=38060 12720 1 180 $X=32350 $Y=12480
X13 1 26 3 27 3 1 sky130_fd_sc_hd__buf_8 $T=40820 29040 0 180 $X=35110 $Y=26080
X14 1 28 3 29 3 1 sky130_fd_sc_hd__buf_8 $T=41280 18160 0 180 $X=35570 $Y=15200
X15 1 30 3 31 3 1 sky130_fd_sc_hd__buf_8 $T=47720 12720 1 0 $X=47530 $Y=9760
X16 1 32 3 33 3 1 sky130_fd_sc_hd__buf_8 $T=62440 12720 1 0 $X=62250 $Y=9760
X17 1 34 3 35 3 1 sky130_fd_sc_hd__buf_8 $T=65660 12720 0 0 $X=65470 $Y=12480
X18 1 36 3 37 3 1 sky130_fd_sc_hd__buf_8 $T=65660 23600 0 0 $X=65470 $Y=23360
X19 1 38 3 39 3 1 sky130_fd_sc_hd__buf_8 $T=73940 12720 1 0 $X=73750 $Y=9760
X20 1 40 3 41 3 1 sky130_fd_sc_hd__buf_8 $T=73940 18160 1 0 $X=73750 $Y=15200
X21 1 42 3 43 3 1 sky130_fd_sc_hd__buf_8 $T=82680 12720 1 0 $X=82490 $Y=9760
X22 1 44 3 45 3 1 sky130_fd_sc_hd__buf_8 $T=91420 12720 1 0 $X=91230 $Y=9760
X23 1 46 3 47 3 1 sky130_fd_sc_hd__buf_8 $T=97400 12720 1 0 $X=97210 $Y=9760
X24 1 48 3 49 3 1 sky130_fd_sc_hd__buf_8 $T=103380 12720 0 0 $X=103190 $Y=12480
X25 1 50 3 51 3 1 sky130_fd_sc_hd__buf_8 $T=103380 18160 1 0 $X=103190 $Y=15200
X26 1 52 3 53 3 1 sky130_fd_sc_hd__buf_8 $T=114880 18160 1 180 $X=109170 $Y=17920
X27 1 54 3 55 3 1 sky130_fd_sc_hd__buf_8 $T=115800 12720 1 180 $X=110090 $Y=12480
X28 1 56 3 57 3 1 sky130_fd_sc_hd__buf_8 $T=123620 12720 0 180 $X=117910 $Y=9760
X29 1 58 3 59 3 1 sky130_fd_sc_hd__buf_8 $T=123620 18160 0 180 $X=117910 $Y=15200
X30 1 60 3 61 3 1 sky130_fd_sc_hd__buf_8 $T=132820 12720 0 0 $X=132630 $Y=12480
X31 1 62 3 63 3 1 sky130_fd_sc_hd__buf_8 $T=138340 12720 1 0 $X=138150 $Y=9760
X32 1 64 3 65 3 1 sky130_fd_sc_hd__buf_8 $T=144780 12720 1 180 $X=139070 $Y=12480
X33 1 66 3 67 3 1 sky130_fd_sc_hd__buf_8 $T=153060 23600 1 180 $X=147350 $Y=23360
X34 1 68 3 69 3 1 sky130_fd_sc_hd__buf_8 $T=148460 12720 1 0 $X=148270 $Y=9760
X35 1 70 3 71 3 1 sky130_fd_sc_hd__buf_8 $T=162260 18160 1 0 $X=162070 $Y=15200
X36 1 72 3 73 3 1 sky130_fd_sc_hd__buf_8 $T=163180 12720 1 0 $X=162990 $Y=9760
X37 1 74 3 75 3 1 sky130_fd_sc_hd__buf_8 $T=176980 18160 1 0 $X=176790 $Y=15200
X38 1 76 3 77 3 1 sky130_fd_sc_hd__buf_8 $T=180200 23600 0 0 $X=180010 $Y=23360
X39 1 23 3 9 78 3 1 sky130_fd_sc_hd__dfxtp_1 $T=48180 34480 0 0 $X=47990 $Y=34240
X40 1 27 3 9 79 3 1 sky130_fd_sc_hd__dfxtp_1 $T=48640 34480 1 0 $X=48450 $Y=31520
X41 1 21 3 9 80 3 1 sky130_fd_sc_hd__dfxtp_1 $T=49560 18160 0 0 $X=49370 $Y=17920
X42 1 19 3 9 81 3 1 sky130_fd_sc_hd__dfxtp_1 $T=49560 23600 0 0 $X=49370 $Y=23360
X43 1 15 3 9 82 3 1 sky130_fd_sc_hd__dfxtp_1 $T=50020 18160 1 0 $X=49830 $Y=15200
X44 1 33 3 11 83 3 1 sky130_fd_sc_hd__dfxtp_1 $T=51400 23600 1 0 $X=51210 $Y=20640
X45 1 31 3 9 84 3 1 sky130_fd_sc_hd__dfxtp_1 $T=59220 18160 1 0 $X=59030 $Y=15200
X46 1 25 3 9 85 3 1 sky130_fd_sc_hd__dfxtp_1 $T=59220 18160 0 0 $X=59030 $Y=17920
X47 1 37 3 9 86 3 1 sky130_fd_sc_hd__dfxtp_1 $T=59220 29040 1 0 $X=59030 $Y=26080
X48 1 29 3 9 87 3 1 sky130_fd_sc_hd__dfxtp_1 $T=59220 29040 0 0 $X=59030 $Y=28800
X49 1 39 3 11 88 3 1 sky130_fd_sc_hd__dfxtp_1 $T=66120 23600 1 0 $X=65930 $Y=20640
X50 1 41 3 11 89 3 1 sky130_fd_sc_hd__dfxtp_1 $T=75320 18160 0 0 $X=75130 $Y=17920
X51 1 35 3 11 90 3 1 sky130_fd_sc_hd__dfxtp_1 $T=77160 23600 0 0 $X=76970 $Y=23360
X52 1 45 3 11 91 3 1 sky130_fd_sc_hd__dfxtp_1 $T=80840 23600 1 0 $X=80650 $Y=20640
X53 1 47 3 11 92 3 1 sky130_fd_sc_hd__dfxtp_1 $T=90960 23600 0 0 $X=90770 $Y=23360
X54 1 43 3 11 93 3 1 sky130_fd_sc_hd__dfxtp_1 $T=93720 18160 0 0 $X=93530 $Y=17920
X55 1 51 3 11 94 3 1 sky130_fd_sc_hd__dfxtp_1 $T=95560 23600 1 0 $X=95370 $Y=20640
X56 1 53 3 12 95 3 1 sky130_fd_sc_hd__dfxtp_1 $T=110280 23600 1 0 $X=110090 $Y=20640
X57 1 49 3 12 96 3 1 sky130_fd_sc_hd__dfxtp_1 $T=118100 18160 0 0 $X=117910 $Y=17920
X58 1 17 3 12 97 3 1 sky130_fd_sc_hd__dfxtp_1 $T=118100 23600 0 0 $X=117910 $Y=23360
X59 1 59 3 12 98 3 1 sky130_fd_sc_hd__dfxtp_1 $T=124540 23600 1 0 $X=124350 $Y=20640
X60 1 77 3 12 99 3 1 sky130_fd_sc_hd__dfxtp_1 $T=124540 29040 1 0 $X=124350 $Y=26080
X61 1 55 3 12 100 3 1 sky130_fd_sc_hd__dfxtp_1 $T=132820 18160 0 0 $X=132630 $Y=17920
X62 1 63 3 12 101 3 1 sky130_fd_sc_hd__dfxtp_1 $T=134660 23600 1 0 $X=134470 $Y=20640
X63 1 67 3 12 102 3 1 sky130_fd_sc_hd__dfxtp_1 $T=135120 29040 1 0 $X=134930 $Y=26080
X64 1 61 3 13 103 3 1 sky130_fd_sc_hd__dfxtp_1 $T=153060 18160 0 0 $X=152870 $Y=17920
X65 1 57 3 13 104 3 1 sky130_fd_sc_hd__dfxtp_1 $T=153520 18160 1 0 $X=153330 $Y=15200
X66 1 71 3 13 105 3 1 sky130_fd_sc_hd__dfxtp_1 $T=153520 23600 1 0 $X=153330 $Y=20640
X67 1 75 3 13 106 3 1 sky130_fd_sc_hd__dfxtp_1 $T=162260 23600 1 0 $X=162070 $Y=20640
X68 1 69 3 13 2 3 1 sky130_fd_sc_hd__dfxtp_1 $T=165480 18160 0 0 $X=165290 $Y=17920
X69 1 65 3 13 107 3 1 sky130_fd_sc_hd__dfxtp_1 $T=169160 18160 1 0 $X=168970 $Y=15200
X70 1 73 3 13 108 3 1 sky130_fd_sc_hd__dfxtp_1 $T=176980 23600 1 0 $X=176790 $Y=20640
X71 80 1 3 7 5 15 25 109 3 1 sky130_fd_sc_hd__a221o_1 $T=44500 18160 1 0 $X=44310 $Y=15200
X72 81 1 3 7 5 17 23 109 3 1 sky130_fd_sc_hd__a221o_1 $T=45880 23600 1 0 $X=45690 $Y=20640
X73 78 1 3 7 5 19 27 109 3 1 sky130_fd_sc_hd__a221o_1 $T=45880 29040 1 0 $X=45690 $Y=26080
X74 79 1 3 7 5 23 29 109 3 1 sky130_fd_sc_hd__a221o_1 $T=45880 29040 0 0 $X=45690 $Y=28800
X75 85 1 3 7 5 21 31 109 3 1 sky130_fd_sc_hd__a221o_1 $T=50480 12720 0 0 $X=50290 $Y=12480
X76 84 1 3 7 5 25 33 109 3 1 sky130_fd_sc_hd__a221o_1 $T=64280 12720 1 180 $X=60410 $Y=12480
X77 86 1 3 7 5 29 35 109 3 1 sky130_fd_sc_hd__a221o_1 $T=72100 18160 0 180 $X=68230 $Y=15200
X78 83 1 3 7 5 31 41 109 3 1 sky130_fd_sc_hd__a221o_1 $T=72100 18160 1 180 $X=68230 $Y=17920
X79 87 1 3 7 5 27 37 109 3 1 sky130_fd_sc_hd__a221o_1 $T=72100 29040 0 180 $X=68230 $Y=26080
X80 90 1 3 7 5 37 39 109 3 1 sky130_fd_sc_hd__a221o_1 $T=73940 29040 0 0 $X=73750 $Y=28800
X81 91 1 3 7 5 39 47 109 3 1 sky130_fd_sc_hd__a221o_1 $T=80380 29040 0 0 $X=80190 $Y=28800
X82 89 1 3 7 5 33 43 109 3 1 sky130_fd_sc_hd__a221o_1 $T=84980 18160 0 180 $X=81110 $Y=15200
X83 88 1 3 7 5 35 45 109 3 1 sky130_fd_sc_hd__a221o_1 $T=82680 18160 0 0 $X=82490 $Y=17920
X84 92 1 3 7 5 45 49 109 3 1 sky130_fd_sc_hd__a221o_1 $T=92800 12720 0 0 $X=92610 $Y=12480
X85 94 1 3 7 5 43 53 109 3 1 sky130_fd_sc_hd__a221o_1 $T=93720 29040 0 0 $X=93530 $Y=28800
X86 93 1 3 7 5 41 51 109 3 1 sky130_fd_sc_hd__a221o_1 $T=98320 18160 0 180 $X=94450 $Y=15200
X87 95 1 3 7 5 51 59 109 3 1 sky130_fd_sc_hd__a221o_1 $T=111200 18160 1 0 $X=111010 $Y=15200
X88 97 1 3 7 5 77 19 109 3 1 sky130_fd_sc_hd__a221o_1 $T=112580 23600 0 0 $X=112390 $Y=23360
X89 96 1 3 7 5 47 55 109 3 1 sky130_fd_sc_hd__a221o_1 $T=118100 12720 0 0 $X=117910 $Y=12480
X90 99 1 3 7 5 75 17 109 3 1 sky130_fd_sc_hd__a221o_1 $T=119480 29040 1 0 $X=119290 $Y=26080
X91 98 1 3 7 5 53 63 109 3 1 sky130_fd_sc_hd__a221o_1 $T=119480 29040 0 0 $X=119290 $Y=28800
X92 100 1 3 7 5 49 57 109 3 1 sky130_fd_sc_hd__a221o_1 $T=125460 18160 1 0 $X=125270 $Y=15200
X93 104 1 3 7 5 55 61 109 3 1 sky130_fd_sc_hd__a221o_1 $T=134660 18160 1 0 $X=134470 $Y=15200
X94 101 1 3 7 5 59 67 109 3 1 sky130_fd_sc_hd__a221o_1 $T=141560 23600 1 180 $X=137690 $Y=23360
X95 102 1 3 7 5 63 71 109 3 1 sky130_fd_sc_hd__a221o_1 $T=141560 29040 1 180 $X=137690 $Y=28800
X96 103 1 3 7 5 57 65 109 3 1 sky130_fd_sc_hd__a221o_1 $T=142480 18160 1 0 $X=142290 $Y=15200
X97 107 1 3 7 5 61 69 109 3 1 sky130_fd_sc_hd__a221o_1 $T=142480 18160 0 0 $X=142290 $Y=17920
X98 105 1 3 7 5 67 75 109 3 1 sky130_fd_sc_hd__a221o_1 $T=158580 23600 1 180 $X=154710 $Y=23360
X99 106 1 3 7 5 71 77 109 3 1 sky130_fd_sc_hd__a221o_1 $T=156740 29040 1 0 $X=156550 $Y=26080
X100 4 1 3 8 6 65 73 109 3 1 sky130_fd_sc_hd__a221o_1 $T=171460 12720 1 180 $X=167590 $Y=12480
X101 108 1 3 7 69 5 3 1 sky130_fd_sc_hd__a21o_1 $T=169160 23600 0 0 $X=168970 $Y=23360
X102 1 82 3 21 7 5 3 1 sky130_fd_sc_hd__or3_1 $T=45420 12720 0 0 $X=45230 $Y=12480
X103 1 109 3 6 3 1 sky130_fd_sc_hd__inv_2 $T=120400 34480 0 180 $X=118830 $Y=31520
X104 110 111 1 3 sky130_fd_sc_hd__tap_1 $T=10000 12720 1 0 $X=9810 $Y=9760
X105 112 113 1 3 sky130_fd_sc_hd__tap_1 $T=10000 12720 0 0 $X=9810 $Y=12480
X106 114 115 1 3 sky130_fd_sc_hd__tap_1 $T=10000 18160 1 0 $X=9810 $Y=15200
X107 116 117 1 3 sky130_fd_sc_hd__tap_1 $T=10000 18160 0 0 $X=9810 $Y=17920
X108 118 119 1 3 sky130_fd_sc_hd__tap_1 $T=10000 23600 1 0 $X=9810 $Y=20640
X109 120 121 1 3 sky130_fd_sc_hd__tap_1 $T=10000 23600 0 0 $X=9810 $Y=23360
X110 122 123 1 3 sky130_fd_sc_hd__tap_1 $T=10000 29040 1 0 $X=9810 $Y=26080
X111 124 125 1 3 sky130_fd_sc_hd__tap_1 $T=10000 29040 0 0 $X=9810 $Y=28800
X112 126 127 1 3 sky130_fd_sc_hd__tap_1 $T=10000 34480 1 0 $X=9810 $Y=31520
X113 128 129 1 3 sky130_fd_sc_hd__tap_1 $T=10000 34480 0 0 $X=9810 $Y=34240
X114 130 131 1 3 sky130_fd_sc_hd__tap_1 $T=10000 39920 1 0 $X=9810 $Y=36960
X115 132 133 1 3 sky130_fd_sc_hd__tap_1 $T=10000 39920 0 0 $X=9810 $Y=39680
X116 134 135 1 3 sky130_fd_sc_hd__tap_1 $T=10000 45360 1 0 $X=9810 $Y=42400
X117 136 137 1 3 sky130_fd_sc_hd__tap_1 $T=10000 45360 0 0 $X=9810 $Y=45120
X118 138 139 1 3 sky130_fd_sc_hd__tap_1 $T=10000 50800 1 0 $X=9810 $Y=47840
X119 140 141 1 3 sky130_fd_sc_hd__tap_1 $T=10000 50800 0 0 $X=9810 $Y=50560
X120 142 143 1 3 sky130_fd_sc_hd__tap_1 $T=10000 56240 1 0 $X=9810 $Y=53280
X121 144 145 1 3 sky130_fd_sc_hd__tap_1 $T=10000 56240 0 0 $X=9810 $Y=56000
X122 146 147 1 3 sky130_fd_sc_hd__tap_1 $T=189860 12720 0 180 $X=189210 $Y=9760
X123 148 149 1 3 sky130_fd_sc_hd__tap_1 $T=189860 12720 1 180 $X=189210 $Y=12480
X124 150 151 1 3 sky130_fd_sc_hd__tap_1 $T=189860 18160 0 180 $X=189210 $Y=15200
X125 152 153 1 3 sky130_fd_sc_hd__tap_1 $T=189860 18160 1 180 $X=189210 $Y=17920
X126 154 155 1 3 sky130_fd_sc_hd__tap_1 $T=189860 23600 0 180 $X=189210 $Y=20640
X127 156 157 1 3 sky130_fd_sc_hd__tap_1 $T=189860 23600 1 180 $X=189210 $Y=23360
X128 158 159 1 3 sky130_fd_sc_hd__tap_1 $T=189860 29040 0 180 $X=189210 $Y=26080
X129 160 161 1 3 sky130_fd_sc_hd__tap_1 $T=189860 29040 1 180 $X=189210 $Y=28800
X130 162 163 1 3 sky130_fd_sc_hd__tap_1 $T=189860 34480 0 180 $X=189210 $Y=31520
X131 164 165 1 3 sky130_fd_sc_hd__tap_1 $T=189860 34480 1 180 $X=189210 $Y=34240
X132 166 167 1 3 sky130_fd_sc_hd__tap_1 $T=189860 39920 0 180 $X=189210 $Y=36960
X133 168 169 1 3 sky130_fd_sc_hd__tap_1 $T=189860 39920 1 180 $X=189210 $Y=39680
X134 170 171 1 3 sky130_fd_sc_hd__tap_1 $T=189860 45360 0 180 $X=189210 $Y=42400
X135 172 173 1 3 sky130_fd_sc_hd__tap_1 $T=189860 45360 1 180 $X=189210 $Y=45120
X136 174 175 1 3 sky130_fd_sc_hd__tap_1 $T=189860 50800 0 180 $X=189210 $Y=47840
X137 176 177 1 3 sky130_fd_sc_hd__tap_1 $T=189860 50800 1 180 $X=189210 $Y=50560
X138 178 179 1 3 sky130_fd_sc_hd__tap_1 $T=189860 56240 0 180 $X=189210 $Y=53280
X139 180 181 1 3 sky130_fd_sc_hd__tap_1 $T=189860 56240 1 180 $X=189210 $Y=56000
X140 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=29320 12720 1 0 $X=29130 $Y=9760
X141 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=29320 12720 0 0 $X=29130 $Y=12480
X142 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=29320 18160 1 0 $X=29130 $Y=15200
X143 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=29320 18160 0 0 $X=29130 $Y=17920
X144 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=29320 23600 1 0 $X=29130 $Y=20640
X145 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=29320 23600 0 0 $X=29130 $Y=23360
X146 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=44040 18160 1 0 $X=43850 $Y=15200
X147 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=44040 18160 0 0 $X=43850 $Y=17920
X148 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=44040 23600 1 0 $X=43850 $Y=20640
X149 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=44040 23600 0 0 $X=43850 $Y=23360
X150 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 12720 1 0 $X=58570 $Y=9760
X151 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 12720 0 0 $X=58570 $Y=12480
X152 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 18160 1 0 $X=58570 $Y=15200
X153 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 18160 0 0 $X=58570 $Y=17920
X154 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 23600 1 0 $X=58570 $Y=20640
X155 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 23600 0 0 $X=58570 $Y=23360
X156 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 29040 1 0 $X=58570 $Y=26080
X157 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 29040 0 0 $X=58570 $Y=28800
X158 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 12720 1 0 $X=73290 $Y=9760
X159 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 12720 0 0 $X=73290 $Y=12480
X160 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 18160 1 0 $X=73290 $Y=15200
X161 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 18160 0 0 $X=73290 $Y=17920
X162 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 23600 1 0 $X=73290 $Y=20640
X163 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 23600 0 0 $X=73290 $Y=23360
X164 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 29040 1 0 $X=73290 $Y=26080
X165 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 29040 0 0 $X=73290 $Y=28800
X166 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 12720 1 0 $X=88010 $Y=9760
X167 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 12720 0 0 $X=88010 $Y=12480
X168 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 18160 1 0 $X=88010 $Y=15200
X169 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 18160 0 0 $X=88010 $Y=17920
X170 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 23600 1 0 $X=88010 $Y=20640
X171 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 23600 0 0 $X=88010 $Y=23360
X172 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 29040 1 0 $X=88010 $Y=26080
X173 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 29040 0 0 $X=88010 $Y=28800
X174 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=102920 12720 1 0 $X=102730 $Y=9760
X175 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=102920 12720 0 0 $X=102730 $Y=12480
X176 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=102920 18160 1 0 $X=102730 $Y=15200
X177 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=102920 18160 0 0 $X=102730 $Y=17920
X178 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=102920 29040 1 0 $X=102730 $Y=26080
X179 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=102920 29040 0 0 $X=102730 $Y=28800
X180 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 12720 1 0 $X=117450 $Y=9760
X181 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 12720 0 0 $X=117450 $Y=12480
X182 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 18160 1 0 $X=117450 $Y=15200
X183 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 18160 0 0 $X=117450 $Y=17920
X184 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 23600 1 0 $X=117450 $Y=20640
X185 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 23600 0 0 $X=117450 $Y=23360
X186 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 29040 1 0 $X=117450 $Y=26080
X187 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 29040 0 0 $X=117450 $Y=28800
X188 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 34480 1 0 $X=117450 $Y=31520
X189 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 34480 0 0 $X=117450 $Y=34240
X190 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 39920 1 0 $X=117450 $Y=36960
X191 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 39920 0 0 $X=117450 $Y=39680
X192 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 45360 1 0 $X=117450 $Y=42400
X193 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 45360 0 0 $X=117450 $Y=45120
X194 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 50800 1 0 $X=117450 $Y=47840
X195 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 50800 0 0 $X=117450 $Y=50560
X196 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 56240 1 0 $X=117450 $Y=53280
X197 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 56240 0 0 $X=117450 $Y=56000
X198 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 12720 1 0 $X=132170 $Y=9760
X199 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 12720 0 0 $X=132170 $Y=12480
X200 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 23600 1 0 $X=132170 $Y=20640
X201 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 23600 0 0 $X=132170 $Y=23360
X202 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 29040 1 0 $X=132170 $Y=26080
X203 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 29040 0 0 $X=132170 $Y=28800
X204 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 34480 1 0 $X=132170 $Y=31520
X205 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 34480 0 0 $X=132170 $Y=34240
X206 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 39920 1 0 $X=132170 $Y=36960
X207 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 39920 0 0 $X=132170 $Y=39680
X208 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 45360 1 0 $X=132170 $Y=42400
X209 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 45360 0 0 $X=132170 $Y=45120
X210 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 50800 1 0 $X=132170 $Y=47840
X211 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 50800 0 0 $X=132170 $Y=50560
X212 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 56240 1 0 $X=132170 $Y=53280
X213 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 56240 0 0 $X=132170 $Y=56000
X214 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 12720 1 0 $X=146890 $Y=9760
X215 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 12720 0 0 $X=146890 $Y=12480
X216 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 18160 1 0 $X=146890 $Y=15200
X217 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 18160 0 0 $X=146890 $Y=17920
X218 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 23600 1 0 $X=146890 $Y=20640
X219 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 23600 0 0 $X=146890 $Y=23360
X220 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 34480 1 0 $X=146890 $Y=31520
X221 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 34480 0 0 $X=146890 $Y=34240
X222 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 39920 1 0 $X=146890 $Y=36960
X223 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 39920 0 0 $X=146890 $Y=39680
X224 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 45360 1 0 $X=146890 $Y=42400
X225 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 45360 0 0 $X=146890 $Y=45120
X226 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 50800 1 0 $X=146890 $Y=47840
X227 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 50800 0 0 $X=146890 $Y=50560
X228 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 56240 1 0 $X=146890 $Y=53280
X229 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 56240 0 0 $X=146890 $Y=56000
X230 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 12720 1 0 $X=161610 $Y=9760
X231 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 12720 0 0 $X=161610 $Y=12480
X232 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 18160 1 0 $X=161610 $Y=15200
X233 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 18160 0 0 $X=161610 $Y=17920
X234 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 23600 1 0 $X=161610 $Y=20640
X235 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 23600 0 0 $X=161610 $Y=23360
X236 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 34480 1 0 $X=161610 $Y=31520
X237 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 34480 0 0 $X=161610 $Y=34240
X238 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 39920 1 0 $X=161610 $Y=36960
X239 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 39920 0 0 $X=161610 $Y=39680
X240 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 45360 1 0 $X=161610 $Y=42400
X241 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 45360 0 0 $X=161610 $Y=45120
X242 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 50800 1 0 $X=161610 $Y=47840
X243 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 50800 0 0 $X=161610 $Y=50560
X244 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 56240 1 0 $X=161610 $Y=53280
X245 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 56240 0 0 $X=161610 $Y=56000
X246 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 18160 1 0 $X=176330 $Y=15200
X247 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 18160 0 0 $X=176330 $Y=17920
X248 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 23600 1 0 $X=176330 $Y=20640
X249 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 23600 0 0 $X=176330 $Y=23360
X250 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 34480 1 0 $X=176330 $Y=31520
X251 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 34480 0 0 $X=176330 $Y=34240
X252 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 39920 1 0 $X=176330 $Y=36960
X253 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 39920 0 0 $X=176330 $Y=39680
X254 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 45360 1 0 $X=176330 $Y=42400
X255 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 45360 0 0 $X=176330 $Y=45120
X256 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 50800 1 0 $X=176330 $Y=47840
X257 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 50800 0 0 $X=176330 $Y=50560
X258 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 56240 1 0 $X=176330 $Y=53280
X259 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 56240 0 0 $X=176330 $Y=56000
X260 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 12720 1 0 $X=188750 $Y=9760
X261 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 12720 0 0 $X=188750 $Y=12480
X262 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 18160 1 0 $X=188750 $Y=15200
X263 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 18160 0 0 $X=188750 $Y=17920
X264 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 23600 1 0 $X=188750 $Y=20640
X265 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 23600 0 0 $X=188750 $Y=23360
X266 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 29040 1 0 $X=188750 $Y=26080
X267 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 29040 0 0 $X=188750 $Y=28800
X268 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 34480 1 0 $X=188750 $Y=31520
X269 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 34480 0 0 $X=188750 $Y=34240
X270 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 39920 1 0 $X=188750 $Y=36960
X271 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 39920 0 0 $X=188750 $Y=39680
X272 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 45360 1 0 $X=188750 $Y=42400
X273 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 45360 0 0 $X=188750 $Y=45120
X274 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 50800 1 0 $X=188750 $Y=47840
X275 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 50800 0 0 $X=188750 $Y=50560
X276 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 56240 1 0 $X=188750 $Y=53280
X277 1 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=188940 56240 0 0 $X=188750 $Y=56000
X278 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 12720 1 0 $X=10270 $Y=9760
X279 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 12720 0 0 $X=10270 $Y=12480
X280 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 18160 1 0 $X=10270 $Y=15200
X281 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 18160 0 0 $X=10270 $Y=17920
X282 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 23600 1 0 $X=10270 $Y=20640
X283 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 23600 0 0 $X=10270 $Y=23360
X284 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 29040 1 0 $X=10270 $Y=26080
X285 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 29040 0 0 $X=10270 $Y=28800
X286 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 34480 1 0 $X=10270 $Y=31520
X287 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 34480 0 0 $X=10270 $Y=34240
X288 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 39920 1 0 $X=10270 $Y=36960
X289 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 39920 0 0 $X=10270 $Y=39680
X290 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 45360 1 0 $X=10270 $Y=42400
X291 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 45360 0 0 $X=10270 $Y=45120
X292 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 50800 1 0 $X=10270 $Y=47840
X293 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 50800 0 0 $X=10270 $Y=50560
X294 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 56240 1 0 $X=10270 $Y=53280
X295 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=10460 56240 0 0 $X=10270 $Y=56000
X296 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=15060 12720 0 0 $X=14870 $Y=12480
X297 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=15060 18160 1 0 $X=14870 $Y=15200
X298 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=15060 23600 0 0 $X=14870 $Y=23360
X299 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=24720 12720 0 0 $X=24530 $Y=12480
X300 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=24720 18160 1 0 $X=24530 $Y=15200
X301 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=26560 23600 0 0 $X=26370 $Y=23360
X302 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=29780 12720 0 0 $X=29590 $Y=12480
X303 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=38060 12720 0 0 $X=37870 $Y=12480
X304 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=41280 18160 1 0 $X=41090 $Y=15200
X305 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=44500 34480 1 0 $X=44310 $Y=31520
X306 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=47720 12720 0 0 $X=47530 $Y=12480
X307 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=54160 12720 0 0 $X=53970 $Y=12480
X308 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=56000 34480 1 0 $X=55810 $Y=31520
X309 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=61520 23600 1 0 $X=61330 $Y=20640
X310 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=62900 23600 0 0 $X=62710 $Y=23360
X311 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=77620 29040 0 0 $X=77430 $Y=28800
X312 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=84060 29040 0 0 $X=83870 $Y=28800
X313 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=88660 12720 1 0 $X=88470 $Y=9760
X314 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=88660 12720 0 0 $X=88470 $Y=12480
X315 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=88660 18160 1 0 $X=88470 $Y=15200
X316 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=98320 18160 1 0 $X=98130 $Y=15200
X317 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=98320 23600 0 0 $X=98130 $Y=23360
X318 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=100160 12720 0 0 $X=99970 $Y=12480
X319 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=103380 18160 0 0 $X=103190 $Y=17920
X320 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=114880 18160 1 0 $X=114690 $Y=15200
X321 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=114880 18160 0 0 $X=114690 $Y=17920
X322 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=121780 23600 1 0 $X=121590 $Y=20640
X323 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=129600 34480 1 0 $X=129410 $Y=31520
X324 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=138340 18160 1 0 $X=138150 $Y=15200
X325 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=142480 29040 1 0 $X=142290 $Y=26080
X326 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=147540 18160 1 0 $X=147350 $Y=15200
X327 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=147540 23600 1 0 $X=147350 $Y=20640
X328 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=157660 12720 1 0 $X=157470 $Y=9760
X329 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=171920 23600 0 0 $X=171730 $Y=23360
X330 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=172380 12720 1 0 $X=172190 $Y=9760
X331 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=184340 23600 1 0 $X=184150 $Y=20640
X332 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 12720 1 0 $X=185990 $Y=9760
X333 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 12720 0 0 $X=185990 $Y=12480
X334 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 18160 1 0 $X=185990 $Y=15200
X335 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 18160 0 0 $X=185990 $Y=17920
X336 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 29040 1 0 $X=185990 $Y=26080
X337 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 29040 0 0 $X=185990 $Y=28800
X338 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 34480 1 0 $X=185990 $Y=31520
X339 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 34480 0 0 $X=185990 $Y=34240
X340 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 39920 1 0 $X=185990 $Y=36960
X341 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 39920 0 0 $X=185990 $Y=39680
X342 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 45360 1 0 $X=185990 $Y=42400
X343 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 45360 0 0 $X=185990 $Y=45120
X344 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 50800 1 0 $X=185990 $Y=47840
X345 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 50800 0 0 $X=185990 $Y=50560
X346 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 56240 1 0 $X=185990 $Y=53280
X347 1 3 3 1 sky130_fd_sc_hd__decap_6 $T=186180 56240 0 0 $X=185990 $Y=56000
X348 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=17820 12720 0 0 $X=17630 $Y=12480
X349 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=17820 18160 1 0 $X=17630 $Y=15200
X350 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=19660 23600 0 0 $X=19470 $Y=23360
X351 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=27940 12720 1 0 $X=27750 $Y=9760
X352 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=27940 18160 0 0 $X=27750 $Y=17920
X353 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=27940 23600 1 0 $X=27750 $Y=20640
X354 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=42660 18160 0 0 $X=42470 $Y=17920
X355 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=42660 23600 1 0 $X=42470 $Y=20640
X356 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=42660 23600 0 0 $X=42470 $Y=23360
X357 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=44500 23600 1 0 $X=44310 $Y=20640
X358 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=44500 29040 1 0 $X=44310 $Y=26080
X359 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=44500 29040 0 0 $X=44310 $Y=28800
X360 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=46340 12720 1 0 $X=46150 $Y=9760
X361 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=47260 34480 1 0 $X=47070 $Y=31520
X362 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=48180 18160 0 0 $X=47990 $Y=17920
X363 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=48180 23600 0 0 $X=47990 $Y=23360
X364 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 18160 1 0 $X=57190 $Y=15200
X365 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 34480 0 0 $X=57190 $Y=34240
X366 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 39920 1 0 $X=57190 $Y=36960
X367 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 39920 0 0 $X=57190 $Y=39680
X368 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 45360 1 0 $X=57190 $Y=42400
X369 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 45360 0 0 $X=57190 $Y=45120
X370 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 50800 1 0 $X=57190 $Y=47840
X371 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 50800 0 0 $X=57190 $Y=50560
X372 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 56240 1 0 $X=57190 $Y=53280
X373 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=57380 56240 0 0 $X=57190 $Y=56000
X374 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=59220 12720 0 0 $X=59030 $Y=12480
X375 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=61060 12720 1 0 $X=60870 $Y=9760
X376 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=64280 12720 0 0 $X=64090 $Y=12480
X377 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=71180 12720 0 0 $X=70990 $Y=12480
X378 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=71180 23600 0 0 $X=70990 $Y=23360
X379 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=72100 18160 1 0 $X=71910 $Y=15200
X380 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=72100 18160 0 0 $X=71910 $Y=17920
X381 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=72100 29040 1 0 $X=71910 $Y=26080
X382 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=72100 29040 0 0 $X=71910 $Y=28800
X383 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=73940 18160 0 0 $X=73750 $Y=17920
X384 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=75780 23600 0 0 $X=75590 $Y=23360
X385 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=81300 12720 1 0 $X=81110 $Y=9760
X386 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=86820 12720 0 0 $X=86630 $Y=12480
X387 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=86820 18160 1 0 $X=86630 $Y=15200
X388 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=86820 29040 1 0 $X=86630 $Y=26080
X389 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=86820 29040 0 0 $X=86630 $Y=28800
X390 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=88660 23600 0 0 $X=88470 $Y=23360
X391 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=91420 12720 0 0 $X=91230 $Y=12480
X392 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=92340 18160 0 0 $X=92150 $Y=17920
X393 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=92340 29040 0 0 $X=92150 $Y=28800
X394 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=93260 18160 1 0 $X=93070 $Y=15200
X395 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=94180 23600 1 0 $X=93990 $Y=20640
X396 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=101540 29040 1 0 $X=101350 $Y=26080
X397 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=107980 18160 0 0 $X=107790 $Y=17920
X398 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=108900 12720 0 0 $X=108710 $Y=12480
X399 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=108900 18160 1 0 $X=108710 $Y=15200
X400 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=108900 23600 1 0 $X=108710 $Y=20640
X401 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=116260 12720 1 0 $X=116070 $Y=9760
X402 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=116260 23600 0 0 $X=116070 $Y=23360
X403 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=118100 29040 1 0 $X=117910 $Y=26080
X404 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=118100 29040 0 0 $X=117910 $Y=28800
X405 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=123160 29040 1 0 $X=122970 $Y=26080
X406 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 12720 1 0 $X=130790 $Y=9760
X407 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 12720 0 0 $X=130790 $Y=12480
X408 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 23600 0 0 $X=130790 $Y=23360
X409 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 34480 0 0 $X=130790 $Y=34240
X410 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 39920 1 0 $X=130790 $Y=36960
X411 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 39920 0 0 $X=130790 $Y=39680
X412 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 45360 1 0 $X=130790 $Y=42400
X413 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 45360 0 0 $X=130790 $Y=45120
X414 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 50800 1 0 $X=130790 $Y=47840
X415 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 50800 0 0 $X=130790 $Y=50560
X416 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 56240 1 0 $X=130790 $Y=53280
X417 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=130980 56240 0 0 $X=130790 $Y=56000
X418 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=132820 29040 1 0 $X=132630 $Y=26080
X419 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=136500 23600 0 0 $X=136310 $Y=23360
X420 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=136500 29040 0 0 $X=136310 $Y=28800
X421 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=140180 18160 0 0 $X=139990 $Y=17920
X422 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=141100 18160 1 0 $X=140910 $Y=15200
X423 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=144780 12720 0 0 $X=144590 $Y=12480
X424 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 12720 1 0 $X=145510 $Y=9760
X425 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 23600 1 0 $X=145510 $Y=20640
X426 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 34480 1 0 $X=145510 $Y=31520
X427 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 34480 0 0 $X=145510 $Y=34240
X428 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 39920 1 0 $X=145510 $Y=36960
X429 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 39920 0 0 $X=145510 $Y=39680
X430 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 45360 1 0 $X=145510 $Y=42400
X431 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 45360 0 0 $X=145510 $Y=45120
X432 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 50800 1 0 $X=145510 $Y=47840
X433 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 50800 0 0 $X=145510 $Y=50560
X434 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 56240 1 0 $X=145510 $Y=53280
X435 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=145700 56240 0 0 $X=145510 $Y=56000
X436 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=152140 18160 1 0 $X=151950 $Y=15200
X437 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=152140 23600 1 0 $X=151950 $Y=20640
X438 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 12720 1 0 $X=160230 $Y=9760
X439 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 12720 0 0 $X=160230 $Y=12480
X440 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 18160 0 0 $X=160230 $Y=17920
X441 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 23600 0 0 $X=160230 $Y=23360
X442 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 34480 1 0 $X=160230 $Y=31520
X443 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 34480 0 0 $X=160230 $Y=34240
X444 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 39920 1 0 $X=160230 $Y=36960
X445 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 39920 0 0 $X=160230 $Y=39680
X446 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 45360 1 0 $X=160230 $Y=42400
X447 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 45360 0 0 $X=160230 $Y=45120
X448 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 50800 1 0 $X=160230 $Y=47840
X449 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 50800 0 0 $X=160230 $Y=50560
X450 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 56240 1 0 $X=160230 $Y=53280
X451 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=160420 56240 0 0 $X=160230 $Y=56000
X452 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=167780 18160 1 0 $X=167590 $Y=15200
X453 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=167780 23600 0 0 $X=167590 $Y=23360
X454 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 12720 1 0 $X=174950 $Y=9760
X455 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 12720 0 0 $X=174950 $Y=12480
X456 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 23600 1 0 $X=174950 $Y=20640
X457 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 34480 1 0 $X=174950 $Y=31520
X458 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 34480 0 0 $X=174950 $Y=34240
X459 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 39920 1 0 $X=174950 $Y=36960
X460 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 39920 0 0 $X=174950 $Y=39680
X461 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 45360 1 0 $X=174950 $Y=42400
X462 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 45360 0 0 $X=174950 $Y=45120
X463 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 50800 1 0 $X=174950 $Y=47840
X464 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 50800 0 0 $X=174950 $Y=50560
X465 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 56240 1 0 $X=174950 $Y=53280
X466 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=175140 56240 0 0 $X=174950 $Y=56000
X467 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=178820 23600 0 0 $X=178630 $Y=23360
X468 1 3 3 1 sky130_fd_sc_hd__decap_3 $T=187560 23600 0 0 $X=187370 $Y=23360
X469 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 12720 1 0 $X=14870 $Y=9760
X470 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 18160 0 0 $X=14870 $Y=17920
X471 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 23600 1 0 $X=14870 $Y=20640
X472 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 29040 1 0 $X=14870 $Y=26080
X473 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 29040 0 0 $X=14870 $Y=28800
X474 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 34480 1 0 $X=14870 $Y=31520
X475 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 34480 0 0 $X=14870 $Y=34240
X476 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 39920 1 0 $X=14870 $Y=36960
X477 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 39920 0 0 $X=14870 $Y=39680
X478 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 45360 1 0 $X=14870 $Y=42400
X479 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 45360 0 0 $X=14870 $Y=45120
X480 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 50800 1 0 $X=14870 $Y=47840
X481 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 50800 0 0 $X=14870 $Y=50560
X482 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 56240 1 0 $X=14870 $Y=53280
X483 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=15060 56240 0 0 $X=14870 $Y=56000
X484 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 12720 1 0 $X=20390 $Y=9760
X485 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 18160 0 0 $X=20390 $Y=17920
X486 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 23600 1 0 $X=20390 $Y=20640
X487 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 29040 1 0 $X=20390 $Y=26080
X488 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 29040 0 0 $X=20390 $Y=28800
X489 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 34480 1 0 $X=20390 $Y=31520
X490 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 34480 0 0 $X=20390 $Y=34240
X491 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 39920 1 0 $X=20390 $Y=36960
X492 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 39920 0 0 $X=20390 $Y=39680
X493 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 45360 1 0 $X=20390 $Y=42400
X494 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 45360 0 0 $X=20390 $Y=45120
X495 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 50800 1 0 $X=20390 $Y=47840
X496 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 50800 0 0 $X=20390 $Y=50560
X497 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 56240 1 0 $X=20390 $Y=53280
X498 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=20580 56240 0 0 $X=20390 $Y=56000
X499 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=29780 18160 0 0 $X=29590 $Y=17920
X500 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=29780 23600 1 0 $X=29590 $Y=20640
X501 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=29780 23600 0 0 $X=29590 $Y=23360
X502 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 12720 1 0 $X=35110 $Y=9760
X503 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 18160 0 0 $X=35110 $Y=17920
X504 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 23600 1 0 $X=35110 $Y=20640
X505 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 23600 0 0 $X=35110 $Y=23360
X506 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 29040 0 0 $X=35110 $Y=28800
X507 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 34480 1 0 $X=35110 $Y=31520
X508 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 34480 0 0 $X=35110 $Y=34240
X509 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 39920 1 0 $X=35110 $Y=36960
X510 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 39920 0 0 $X=35110 $Y=39680
X511 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 45360 1 0 $X=35110 $Y=42400
X512 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 45360 0 0 $X=35110 $Y=45120
X513 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 50800 1 0 $X=35110 $Y=47840
X514 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 50800 0 0 $X=35110 $Y=50560
X515 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 56240 1 0 $X=35110 $Y=53280
X516 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=35300 56240 0 0 $X=35110 $Y=56000
X517 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=44500 39920 1 0 $X=44310 $Y=36960
X518 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=44500 39920 0 0 $X=44310 $Y=39680
X519 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=44500 45360 1 0 $X=44310 $Y=42400
X520 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=44500 45360 0 0 $X=44310 $Y=45120
X521 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=44500 50800 1 0 $X=44310 $Y=47840
X522 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=44500 50800 0 0 $X=44310 $Y=50560
X523 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=44500 56240 1 0 $X=44310 $Y=53280
X524 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=44500 56240 0 0 $X=44310 $Y=56000
X525 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=49560 29040 1 0 $X=49370 $Y=26080
X526 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=49560 29040 0 0 $X=49370 $Y=28800
X527 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=50020 39920 1 0 $X=49830 $Y=36960
X528 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=50020 39920 0 0 $X=49830 $Y=39680
X529 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=50020 45360 1 0 $X=49830 $Y=42400
X530 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=50020 45360 0 0 $X=49830 $Y=45120
X531 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=50020 50800 1 0 $X=49830 $Y=47840
X532 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=50020 50800 0 0 $X=49830 $Y=50560
X533 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=50020 56240 1 0 $X=49830 $Y=53280
X534 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=50020 56240 0 0 $X=49830 $Y=56000
X535 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=53240 12720 1 0 $X=53050 $Y=9760
X536 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 34480 1 0 $X=64550 $Y=31520
X537 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 34480 0 0 $X=64550 $Y=34240
X538 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 39920 1 0 $X=64550 $Y=36960
X539 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 39920 0 0 $X=64550 $Y=39680
X540 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 45360 1 0 $X=64550 $Y=42400
X541 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 45360 0 0 $X=64550 $Y=45120
X542 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 50800 1 0 $X=64550 $Y=47840
X543 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 50800 0 0 $X=64550 $Y=50560
X544 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 56240 1 0 $X=64550 $Y=53280
X545 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=64740 56240 0 0 $X=64550 $Y=56000
X546 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=66580 29040 0 0 $X=66390 $Y=28800
X547 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=67960 12720 1 0 $X=67770 $Y=9760
X548 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 12720 0 0 $X=73750 $Y=12480
X549 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 23600 1 0 $X=73750 $Y=20640
X550 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 29040 1 0 $X=73750 $Y=26080
X551 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 34480 1 0 $X=73750 $Y=31520
X552 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 34480 0 0 $X=73750 $Y=34240
X553 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 39920 1 0 $X=73750 $Y=36960
X554 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 39920 0 0 $X=73750 $Y=39680
X555 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 45360 1 0 $X=73750 $Y=42400
X556 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 45360 0 0 $X=73750 $Y=45120
X557 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 50800 1 0 $X=73750 $Y=47840
X558 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 50800 0 0 $X=73750 $Y=50560
X559 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 56240 1 0 $X=73750 $Y=53280
X560 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=73940 56240 0 0 $X=73750 $Y=56000
X561 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 12720 0 0 $X=79270 $Y=12480
X562 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 29040 1 0 $X=79270 $Y=26080
X563 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 34480 1 0 $X=79270 $Y=31520
X564 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 34480 0 0 $X=79270 $Y=34240
X565 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 39920 1 0 $X=79270 $Y=36960
X566 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 39920 0 0 $X=79270 $Y=39680
X567 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 45360 1 0 $X=79270 $Y=42400
X568 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 45360 0 0 $X=79270 $Y=45120
X569 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 50800 1 0 $X=79270 $Y=47840
X570 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 50800 0 0 $X=79270 $Y=50560
X571 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 56240 1 0 $X=79270 $Y=53280
X572 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=79460 56240 0 0 $X=79270 $Y=56000
X573 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=88660 23600 1 0 $X=88470 $Y=20640
X574 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=88660 29040 1 0 $X=88470 $Y=26080
X575 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 29040 1 0 $X=93990 $Y=26080
X576 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 34480 1 0 $X=93990 $Y=31520
X577 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 34480 0 0 $X=93990 $Y=34240
X578 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 39920 1 0 $X=93990 $Y=36960
X579 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 39920 0 0 $X=93990 $Y=39680
X580 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 45360 1 0 $X=93990 $Y=42400
X581 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 45360 0 0 $X=93990 $Y=45120
X582 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 50800 1 0 $X=93990 $Y=47840
X583 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 50800 0 0 $X=93990 $Y=50560
X584 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 56240 1 0 $X=93990 $Y=53280
X585 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=94180 56240 0 0 $X=93990 $Y=56000
X586 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=97400 29040 0 0 $X=97210 $Y=28800
X587 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 12720 1 0 $X=103190 $Y=9760
X588 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 29040 1 0 $X=103190 $Y=26080
X589 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 29040 0 0 $X=103190 $Y=28800
X590 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 34480 1 0 $X=103190 $Y=31520
X591 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 34480 0 0 $X=103190 $Y=34240
X592 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 39920 1 0 $X=103190 $Y=36960
X593 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 39920 0 0 $X=103190 $Y=39680
X594 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 45360 1 0 $X=103190 $Y=42400
X595 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 45360 0 0 $X=103190 $Y=45120
X596 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 50800 1 0 $X=103190 $Y=47840
X597 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 50800 0 0 $X=103190 $Y=50560
X598 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 56240 1 0 $X=103190 $Y=53280
X599 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=103380 56240 0 0 $X=103190 $Y=56000
X600 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 12720 1 0 $X=108710 $Y=9760
X601 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 29040 1 0 $X=108710 $Y=26080
X602 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 29040 0 0 $X=108710 $Y=28800
X603 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 34480 1 0 $X=108710 $Y=31520
X604 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 34480 0 0 $X=108710 $Y=34240
X605 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 39920 1 0 $X=108710 $Y=36960
X606 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 39920 0 0 $X=108710 $Y=39680
X607 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 45360 1 0 $X=108710 $Y=42400
X608 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 45360 0 0 $X=108710 $Y=45120
X609 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 50800 1 0 $X=108710 $Y=47840
X610 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 50800 0 0 $X=108710 $Y=50560
X611 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 56240 1 0 $X=108710 $Y=53280
X612 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=108900 56240 0 0 $X=108710 $Y=56000
X613 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 34480 0 0 $X=117910 $Y=34240
X614 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 39920 1 0 $X=117910 $Y=36960
X615 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 39920 0 0 $X=117910 $Y=39680
X616 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 45360 1 0 $X=117910 $Y=42400
X617 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 45360 0 0 $X=117910 $Y=45120
X618 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 50800 1 0 $X=117910 $Y=47840
X619 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 50800 0 0 $X=117910 $Y=50560
X620 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 56240 1 0 $X=117910 $Y=53280
X621 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=118100 56240 0 0 $X=117910 $Y=56000
X622 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=120400 34480 1 0 $X=120210 $Y=31520
X623 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=121780 12720 0 0 $X=121590 $Y=12480
X624 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123160 29040 0 0 $X=122970 $Y=28800
X625 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 12720 1 0 $X=123430 $Y=9760
X626 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 34480 0 0 $X=123430 $Y=34240
X627 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 39920 1 0 $X=123430 $Y=36960
X628 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 39920 0 0 $X=123430 $Y=39680
X629 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 45360 1 0 $X=123430 $Y=42400
X630 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 45360 0 0 $X=123430 $Y=45120
X631 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 50800 1 0 $X=123430 $Y=47840
X632 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 50800 0 0 $X=123430 $Y=50560
X633 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 56240 1 0 $X=123430 $Y=53280
X634 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=123620 56240 0 0 $X=123430 $Y=56000
X635 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=125460 18160 0 0 $X=125270 $Y=17920
X636 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=125460 23600 0 0 $X=125270 $Y=23360
X637 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 12720 1 0 $X=132630 $Y=9760
X638 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 34480 1 0 $X=132630 $Y=31520
X639 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 34480 0 0 $X=132630 $Y=34240
X640 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 39920 1 0 $X=132630 $Y=36960
X641 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 39920 0 0 $X=132630 $Y=39680
X642 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 45360 1 0 $X=132630 $Y=42400
X643 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 45360 0 0 $X=132630 $Y=45120
X644 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 50800 1 0 $X=132630 $Y=47840
X645 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 50800 0 0 $X=132630 $Y=50560
X646 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 56240 1 0 $X=132630 $Y=53280
X647 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=132820 56240 0 0 $X=132630 $Y=56000
X648 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 34480 1 0 $X=138150 $Y=31520
X649 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 34480 0 0 $X=138150 $Y=34240
X650 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 39920 1 0 $X=138150 $Y=36960
X651 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 39920 0 0 $X=138150 $Y=39680
X652 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 45360 1 0 $X=138150 $Y=42400
X653 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 45360 0 0 $X=138150 $Y=45120
X654 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 50800 1 0 $X=138150 $Y=47840
X655 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 50800 0 0 $X=138150 $Y=50560
X656 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 56240 1 0 $X=138150 $Y=53280
X657 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=138340 56240 0 0 $X=138150 $Y=56000
X658 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=141560 23600 0 0 $X=141370 $Y=23360
X659 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=141560 29040 0 0 $X=141370 $Y=28800
X660 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 12720 0 0 $X=147350 $Y=12480
X661 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 18160 0 0 $X=147350 $Y=17920
X662 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 34480 1 0 $X=147350 $Y=31520
X663 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 34480 0 0 $X=147350 $Y=34240
X664 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 39920 1 0 $X=147350 $Y=36960
X665 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 39920 0 0 $X=147350 $Y=39680
X666 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 45360 1 0 $X=147350 $Y=42400
X667 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 45360 0 0 $X=147350 $Y=45120
X668 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 50800 1 0 $X=147350 $Y=47840
X669 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 50800 0 0 $X=147350 $Y=50560
X670 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 56240 1 0 $X=147350 $Y=53280
X671 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=147540 56240 0 0 $X=147350 $Y=56000
X672 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 12720 0 0 $X=152870 $Y=12480
X673 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 29040 0 0 $X=152870 $Y=28800
X674 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 34480 1 0 $X=152870 $Y=31520
X675 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 34480 0 0 $X=152870 $Y=34240
X676 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 39920 1 0 $X=152870 $Y=36960
X677 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 39920 0 0 $X=152870 $Y=39680
X678 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 45360 1 0 $X=152870 $Y=42400
X679 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 45360 0 0 $X=152870 $Y=45120
X680 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 50800 1 0 $X=152870 $Y=47840
X681 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 50800 0 0 $X=152870 $Y=50560
X682 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 56240 1 0 $X=152870 $Y=53280
X683 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=153060 56240 0 0 $X=152870 $Y=56000
X684 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 12720 0 0 $X=162070 $Y=12480
X685 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 23600 0 0 $X=162070 $Y=23360
X686 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 29040 1 0 $X=162070 $Y=26080
X687 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 29040 0 0 $X=162070 $Y=28800
X688 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 34480 1 0 $X=162070 $Y=31520
X689 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 34480 0 0 $X=162070 $Y=34240
X690 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 39920 1 0 $X=162070 $Y=36960
X691 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 39920 0 0 $X=162070 $Y=39680
X692 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 45360 1 0 $X=162070 $Y=42400
X693 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 45360 0 0 $X=162070 $Y=45120
X694 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 50800 1 0 $X=162070 $Y=47840
X695 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 50800 0 0 $X=162070 $Y=50560
X696 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 56240 1 0 $X=162070 $Y=53280
X697 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=162260 56240 0 0 $X=162070 $Y=56000
X698 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 29040 1 0 $X=167590 $Y=26080
X699 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 29040 0 0 $X=167590 $Y=28800
X700 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 34480 1 0 $X=167590 $Y=31520
X701 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 34480 0 0 $X=167590 $Y=34240
X702 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 39920 1 0 $X=167590 $Y=36960
X703 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 39920 0 0 $X=167590 $Y=39680
X704 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 45360 1 0 $X=167590 $Y=42400
X705 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 45360 0 0 $X=167590 $Y=45120
X706 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 50800 1 0 $X=167590 $Y=47840
X707 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 50800 0 0 $X=167590 $Y=50560
X708 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 56240 1 0 $X=167590 $Y=53280
X709 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=167780 56240 0 0 $X=167590 $Y=56000
X710 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 18160 0 0 $X=176790 $Y=17920
X711 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 34480 1 0 $X=176790 $Y=31520
X712 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 34480 0 0 $X=176790 $Y=34240
X713 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 39920 1 0 $X=176790 $Y=36960
X714 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 39920 0 0 $X=176790 $Y=39680
X715 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 45360 1 0 $X=176790 $Y=42400
X716 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 45360 0 0 $X=176790 $Y=45120
X717 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 50800 1 0 $X=176790 $Y=47840
X718 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 50800 0 0 $X=176790 $Y=50560
X719 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 56240 1 0 $X=176790 $Y=53280
X720 1 3 3 1 sky130_fd_sc_hd__decap_12 $T=176980 56240 0 0 $X=176790 $Y=56000
X721 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=17820 23600 0 0 $X=17630 $Y=23360
X722 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=26100 12720 1 0 $X=25910 $Y=9760
X723 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=26100 18160 0 0 $X=25910 $Y=17920
X724 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=26100 23600 1 0 $X=25910 $Y=20640
X725 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=27480 12720 0 0 $X=27290 $Y=12480
X726 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=27480 18160 1 0 $X=27290 $Y=15200
X727 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 12720 1 0 $X=40630 $Y=9760
X728 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 12720 0 0 $X=40630 $Y=12480
X729 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 18160 0 0 $X=40630 $Y=17920
X730 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 23600 1 0 $X=40630 $Y=20640
X731 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 23600 0 0 $X=40630 $Y=23360
X732 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 29040 1 0 $X=40630 $Y=26080
X733 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 29040 0 0 $X=40630 $Y=28800
X734 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 34480 1 0 $X=40630 $Y=31520
X735 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 34480 0 0 $X=40630 $Y=34240
X736 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 39920 1 0 $X=40630 $Y=36960
X737 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 39920 0 0 $X=40630 $Y=39680
X738 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 45360 1 0 $X=40630 $Y=42400
X739 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 45360 0 0 $X=40630 $Y=45120
X740 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 50800 1 0 $X=40630 $Y=47840
X741 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 50800 0 0 $X=40630 $Y=50560
X742 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 56240 1 0 $X=40630 $Y=53280
X743 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=40820 56240 0 0 $X=40630 $Y=56000
X744 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=44500 12720 1 0 $X=44310 $Y=9760
X745 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=48180 18160 1 0 $X=47990 $Y=15200
X746 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=49560 23600 1 0 $X=49370 $Y=20640
X747 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 34480 0 0 $X=55350 $Y=34240
X748 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 39920 1 0 $X=55350 $Y=36960
X749 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 39920 0 0 $X=55350 $Y=39680
X750 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 45360 1 0 $X=55350 $Y=42400
X751 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 45360 0 0 $X=55350 $Y=45120
X752 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 50800 1 0 $X=55350 $Y=47840
X753 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 50800 0 0 $X=55350 $Y=50560
X754 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 56240 1 0 $X=55350 $Y=53280
X755 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=55540 56240 0 0 $X=55350 $Y=56000
X756 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=56920 12720 0 0 $X=56730 $Y=12480
X757 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=56920 18160 0 0 $X=56730 $Y=17920
X758 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=56920 23600 0 0 $X=56730 $Y=23360
X759 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=59220 12720 1 0 $X=59030 $Y=9760
X760 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=64280 23600 1 0 $X=64090 $Y=20640
X761 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=66580 18160 1 0 $X=66390 $Y=15200
X762 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=66580 18160 0 0 $X=66390 $Y=17920
X763 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=66580 29040 1 0 $X=66390 $Y=26080
X764 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 34480 1 0 $X=70070 $Y=31520
X765 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 34480 0 0 $X=70070 $Y=34240
X766 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 39920 1 0 $X=70070 $Y=36960
X767 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 39920 0 0 $X=70070 $Y=39680
X768 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 45360 1 0 $X=70070 $Y=42400
X769 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 45360 0 0 $X=70070 $Y=45120
X770 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 50800 1 0 $X=70070 $Y=47840
X771 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 50800 0 0 $X=70070 $Y=50560
X772 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 56240 1 0 $X=70070 $Y=53280
X773 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=70260 56240 0 0 $X=70070 $Y=56000
X774 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=73940 23600 0 0 $X=73750 $Y=23360
X775 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=79460 12720 1 0 $X=79270 $Y=9760
X776 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=79460 18160 1 0 $X=79270 $Y=15200
X777 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=84980 12720 0 0 $X=84790 $Y=12480
X778 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=84980 18160 1 0 $X=84790 $Y=15200
X779 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=84980 29040 1 0 $X=84790 $Y=26080
X780 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=86360 18160 0 0 $X=86170 $Y=17920
X781 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=91420 18160 1 0 $X=91230 $Y=15200
X782 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 29040 1 0 $X=99510 $Y=26080
X783 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 34480 1 0 $X=99510 $Y=31520
X784 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 34480 0 0 $X=99510 $Y=34240
X785 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 39920 1 0 $X=99510 $Y=36960
X786 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 39920 0 0 $X=99510 $Y=39680
X787 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 45360 1 0 $X=99510 $Y=42400
X788 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 45360 0 0 $X=99510 $Y=45120
X789 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 50800 1 0 $X=99510 $Y=47840
X790 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 50800 0 0 $X=99510 $Y=50560
X791 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 56240 1 0 $X=99510 $Y=53280
X792 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=99700 56240 0 0 $X=99510 $Y=56000
X793 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=101080 18160 1 0 $X=100890 $Y=15200
X794 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=101080 18160 0 0 $X=100890 $Y=17920
X795 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=101080 23600 0 0 $X=100890 $Y=23360
X796 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=106140 18160 0 0 $X=105950 $Y=17920
X797 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=114420 12720 1 0 $X=114230 $Y=9760
X798 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=115800 12720 0 0 $X=115610 $Y=12480
X799 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=123620 18160 1 0 $X=123430 $Y=15200
X800 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 12720 1 0 $X=128950 $Y=9760
X801 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 18160 1 0 $X=128950 $Y=15200
X802 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 34480 0 0 $X=128950 $Y=34240
X803 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 39920 1 0 $X=128950 $Y=36960
X804 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 39920 0 0 $X=128950 $Y=39680
X805 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 45360 1 0 $X=128950 $Y=42400
X806 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 45360 0 0 $X=128950 $Y=45120
X807 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 50800 1 0 $X=128950 $Y=47840
X808 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 50800 0 0 $X=128950 $Y=50560
X809 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 56240 1 0 $X=128950 $Y=53280
X810 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=129140 56240 0 0 $X=128950 $Y=56000
X811 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=132820 18160 1 0 $X=132630 $Y=15200
X812 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 12720 1 0 $X=143670 $Y=9760
X813 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 34480 1 0 $X=143670 $Y=31520
X814 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 34480 0 0 $X=143670 $Y=34240
X815 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 39920 1 0 $X=143670 $Y=36960
X816 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 39920 0 0 $X=143670 $Y=39680
X817 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 45360 1 0 $X=143670 $Y=42400
X818 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 45360 0 0 $X=143670 $Y=45120
X819 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 50800 1 0 $X=143670 $Y=47840
X820 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 50800 0 0 $X=143670 $Y=50560
X821 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 56240 1 0 $X=143670 $Y=53280
X822 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=143860 56240 0 0 $X=143670 $Y=56000
X823 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=145240 29040 1 0 $X=145050 $Y=26080
X824 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=150300 18160 1 0 $X=150110 $Y=15200
X825 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=150300 23600 1 0 $X=150110 $Y=20640
X826 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=153060 23600 0 0 $X=152870 $Y=23360
X827 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 12720 0 0 $X=158390 $Y=12480
X828 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 23600 0 0 $X=158390 $Y=23360
X829 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 29040 0 0 $X=158390 $Y=28800
X830 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 34480 1 0 $X=158390 $Y=31520
X831 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 34480 0 0 $X=158390 $Y=34240
X832 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 39920 1 0 $X=158390 $Y=36960
X833 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 39920 0 0 $X=158390 $Y=39680
X834 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 45360 1 0 $X=158390 $Y=42400
X835 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 45360 0 0 $X=158390 $Y=45120
X836 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 50800 1 0 $X=158390 $Y=47840
X837 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 50800 0 0 $X=158390 $Y=50560
X838 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 56240 1 0 $X=158390 $Y=53280
X839 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=158580 56240 0 0 $X=158390 $Y=56000
X840 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 23600 1 0 $X=173110 $Y=20640
X841 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 34480 1 0 $X=173110 $Y=31520
X842 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 34480 0 0 $X=173110 $Y=34240
X843 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 39920 1 0 $X=173110 $Y=36960
X844 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 39920 0 0 $X=173110 $Y=39680
X845 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 45360 1 0 $X=173110 $Y=42400
X846 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 45360 0 0 $X=173110 $Y=45120
X847 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 50800 1 0 $X=173110 $Y=47840
X848 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 50800 0 0 $X=173110 $Y=50560
X849 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 56240 1 0 $X=173110 $Y=53280
X850 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=173300 56240 0 0 $X=173110 $Y=56000
X851 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=174680 18160 0 0 $X=174490 $Y=17920
X852 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=174680 23600 0 0 $X=174490 $Y=23360
X853 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=176980 23600 0 0 $X=176790 $Y=23360
X854 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=185720 23600 0 0 $X=185530 $Y=23360
X855 1 3 3 1 sky130_fd_sc_hd__decap_4 $T=187100 23600 1 0 $X=186910 $Y=20640
X856 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=44500 18160 0 0 $X=44310 $Y=17920
X857 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=44500 23600 0 0 $X=44310 $Y=23360
X858 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=44500 34480 0 0 $X=44310 $Y=34240
X859 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=55080 29040 1 0 $X=54890 $Y=26080
X860 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=55080 29040 0 0 $X=54890 $Y=28800
X861 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=59220 23600 0 0 $X=59030 $Y=23360
X862 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=84520 23600 0 0 $X=84330 $Y=23360
X863 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=88660 18160 0 0 $X=88470 $Y=17920
X864 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=88660 29040 0 0 $X=88470 $Y=28800
X865 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=96480 12720 0 0 $X=96290 $Y=12480
X866 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=108900 23600 0 0 $X=108710 $Y=23360
X867 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=118100 23600 1 0 $X=117910 $Y=20640
X868 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=125920 34480 1 0 $X=125730 $Y=31520
X869 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=127300 12720 0 0 $X=127110 $Y=12480
X870 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=128680 29040 0 0 $X=128490 $Y=28800
X871 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=132820 23600 0 0 $X=132630 $Y=23360
X872 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=132820 29040 0 0 $X=132630 $Y=28800
X873 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=142020 23600 1 0 $X=141830 $Y=20640
X874 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=153060 29040 1 0 $X=152870 $Y=26080
X875 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=153980 12720 1 0 $X=153790 $Y=9760
X876 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=168700 12720 1 0 $X=168510 $Y=9760
X877 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=171460 12720 0 0 $X=171270 $Y=12480
X878 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 12720 1 0 $X=182310 $Y=9760
X879 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 12720 0 0 $X=182310 $Y=12480
X880 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 18160 1 0 $X=182310 $Y=15200
X881 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 18160 0 0 $X=182310 $Y=17920
X882 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 29040 1 0 $X=182310 $Y=26080
X883 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 29040 0 0 $X=182310 $Y=28800
X884 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 34480 1 0 $X=182310 $Y=31520
X885 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 34480 0 0 $X=182310 $Y=34240
X886 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 39920 1 0 $X=182310 $Y=36960
X887 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 39920 0 0 $X=182310 $Y=39680
X888 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 45360 1 0 $X=182310 $Y=42400
X889 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 45360 0 0 $X=182310 $Y=45120
X890 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 50800 1 0 $X=182310 $Y=47840
X891 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 50800 0 0 $X=182310 $Y=50560
X892 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 56240 1 0 $X=182310 $Y=53280
X893 1 3 3 1 sky130_fd_sc_hd__decap_8 $T=182500 56240 0 0 $X=182310 $Y=56000
X894 1 3 3 1 sky130_fd_sc_hd__fill_1 $T=35300 18160 1 0 $X=35110 $Y=15200
X895 1 3 3 1 sky130_fd_sc_hd__fill_1 $T=96940 12720 1 0 $X=96750 $Y=9760
X896 1 3 3 1 sky130_fd_sc_hd__fill_1 $T=131900 23600 1 0 $X=131710 $Y=20640
X897 1 3 3 1 sky130_fd_sc_hd__fill_1 $T=131900 29040 1 0 $X=131710 $Y=26080
X898 1 3 3 1 sky130_fd_sc_hd__fill_1 $T=132820 23600 1 0 $X=132630 $Y=20640
X899 1 3 3 1 sky130_fd_sc_hd__fill_1 $T=169620 23600 1 0 $X=169430 $Y=20640
X900 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=44500 12720 0 0 $X=44310 $Y=12480
X901 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=59220 23600 1 0 $X=59030 $Y=20640
X902 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=72560 12720 0 0 $X=72370 $Y=12480
X903 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=72560 23600 0 0 $X=72370 $Y=23360
X904 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=90040 23600 0 0 $X=89850 $Y=23360
X905 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=110280 18160 1 0 $X=110090 $Y=15200
X906 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=118100 34480 1 0 $X=117910 $Y=31520
X907 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=134200 29040 1 0 $X=134010 $Y=26080
X908 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=138340 12720 0 0 $X=138150 $Y=12480
X909 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=141560 18160 0 0 $X=141370 $Y=17920
X910 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=146160 12720 0 0 $X=145970 $Y=12480
X911 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=146160 18160 1 0 $X=145970 $Y=15200
X912 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=146160 18160 0 0 $X=145970 $Y=17920
X913 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=147540 12720 1 0 $X=147350 $Y=9760
X914 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=160880 18160 1 0 $X=160690 $Y=15200
X915 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=160880 23600 1 0 $X=160690 $Y=20640
X916 1 3 3 1 sky130_fd_sc_hd__fill_2 $T=162260 12720 1 0 $X=162070 $Y=9760
X917 15 L1M1_PR $T=20350 13910 0 0 $X=20205 $Y=13795
X918 17 L1M1_PR $T=20350 16970 0 0 $X=20205 $Y=16855
X919 14 L1M1_PR $T=21270 14250 0 0 $X=21125 $Y=14135
X920 16 L1M1_PR $T=21270 16630 0 0 $X=21125 $Y=16515
X921 19 L1M1_PR $T=22190 24790 0 0 $X=22045 $Y=24675
X922 18 L1M1_PR $T=23110 25130 0 0 $X=22965 $Y=25015
X923 21 L1M1_PR $T=30930 11530 0 0 $X=30785 $Y=11415
X924 23 L1M1_PR $T=30930 16970 0 0 $X=30785 $Y=16855
X925 20 L1M1_PR $T=31850 11190 0 0 $X=31705 $Y=11075
X926 22 L1M1_PR $T=31850 16630 0 0 $X=31705 $Y=16515
X927 24 L1M1_PR $T=35070 14250 0 0 $X=34925 $Y=14135
X928 25 L1M1_PR $T=37830 13910 0 0 $X=37685 $Y=13795
X929 26 L1M1_PR $T=37830 27510 0 0 $X=37685 $Y=27395
X930 28 L1M1_PR $T=39210 16630 0 0 $X=39065 $Y=16515
X931 29 L1M1_PR $T=40590 16970 0 0 $X=40445 $Y=16855
X932 27 L1M1_PR $T=40590 27850 0 0 $X=40445 $Y=27735
X933 7 L1M1_PR $T=44730 16970 0 0 $X=44585 $Y=16855
X934 5 L1M1_PR $T=45420 16970 0 0 $X=45275 $Y=16855
X935 7 L1M1_PR $T=45650 14930 0 0 $X=45505 $Y=14815
X936 21 L1M1_PR $T=45675 13910 0 0 $X=45530 $Y=13795
X937 5 L1M1_PR $T=46110 13910 0 0 $X=45965 $Y=13795
X938 15 L1M1_PR $T=46110 17310 0 0 $X=45965 $Y=17195
X939 7 L1M1_PR $T=46110 22410 0 0 $X=45965 $Y=22295
X940 7 L1M1_PR $T=46110 27850 0 0 $X=45965 $Y=27735
X941 7 L1M1_PR $T=46110 30230 0 0 $X=45965 $Y=30115
X942 25 L1M1_PR $T=46570 16970 0 0 $X=46425 $Y=16855
X943 5 L1M1_PR $T=46800 22410 0 0 $X=46655 $Y=22295
X944 5 L1M1_PR $T=46800 27850 0 0 $X=46655 $Y=27735
X945 5 L1M1_PR $T=46800 30230 0 0 $X=46655 $Y=30115
X946 109 L1M1_PR $T=47260 16970 0 0 $X=47115 $Y=16855
X947 19 L1M1_PR $T=47260 27850 0 0 $X=47115 $Y=27735
X948 82 L1M1_PR $T=47490 14930 0 0 $X=47345 $Y=14815
X949 17 L1M1_PR $T=47490 22750 0 0 $X=47345 $Y=22635
X950 23 L1M1_PR $T=47490 30230 0 0 $X=47345 $Y=30115
X951 80 L1M1_PR $T=47950 17650 0 0 $X=47805 $Y=17535
X952 23 L1M1_PR $T=47950 22410 0 0 $X=47805 $Y=22295
X953 27 L1M1_PR $T=47950 28190 0 0 $X=47805 $Y=28075
X954 29 L1M1_PR $T=47950 29890 0 0 $X=47805 $Y=29775
X955 9 L1M1_PR $T=48410 36010 0 0 $X=48265 $Y=35895
X956 109 L1M1_PR $T=48640 22410 0 0 $X=48495 $Y=22295
X957 109 L1M1_PR $T=48640 27850 0 0 $X=48495 $Y=27735
X958 109 L1M1_PR $T=48640 30230 0 0 $X=48495 $Y=30115
X959 31 L1M1_PR $T=48870 11530 0 0 $X=48725 $Y=11415
X960 9 L1M1_PR $T=48870 32950 0 0 $X=48725 $Y=32835
X961 81 L1M1_PR $T=49330 23090 0 0 $X=49185 $Y=22975
X962 78 L1M1_PR $T=49330 28530 0 0 $X=49185 $Y=28415
X963 79 L1M1_PR $T=49330 31250 0 0 $X=49185 $Y=31135
X964 30 L1M1_PR $T=49715 11190 0 0 $X=49570 $Y=11075
X965 78 L1M1_PR $T=49715 35330 0 0 $X=49570 $Y=35215
X966 9 L1M1_PR $T=49790 19350 0 0 $X=49645 $Y=19235
X967 9 L1M1_PR $T=49790 24790 0 0 $X=49645 $Y=24675
X968 79 L1M1_PR $T=50175 33290 0 0 $X=50030 $Y=33175
X969 9 L1M1_PR $T=50250 16970 0 0 $X=50105 $Y=16855
X970 7 L1M1_PR $T=50740 13910 0 0 $X=50595 $Y=13795
X971 80 L1M1_PR $T=51095 19010 0 0 $X=50950 $Y=18895
X972 81 L1M1_PR $T=51095 24450 0 0 $X=50950 $Y=24335
X973 5 L1M1_PR $T=51175 13910 0 0 $X=51030 $Y=13795
X974 82 L1M1_PR $T=51555 16970 0 0 $X=51410 $Y=16855
X975 11 L1M1_PR $T=51630 22410 0 0 $X=51485 $Y=22295
X976 21 L1M1_PR $T=52090 13570 0 0 $X=51945 $Y=13455
X977 31 L1M1_PR $T=52550 13570 0 0 $X=52405 $Y=13455
X978 83 L1M1_PR $T=52935 22750 0 0 $X=52790 $Y=22635
X979 109 L1M1_PR $T=53240 13910 0 0 $X=53095 $Y=13795
X980 85 L1M1_PR $T=53930 14930 0 0 $X=53785 $Y=14815
X981 23 L1M1_PR $T=55310 34990 0 0 $X=55165 $Y=34875
X982 27 L1M1_PR $T=55770 32270 0 0 $X=55625 $Y=32155
X983 21 L1M1_PR $T=56690 18670 0 0 $X=56545 $Y=18555
X984 19 L1M1_PR $T=56690 24110 0 0 $X=56545 $Y=23995
X985 15 L1M1_PR $T=57150 15950 0 0 $X=57005 $Y=15835
X986 33 L1M1_PR $T=58530 21390 0 0 $X=58385 $Y=21275
X987 9 L1M1_PR $T=59450 16970 0 0 $X=59305 $Y=16855
X988 9 L1M1_PR $T=59450 19350 0 0 $X=59305 $Y=19235
X989 9 L1M1_PR $T=59450 27850 0 0 $X=59305 $Y=27735
X990 9 L1M1_PR $T=59450 30230 0 0 $X=59305 $Y=30115
X991 9 L1M1_PR $T=60370 23090 0 0 $X=60225 $Y=22975
X992 84 L1M1_PR $T=60755 16970 0 0 $X=60610 $Y=16855
X993 85 L1M1_PR $T=60755 19010 0 0 $X=60610 $Y=18895
X994 86 L1M1_PR $T=60755 27850 0 0 $X=60610 $Y=27735
X995 87 L1M1_PR $T=60755 29890 0 0 $X=60610 $Y=29775
X996 84 L1M1_PR $T=60830 14930 0 0 $X=60685 $Y=14815
X997 10 L1M1_PR $T=61290 22410 0 0 $X=61145 $Y=22295
X998 109 L1M1_PR $T=61520 13910 0 0 $X=61375 $Y=13795
X999 33 L1M1_PR $T=62210 13570 0 0 $X=62065 $Y=13455
X1000 33 L1M1_PR $T=62670 11530 0 0 $X=62525 $Y=11415
X1001 25 L1M1_PR $T=62670 13910 0 0 $X=62525 $Y=13795
X1002 5 L1M1_PR $T=63360 13910 0 0 $X=63215 $Y=13795
X1003 7 L1M1_PR $T=64050 13910 0 0 $X=63905 $Y=13795
X1004 32 L1M1_PR $T=65430 11190 0 0 $X=65285 $Y=11075
X1005 37 L1M1_PR $T=65890 24790 0 0 $X=65745 $Y=24675
X1006 31 L1M1_PR $T=66350 15950 0 0 $X=66205 $Y=15835
X1007 25 L1M1_PR $T=66350 18670 0 0 $X=66205 $Y=18555
X1008 11 L1M1_PR $T=66350 22410 0 0 $X=66205 $Y=22295
X1009 37 L1M1_PR $T=66350 26830 0 0 $X=66205 $Y=26715
X1010 29 L1M1_PR $T=66350 31250 0 0 $X=66205 $Y=31135
X1011 35 L1M1_PR $T=66810 13910 0 0 $X=66665 $Y=13795
X1012 88 L1M1_PR $T=67655 22410 0 0 $X=67510 $Y=22295
X1013 34 L1M1_PR $T=68190 14250 0 0 $X=68045 $Y=14135
X1014 86 L1M1_PR $T=68650 17650 0 0 $X=68505 $Y=17535
X1015 83 L1M1_PR $T=68650 20370 0 0 $X=68505 $Y=20255
X1016 87 L1M1_PR $T=68650 28530 0 0 $X=68505 $Y=28415
X1017 109 L1M1_PR $T=69340 16970 0 0 $X=69195 $Y=16855
X1018 109 L1M1_PR $T=69340 19350 0 0 $X=69195 $Y=19235
X1019 109 L1M1_PR $T=69340 27850 0 0 $X=69195 $Y=27735
X1020 35 L1M1_PR $T=70030 16970 0 0 $X=69885 $Y=16855
X1021 41 L1M1_PR $T=70030 19010 0 0 $X=69885 $Y=18895
X1022 36 L1M1_PR $T=70030 24450 0 0 $X=69885 $Y=24335
X1023 37 L1M1_PR $T=70030 27850 0 0 $X=69885 $Y=27735
X1024 29 L1M1_PR $T=70490 17310 0 0 $X=70345 $Y=17195
X1025 31 L1M1_PR $T=70490 19350 0 0 $X=70345 $Y=19235
X1026 27 L1M1_PR $T=70490 28190 0 0 $X=70345 $Y=28075
X1027 5 L1M1_PR $T=71180 27850 0 0 $X=71035 $Y=27735
X1028 5 L1M1_PR $T=71265 16970 0 0 $X=71120 $Y=16855
X1029 5 L1M1_PR $T=71265 19350 0 0 $X=71120 $Y=19235
X1030 7 L1M1_PR $T=71835 16970 0 0 $X=71690 $Y=16855
X1031 7 L1M1_PR $T=71870 19350 0 0 $X=71725 $Y=19235
X1032 7 L1M1_PR $T=71870 27850 0 0 $X=71725 $Y=27735
X1033 39 L1M1_PR $T=73250 23090 0 0 $X=73105 $Y=22975
X1034 39 L1M1_PR $T=74170 11530 0 0 $X=74025 $Y=11415
X1035 41 L1M1_PR $T=74170 16970 0 0 $X=74025 $Y=16855
X1036 7 L1M1_PR $T=74170 30230 0 0 $X=74025 $Y=30115
X1037 5 L1M1_PR $T=74860 30230 0 0 $X=74715 $Y=30115
X1038 11 L1M1_PR $T=75550 19350 0 0 $X=75405 $Y=19235
X1039 37 L1M1_PR $T=75550 29890 0 0 $X=75405 $Y=29775
X1040 39 L1M1_PR $T=76010 29890 0 0 $X=75865 $Y=29775
X1041 40 L1M1_PR $T=76470 16630 0 0 $X=76325 $Y=16515
X1042 109 L1M1_PR $T=76700 30230 0 0 $X=76555 $Y=30115
X1043 89 L1M1_PR $T=76855 19010 0 0 $X=76710 $Y=18895
X1044 11 L1M1_PR $T=77390 25130 0 0 $X=77245 $Y=25015
X1045 90 L1M1_PR $T=77390 29550 0 0 $X=77245 $Y=29435
X1046 38 L1M1_PR $T=78310 11190 0 0 $X=78165 $Y=11075
X1047 90 L1M1_PR $T=78695 24450 0 0 $X=78550 $Y=24335
X1048 10 L1M1_PR $T=79690 22410 0 0 $X=79545 $Y=22295
X1049 11 L1M1_PR $T=80610 23090 0 0 $X=80465 $Y=22975
X1050 7 L1M1_PR $T=80610 30230 0 0 $X=80465 $Y=30115
X1051 11 L1M1_PR $T=81070 22410 0 0 $X=80925 $Y=22295
X1052 5 L1M1_PR $T=81300 30230 0 0 $X=81155 $Y=30115
X1053 89 L1M1_PR $T=81530 17650 0 0 $X=81385 $Y=17535
X1054 39 L1M1_PR $T=81990 29830 0 0 $X=81845 $Y=29715
X1055 109 L1M1_PR $T=82220 16970 0 0 $X=82075 $Y=16855
X1056 91 L1M1_PR $T=82405 22750 0 0 $X=82260 $Y=22635
X1057 41 L1M1_PR $T=82450 18670 0 0 $X=82305 $Y=18555
X1058 47 L1M1_PR $T=82490 29890 0 0 $X=82345 $Y=29775
X1059 43 L1M1_PR $T=82910 11530 0 0 $X=82765 $Y=11415
X1060 43 L1M1_PR $T=82910 16970 0 0 $X=82765 $Y=16855
X1061 7 L1M1_PR $T=82910 19350 0 0 $X=82765 $Y=19235
X1062 109 L1M1_PR $T=83140 30230 0 0 $X=82995 $Y=30115
X1063 33 L1M1_PR $T=83370 16970 0 0 $X=83225 $Y=16855
X1064 5 L1M1_PR $T=83600 19350 0 0 $X=83455 $Y=19235
X1065 91 L1M1_PR $T=83830 29550 0 0 $X=83685 $Y=29435
X1066 5 L1M1_PR $T=84060 16970 0 0 $X=83915 $Y=16855
X1067 35 L1M1_PR $T=84290 19010 0 0 $X=84145 $Y=18895
X1068 35 L1M1_PR $T=84290 24110 0 0 $X=84145 $Y=23995
X1069 7 L1M1_PR $T=84750 16970 0 0 $X=84605 $Y=16855
X1070 45 L1M1_PR $T=84750 19350 0 0 $X=84605 $Y=19235
X1071 109 L1M1_PR $T=85440 19350 0 0 $X=85295 $Y=19235
X1072 88 L1M1_PR $T=86130 20370 0 0 $X=85985 $Y=20255
X1073 42 L1M1_PR $T=87050 11190 0 0 $X=86905 $Y=11075
X1074 45 L1M1_PR $T=87970 21390 0 0 $X=87825 $Y=21275
X1075 11 L1M1_PR $T=91190 24790 0 0 $X=91045 $Y=24675
X1076 45 L1M1_PR $T=91650 11530 0 0 $X=91505 $Y=11415
X1077 92 L1M1_PR $T=92495 24450 0 0 $X=92350 $Y=24335
X1078 7 L1M1_PR $T=93030 13910 0 0 $X=92885 $Y=13795
X1079 44 L1M1_PR $T=93490 11190 0 0 $X=93345 $Y=11075
X1080 5 L1M1_PR $T=93720 13910 0 0 $X=93575 $Y=13795
X1081 11 L1M1_PR $T=93950 19690 0 0 $X=93805 $Y=19575
X1082 7 L1M1_PR $T=93950 30230 0 0 $X=93805 $Y=30115
X1083 45 L1M1_PR $T=94410 13910 0 0 $X=94265 $Y=13795
X1084 5 L1M1_PR $T=94640 30230 0 0 $X=94495 $Y=30115
X1085 49 L1M1_PR $T=94870 13570 0 0 $X=94725 $Y=13455
X1086 93 L1M1_PR $T=94870 17650 0 0 $X=94725 $Y=17535
X1087 93 L1M1_PR $T=95255 19010 0 0 $X=95110 $Y=18895
X1088 43 L1M1_PR $T=95330 29890 0 0 $X=95185 $Y=29775
X1089 109 L1M1_PR $T=95560 13910 0 0 $X=95415 $Y=13795
X1090 109 L1M1_PR $T=95560 16970 0 0 $X=95415 $Y=16855
X1091 11 L1M1_PR $T=95790 22410 0 0 $X=95645 $Y=22295
X1092 53 L1M1_PR $T=95790 30230 0 0 $X=95645 $Y=30115
X1093 92 L1M1_PR $T=96245 13230 0 0 $X=96100 $Y=13115
X1094 51 L1M1_PR $T=96250 16970 0 0 $X=96105 $Y=16855
X1095 109 L1M1_PR $T=96480 30230 0 0 $X=96335 $Y=30115
X1096 41 L1M1_PR $T=96710 17310 0 0 $X=96565 $Y=17195
X1097 94 L1M1_PR $T=97095 22750 0 0 $X=96950 $Y=22635
X1098 94 L1M1_PR $T=97170 29550 0 0 $X=97025 $Y=29435
X1099 5 L1M1_PR $T=97485 16970 0 0 $X=97340 $Y=16855
X1100 7 L1M1_PR $T=98090 16970 0 0 $X=97945 $Y=16855
X1101 47 L1M1_PR $T=98090 24110 0 0 $X=97945 $Y=23995
X1102 47 L1M1_PR $T=98550 11530 0 0 $X=98405 $Y=11415
X1103 46 L1M1_PR $T=99470 11190 0 0 $X=99325 $Y=11075
X1104 43 L1M1_PR $T=100850 18670 0 0 $X=100705 $Y=18555
X1105 43 L1M1_PR $T=100850 20370 0 0 $X=100705 $Y=20255
X1106 51 L1M1_PR $T=102690 21390 0 0 $X=102545 $Y=21275
X1107 49 L1M1_PR $T=103610 13910 0 0 $X=103465 $Y=13795
X1108 51 L1M1_PR $T=103610 16970 0 0 $X=103465 $Y=16855
X1109 48 L1M1_PR $T=105450 14250 0 0 $X=105305 $Y=14135
X1110 50 L1M1_PR $T=105450 16630 0 0 $X=105305 $Y=16515
X1111 52 L1M1_PR $T=110510 19010 0 0 $X=110365 $Y=18895
X1112 12 L1M1_PR $T=110510 22410 0 0 $X=110365 $Y=22295
X1113 7 L1M1_PR $T=111430 16970 0 0 $X=111285 $Y=16855
X1114 95 L1M1_PR $T=111815 22750 0 0 $X=111670 $Y=22635
X1115 5 L1M1_PR $T=112120 16970 0 0 $X=111975 $Y=16855
X1116 51 L1M1_PR $T=112810 16970 0 0 $X=112665 $Y=16855
X1117 7 L1M1_PR $T=112810 24790 0 0 $X=112665 $Y=24675
X1118 59 L1M1_PR $T=113270 17310 0 0 $X=113125 $Y=17195
X1119 5 L1M1_PR $T=113500 24790 0 0 $X=113355 $Y=24675
X1120 54 L1M1_PR $T=113730 14250 0 0 $X=113585 $Y=14135
X1121 109 L1M1_PR $T=113960 16970 0 0 $X=113815 $Y=16855
X1122 77 L1M1_PR $T=114190 24450 0 0 $X=114045 $Y=24335
X1123 95 L1M1_PR $T=114650 17650 0 0 $X=114505 $Y=17535
X1124 53 L1M1_PR $T=114650 19350 0 0 $X=114505 $Y=19235
X1125 19 L1M1_PR $T=114650 24790 0 0 $X=114505 $Y=24675
X1126 109 L1M1_PR $T=115340 24790 0 0 $X=115195 $Y=24675
X1127 55 L1M1_PR $T=115570 13910 0 0 $X=115425 $Y=13795
X1128 97 L1M1_PR $T=116030 24110 0 0 $X=115885 $Y=23995
X1129 53 L1M1_PR $T=117410 21390 0 0 $X=117265 $Y=21275
X1130 7 L1M1_PR $T=118330 13910 0 0 $X=118185 $Y=13795
X1131 12 L1M1_PR $T=118330 19690 0 0 $X=118185 $Y=19575
X1132 12 L1M1_PR $T=118330 24790 0 0 $X=118185 $Y=24675
X1133 5 L1M1_PR $T=119070 13910 0 0 $X=118925 $Y=13795
X1134 47 L1M1_PR $T=119635 13570 0 0 $X=119490 $Y=13455
X1135 96 L1M1_PR $T=119635 19010 0 0 $X=119490 $Y=18895
X1136 97 L1M1_PR $T=119635 24450 0 0 $X=119490 $Y=24335
X1137 109 L1M1_PR $T=119635 32270 0 0 $X=119490 $Y=32155
X1138 7 L1M1_PR $T=119710 27850 0 0 $X=119565 $Y=27735
X1139 7 L1M1_PR $T=119710 30230 0 0 $X=119565 $Y=30115
X1140 55 L1M1_PR $T=120170 13570 0 0 $X=120025 $Y=13455
X1141 6 L1M1_PR $T=120170 33290 0 0 $X=120025 $Y=33175
X1142 5 L1M1_PR $T=120400 27850 0 0 $X=120255 $Y=27735
X1143 5 L1M1_PR $T=120400 30230 0 0 $X=120255 $Y=30115
X1144 58 L1M1_PR $T=120630 16630 0 0 $X=120485 $Y=16515
X1145 109 L1M1_PR $T=120910 13910 0 0 $X=120765 $Y=13795
X1146 75 L1M1_PR $T=121090 27850 0 0 $X=120945 $Y=27735
X1147 53 L1M1_PR $T=121090 29890 0 0 $X=120945 $Y=29775
X1148 56 L1M1_PR $T=121550 11190 0 0 $X=121405 $Y=11075
X1149 96 L1M1_PR $T=121550 13230 0 0 $X=121405 $Y=13115
X1150 17 L1M1_PR $T=121550 28190 0 0 $X=121405 $Y=28075
X1151 63 L1M1_PR $T=121550 29890 0 0 $X=121405 $Y=29775
X1152 109 L1M1_PR $T=122240 27850 0 0 $X=122095 $Y=27735
X1153 109 L1M1_PR $T=122240 30230 0 0 $X=122095 $Y=30115
X1154 59 L1M1_PR $T=122470 16970 0 0 $X=122325 $Y=16855
X1155 57 L1M1_PR $T=122930 11530 0 0 $X=122785 $Y=11415
X1156 99 L1M1_PR $T=122930 28530 0 0 $X=122785 $Y=28415
X1157 98 L1M1_PR $T=122930 29550 0 0 $X=122785 $Y=29435
X1158 12 L1M1_PR $T=124770 22410 0 0 $X=124625 $Y=22295
X1159 12 L1M1_PR $T=124770 27510 0 0 $X=124625 $Y=27395
X1160 49 L1M1_PR $T=125230 18670 0 0 $X=125085 $Y=18555
X1161 17 L1M1_PR $T=125230 25810 0 0 $X=125085 $Y=25695
X1162 7 L1M1_PR $T=125690 16970 0 0 $X=125545 $Y=16855
X1163 98 L1M1_PR $T=126075 22750 0 0 $X=125930 $Y=22635
X1164 99 L1M1_PR $T=126075 28190 0 0 $X=125930 $Y=28075
X1165 5 L1M1_PR $T=126290 16970 0 0 $X=126145 $Y=16855
X1166 49 L1M1_PR $T=127070 17310 0 0 $X=126925 $Y=17195
X1167 57 L1M1_PR $T=127530 16970 0 0 $X=127385 $Y=16855
X1168 109 L1M1_PR $T=128220 16970 0 0 $X=128075 $Y=16855
X1169 100 L1M1_PR $T=128910 17650 0 0 $X=128765 $Y=17535
X1170 59 L1M1_PR $T=131670 21390 0 0 $X=131525 $Y=21275
X1171 77 L1M1_PR $T=131670 26830 0 0 $X=131525 $Y=26715
X1172 77 L1M1_PR $T=131670 28530 0 0 $X=131525 $Y=28415
X1173 12 L1M1_PR $T=133050 19690 0 0 $X=132905 $Y=19575
X1174 10 L1M1_PR $T=133510 22410 0 0 $X=133365 $Y=22295
X1175 61 L1M1_PR $T=133970 13910 0 0 $X=133825 $Y=13795
X1176 100 L1M1_PR $T=134355 19350 0 0 $X=134210 $Y=19235
X1177 12 L1M1_PR $T=134430 23090 0 0 $X=134285 $Y=22975
X1178 60 L1M1_PR $T=134890 14250 0 0 $X=134745 $Y=14135
X1179 7 L1M1_PR $T=134890 16970 0 0 $X=134745 $Y=16855
X1180 12 L1M1_PR $T=134890 22410 0 0 $X=134745 $Y=22295
X1181 12 L1M1_PR $T=135350 27510 0 0 $X=135205 $Y=27395
X1182 5 L1M1_PR $T=135580 16970 0 0 $X=135435 $Y=16855
X1183 101 L1M1_PR $T=136195 22750 0 0 $X=136050 $Y=22635
X1184 55 L1M1_PR $T=136270 17310 0 0 $X=136125 $Y=17195
X1185 61 L1M1_PR $T=136655 16970 0 0 $X=136510 $Y=16855
X1186 102 L1M1_PR $T=136655 28190 0 0 $X=136510 $Y=28075
X1187 109 L1M1_PR $T=137420 16970 0 0 $X=137275 $Y=16855
X1188 104 L1M1_PR $T=138110 17650 0 0 $X=137965 $Y=17535
X1189 101 L1M1_PR $T=138110 24110 0 0 $X=137965 $Y=23995
X1190 102 L1M1_PR $T=138110 29550 0 0 $X=137965 $Y=29435
X1191 109 L1M1_PR $T=138800 24790 0 0 $X=138655 $Y=24675
X1192 109 L1M1_PR $T=138800 30230 0 0 $X=138655 $Y=30115
X1193 63 L1M1_PR $T=139490 11530 0 0 $X=139345 $Y=11415
X1194 67 L1M1_PR $T=139490 24450 0 0 $X=139345 $Y=24335
X1195 71 L1M1_PR $T=139490 30230 0 0 $X=139345 $Y=30115
X1196 55 L1M1_PR $T=139950 18670 0 0 $X=139805 $Y=18555
X1197 59 L1M1_PR $T=139950 24790 0 0 $X=139805 $Y=24675
X1198 63 L1M1_PR $T=139950 29890 0 0 $X=139805 $Y=29775
X1199 62 L1M1_PR $T=140410 11190 0 0 $X=140265 $Y=11075
X1200 5 L1M1_PR $T=140640 24790 0 0 $X=140495 $Y=24675
X1201 5 L1M1_PR $T=140640 30230 0 0 $X=140495 $Y=30115
X1202 7 L1M1_PR $T=141330 24790 0 0 $X=141185 $Y=24675
X1203 7 L1M1_PR $T=141330 30230 0 0 $X=141185 $Y=30115
X1204 63 L1M1_PR $T=141790 23090 0 0 $X=141645 $Y=22975
X1205 67 L1M1_PR $T=142250 26830 0 0 $X=142105 $Y=26715
X1206 64 L1M1_PR $T=142710 14250 0 0 $X=142565 $Y=14135
X1207 7 L1M1_PR $T=142710 16970 0 0 $X=142565 $Y=16855
X1208 7 L1M1_PR $T=142710 19350 0 0 $X=142565 $Y=19235
X1209 5 L1M1_PR $T=143175 16970 0 0 $X=143030 $Y=16855
X1210 5 L1M1_PR $T=143400 19350 0 0 $X=143255 $Y=19235
X1211 57 L1M1_PR $T=144090 16970 0 0 $X=143945 $Y=16855
X1212 61 L1M1_PR $T=144090 19350 0 0 $X=143945 $Y=19235
X1213 65 L1M1_PR $T=144550 13910 0 0 $X=144405 $Y=13795
X1214 69 L1M1_PR $T=144550 19350 0 0 $X=144405 $Y=19235
X1215 65 L1M1_PR $T=144695 16970 0 0 $X=144550 $Y=16855
X1216 109 L1M1_PR $T=145240 19350 0 0 $X=145095 $Y=19235
X1217 109 L1M1_PR $T=145290 16970 0 0 $X=145145 $Y=16855
X1218 103 L1M1_PR $T=145930 17650 0 0 $X=145785 $Y=17535
X1219 107 L1M1_PR $T=145930 18670 0 0 $X=145785 $Y=18555
X1220 69 L1M1_PR $T=148690 11530 0 0 $X=148545 $Y=11415
X1221 66 L1M1_PR $T=150990 25130 0 0 $X=150845 $Y=25015
X1222 67 L1M1_PR $T=151910 24790 0 0 $X=151765 $Y=24675
X1223 68 L1M1_PR $T=152830 11190 0 0 $X=152685 $Y=11075
X1224 13 L1M1_PR $T=153290 19350 0 0 $X=153145 $Y=19235
X1225 13 L1M1_PR $T=153750 16970 0 0 $X=153605 $Y=16855
X1226 13 L1M1_PR $T=153750 22070 0 0 $X=153605 $Y=21955
X1227 103 L1M1_PR $T=154595 19010 0 0 $X=154450 $Y=18895
X1228 104 L1M1_PR $T=155055 16970 0 0 $X=154910 $Y=16855
X1229 105 L1M1_PR $T=155055 22750 0 0 $X=154910 $Y=22635
X1230 105 L1M1_PR $T=155130 24110 0 0 $X=154985 $Y=23995
X1231 109 L1M1_PR $T=155820 24790 0 0 $X=155675 $Y=24675
X1232 75 L1M1_PR $T=156510 24450 0 0 $X=156365 $Y=24335
X1233 67 L1M1_PR $T=156970 24790 0 0 $X=156825 $Y=24675
X1234 7 L1M1_PR $T=156970 27850 0 0 $X=156825 $Y=27735
X1235 5 L1M1_PR $T=157660 24790 0 0 $X=157515 $Y=24675
X1236 5 L1M1_PR $T=157660 27850 0 0 $X=157515 $Y=27735
X1237 7 L1M1_PR $T=158350 24790 0 0 $X=158205 $Y=24675
X1238 71 L1M1_PR $T=158350 28190 0 0 $X=158205 $Y=28075
X1239 77 L1M1_PR $T=158810 28190 0 0 $X=158665 $Y=28075
X1240 109 L1M1_PR $T=159500 27850 0 0 $X=159355 $Y=27735
X1241 61 L1M1_PR $T=160190 20370 0 0 $X=160045 $Y=20255
X1242 106 L1M1_PR $T=160190 26830 0 0 $X=160045 $Y=26715
X1243 57 L1M1_PR $T=160650 15950 0 0 $X=160505 $Y=15835
X1244 71 L1M1_PR $T=160650 23090 0 0 $X=160505 $Y=22975
X1245 71 L1M1_PR $T=162490 16970 0 0 $X=162345 $Y=16855
X1246 4 L1M1_PR $T=162490 19350 0 0 $X=162345 $Y=19235
X1247 13 L1M1_PR $T=162490 22410 0 0 $X=162345 $Y=22295
X1248 106 L1M1_PR $T=163795 22750 0 0 $X=163650 $Y=22635
X1249 73 L1M1_PR $T=164330 11530 0 0 $X=164185 $Y=11415
X1250 70 L1M1_PR $T=164790 16630 0 0 $X=164645 $Y=16515
X1251 72 L1M1_PR $T=165250 11190 0 0 $X=165105 $Y=11075
X1252 2 L1M1_PR $T=165250 19010 0 0 $X=165105 $Y=18895
X1253 13 L1M1_PR $T=165710 19350 0 0 $X=165565 $Y=19235
X1254 2 L1M1_PR $T=167015 19010 0 0 $X=166870 $Y=18895
X1255 4 L1M1_PR $T=168010 14930 0 0 $X=167865 $Y=14815
X1256 109 L1M1_PR $T=168700 13910 0 0 $X=168555 $Y=13795
X1257 73 L1M1_PR $T=169390 13570 0 0 $X=169245 $Y=13455
X1258 13 L1M1_PR $T=169390 16970 0 0 $X=169245 $Y=16855
X1259 75 L1M1_PR $T=169390 21390 0 0 $X=169245 $Y=21275
X1260 75 L1M1_PR $T=169390 23090 0 0 $X=169245 $Y=22975
X1261 108 L1M1_PR $T=169390 24450 0 0 $X=169245 $Y=24335
X1262 65 L1M1_PR $T=169850 13910 0 0 $X=169705 $Y=13795
X1263 10 L1M1_PR $T=170310 22410 0 0 $X=170165 $Y=22295
X1264 7 L1M1_PR $T=170310 24790 0 0 $X=170165 $Y=24675
X1265 6 L1M1_PR $T=170540 13910 0 0 $X=170395 $Y=13795
X1266 107 L1M1_PR $T=170725 16970 0 0 $X=170580 $Y=16855
X1267 8 L1M1_PR $T=171230 13910 0 0 $X=171085 $Y=13795
X1268 13 L1M1_PR $T=171230 21730 0 0 $X=171085 $Y=21615
X1269 69 L1M1_PR $T=171230 24110 0 0 $X=171085 $Y=23995
X1270 5 L1M1_PR $T=171690 24790 0 0 $X=171545 $Y=24675
X1271 6 L1M1_PR $T=172150 22750 0 0 $X=172005 $Y=22635
X1272 69 L1M1_PR $T=172610 20030 0 0 $X=172465 $Y=19915
X1273 5 L1M1_PR $T=173070 22750 0 0 $X=172925 $Y=22635
X1274 8 L1M1_PR $T=173530 19350 0 0 $X=173385 $Y=19235
X1275 7 L1M1_PR $T=173990 20370 0 0 $X=173845 $Y=20255
X1276 65 L1M1_PR $T=176290 15950 0 0 $X=176145 $Y=15835
X1277 75 L1M1_PR $T=177210 16970 0 0 $X=177065 $Y=16855
X1278 13 L1M1_PR $T=177210 22070 0 0 $X=177065 $Y=21955
X1279 108 L1M1_PR $T=178515 22750 0 0 $X=178370 $Y=22635
X1280 74 L1M1_PR $T=179050 16630 0 0 $X=178905 $Y=16515
X1281 77 L1M1_PR $T=181350 24790 0 0 $X=181205 $Y=24675
X1282 73 L1M1_PR $T=184110 21390 0 0 $X=183965 $Y=21275
X1283 76 L1M1_PR $T=184570 24450 0 0 $X=184425 $Y=24335
X1284 5 M1M2_PR_M $T=43350 13570 0 0 $X=43190 $Y=13440
X1285 15 M1M2_PR_M $T=43350 14250 0 0 $X=43190 $Y=14120
X1286 7 M1M2_PR_M $T=43350 16290 0 0 $X=43190 $Y=16160
X1287 19 M1M2_PR_M $T=46110 24450 0 0 $X=45950 $Y=24320
X1288 21 M1M2_PR_M $T=48870 13570 0 0 $X=48710 $Y=13440
X1289 29 M1M2_PR_M $T=70950 17650 0 0 $X=70790 $Y=17520
X1290 7 M1M2_PR_M $T=109590 14590 0 0 $X=109430 $Y=14460
X1291 5 M1M2_PR_M $T=112350 27170 0 0 $X=112190 $Y=27040
X1292 7 M1M2_PR_M $T=128910 16290 0 0 $X=128750 $Y=16160
X1293 109 M1M2_PR_M $T=148230 16970 0 0 $X=148070 $Y=16840
X1294 16 M1M2_PR $T=10230 16630 0 0 $X=10070 $Y=16470
X1295 14 M1M2_PR $T=15750 14250 0 0 $X=15590 $Y=14090
X1296 18 M1M2_PR $T=18510 25130 0 0 $X=18350 $Y=24970
X1297 20 M1M2_PR $T=26790 11190 0 0 $X=26630 $Y=11030
X1298 22 M1M2_PR $T=29550 16630 0 0 $X=29390 $Y=16470
X1299 17 M1M2_PR $T=29550 17310 0 0 $X=29390 $Y=17150
X1300 17 M1M2_PR $T=29550 22750 0 0 $X=29390 $Y=22590
X1301 23 M1M2_PR $T=32310 17310 0 0 $X=32150 $Y=17150
X1302 23 M1M2_PR $T=32310 21390 0 0 $X=32150 $Y=21230
X1303 24 M1M2_PR $T=35070 14250 0 0 $X=34910 $Y=14090
X1304 15 M1M2_PR $T=35070 14930 0 0 $X=34910 $Y=14770
X1305 15 M1M2_PR $T=35070 17650 0 0 $X=34910 $Y=17490
X1306 26 M1M2_PR $T=37830 27510 0 0 $X=37670 $Y=27350
X1307 28 M1M2_PR $T=40590 650 0 0 $X=40430 $Y=490
X1308 28 M1M2_PR $T=40590 16290 0 0 $X=40430 $Y=16130
X1309 29 M1M2_PR $T=40590 16970 0 0 $X=40430 $Y=16810
X1310 17 M1M2_PR $T=40590 22750 0 0 $X=40430 $Y=22590
X1311 29 M1M2_PR $T=40590 29890 0 0 $X=40430 $Y=29730
X1312 17 M1M2_PR $T=40590 38390 0 0 $X=40430 $Y=38230
X1313 15 M1M2_PR $T=42890 9490 0 0 $X=42730 $Y=9330
X1314 7 M1M2_PR $T=43350 14930 0 0 $X=43190 $Y=14770
X1315 5 M1M2_PR $T=43350 17310 0 0 $X=43190 $Y=17150
X1316 5 M1M2_PR $T=43350 22070 0 0 $X=43190 $Y=21910
X1317 5 M1M2_PR $T=43350 27510 0 0 $X=43190 $Y=27350
X1318 5 M1M2_PR $T=43350 30570 0 0 $X=43190 $Y=30410
X1319 21 M1M2_PR $T=46110 11530 0 0 $X=45950 $Y=11370
X1320 25 M1M2_PR $T=46110 13230 0 0 $X=45950 $Y=13070
X1321 21 M1M2_PR $T=46110 14590 0 0 $X=45950 $Y=14430
X1322 25 M1M2_PR $T=46110 15950 0 0 $X=45950 $Y=15790
X1323 7 M1M2_PR $T=46110 16630 0 0 $X=45950 $Y=16470
X1324 7 M1M2_PR $T=46110 22410 0 0 $X=45950 $Y=22250
X1325 23 M1M2_PR $T=46110 23090 0 0 $X=45950 $Y=22930
X1326 19 M1M2_PR $T=46110 26830 0 0 $X=45950 $Y=26670
X1327 7 M1M2_PR $T=46110 27850 0 0 $X=45950 $Y=27690
X1328 7 M1M2_PR $T=46110 29550 0 0 $X=45950 $Y=29390
X1329 7 M1M2_PR $T=46110 30230 0 0 $X=45950 $Y=30070
X1330 23 M1M2_PR $T=46110 30910 0 0 $X=45950 $Y=30750
X1331 28 M1M2_PR $T=48410 650 0 0 $X=48250 $Y=490
X1332 15 M1M2_PR $T=48410 9490 0 0 $X=48250 $Y=9330
X1333 21 M1M2_PR $T=48525 14590 0 0 $X=48365 $Y=14430
X1334 21 M1M2_PR $T=48525 18670 0 0 $X=48365 $Y=18510
X1335 30 M1M2_PR $T=48870 10510 0 0 $X=48710 $Y=10350
X1336 15 M1M2_PR $T=48870 15950 0 0 $X=48710 $Y=15790
X1337 9 M1M2_PR $T=48870 16970 0 0 $X=48710 $Y=16810
X1338 9 M1M2_PR $T=48870 19350 0 0 $X=48710 $Y=19190
X1339 9 M1M2_PR $T=48870 24790 0 0 $X=48710 $Y=24630
X1340 9 M1M2_PR $T=48870 32950 0 0 $X=48710 $Y=32790
X1341 9 M1M2_PR $T=48870 35670 0 0 $X=48710 $Y=35510
X1342 31 M1M2_PR $T=51630 12210 0 0 $X=51470 $Y=12050
X1343 31 M1M2_PR $T=51630 13230 0 0 $X=51470 $Y=13070
X1344 7 M1M2_PR $T=51630 14250 0 0 $X=51470 $Y=14090
X1345 82 M1M2_PR $T=51630 14930 0 0 $X=51470 $Y=14770
X1346 82 M1M2_PR $T=51630 16970 0 0 $X=51470 $Y=16810
X1347 80 M1M2_PR $T=51630 17650 0 0 $X=51470 $Y=17490
X1348 80 M1M2_PR $T=51630 19010 0 0 $X=51470 $Y=18850
X1349 109 M1M2_PR $T=51630 21390 0 0 $X=51470 $Y=21230
X1350 81 M1M2_PR $T=51630 23090 0 0 $X=51470 $Y=22930
X1351 81 M1M2_PR $T=51630 24450 0 0 $X=51470 $Y=24290
X1352 109 M1M2_PR $T=51630 27510 0 0 $X=51470 $Y=27350
X1353 78 M1M2_PR $T=51630 28530 0 0 $X=51470 $Y=28370
X1354 79 M1M2_PR $T=51630 31250 0 0 $X=51470 $Y=31090
X1355 79 M1M2_PR $T=51630 33290 0 0 $X=51470 $Y=33130
X1356 78 M1M2_PR $T=51630 35330 0 0 $X=51470 $Y=35170
X1357 85 M1M2_PR $T=54390 14930 0 0 $X=54230 $Y=14770
X1358 85 M1M2_PR $T=54390 19010 0 0 $X=54230 $Y=18850
X1359 83 M1M2_PR $T=54390 20370 0 0 $X=54230 $Y=20210
X1360 83 M1M2_PR $T=54390 22750 0 0 $X=54230 $Y=22590
X1361 109 M1M2_PR $T=54390 27510 0 0 $X=54230 $Y=27350
X1362 109 M1M2_PR $T=54390 30230 0 0 $X=54230 $Y=30070
X1363 23 M1M2_PR $T=54390 30910 0 0 $X=54230 $Y=30750
X1364 23 M1M2_PR $T=54390 34990 0 0 $X=54230 $Y=34830
X1365 109 M1M2_PR $T=57150 13910 0 0 $X=56990 $Y=13750
X1366 109 M1M2_PR $T=57150 17310 0 0 $X=56990 $Y=17150
X1367 109 M1M2_PR $T=57150 18670 0 0 $X=56990 $Y=18510
X1368 109 M1M2_PR $T=57150 21390 0 0 $X=56990 $Y=21230
X1369 36 M1M2_PR $T=57150 24110 0 0 $X=56990 $Y=23950
X1370 27 M1M2_PR $T=57150 28190 0 0 $X=56990 $Y=28030
X1371 27 M1M2_PR $T=57150 32270 0 0 $X=56990 $Y=32110
X1372 5 M1M2_PR $T=59910 14250 0 0 $X=59750 $Y=14090
X1373 9 M1M2_PR $T=59910 16970 0 0 $X=59750 $Y=16810
X1374 9 M1M2_PR $T=59910 19350 0 0 $X=59750 $Y=19190
X1375 9 M1M2_PR $T=59910 23090 0 0 $X=59750 $Y=22930
X1376 9 M1M2_PR $T=59910 27850 0 0 $X=59750 $Y=27690
X1377 9 M1M2_PR $T=59910 30230 0 0 $X=59750 $Y=30070
X1378 33 M1M2_PR $T=62670 11530 0 0 $X=62510 $Y=11370
X1379 33 M1M2_PR $T=62670 13230 0 0 $X=62510 $Y=13070
X1380 25 M1M2_PR $T=62670 13910 0 0 $X=62510 $Y=13750
X1381 84 M1M2_PR $T=62670 14930 0 0 $X=62510 $Y=14770
X1382 84 M1M2_PR $T=62670 16970 0 0 $X=62510 $Y=16810
X1383 25 M1M2_PR $T=62670 18670 0 0 $X=62510 $Y=18510
X1384 33 M1M2_PR $T=62670 21390 0 0 $X=62510 $Y=21230
X1385 37 M1M2_PR $T=62670 25470 0 0 $X=62510 $Y=25310
X1386 37 M1M2_PR $T=62670 26830 0 0 $X=62510 $Y=26670
X1387 87 M1M2_PR $T=62670 28530 0 0 $X=62510 $Y=28370
X1388 87 M1M2_PR $T=62670 29890 0 0 $X=62510 $Y=29730
X1389 32 M1M2_PR $T=65430 11190 0 0 $X=65270 $Y=11030
X1390 31 M1M2_PR $T=65430 12210 0 0 $X=65270 $Y=12050
X1391 31 M1M2_PR $T=65430 15950 0 0 $X=65270 $Y=15790
X1392 31 M1M2_PR $T=65430 19690 0 0 $X=65270 $Y=19530
X1393 11 M1M2_PR $T=65430 22410 0 0 $X=65270 $Y=22250
X1394 109 M1M2_PR $T=65430 27510 0 0 $X=65270 $Y=27350
X1395 109 M1M2_PR $T=65430 32610 0 0 $X=65270 $Y=32450
X1396 34 M1M2_PR $T=68190 14250 0 0 $X=68030 $Y=14090
X1397 35 M1M2_PR $T=68190 14930 0 0 $X=68030 $Y=14770
X1398 35 M1M2_PR $T=68190 16630 0 0 $X=68030 $Y=16470
X1399 86 M1M2_PR $T=68190 17650 0 0 $X=68030 $Y=17490
X1400 35 M1M2_PR $T=68190 24110 0 0 $X=68030 $Y=23950
X1401 86 M1M2_PR $T=68190 27850 0 0 $X=68030 $Y=27690
X1402 7 M1M2_PR $T=70950 13910 0 0 $X=70790 $Y=13750
X1403 7 M1M2_PR $T=70950 16290 0 0 $X=70790 $Y=16130
X1404 29 M1M2_PR $T=70950 31250 0 0 $X=70790 $Y=31090
X1405 39 M1M2_PR $T=73710 11530 0 0 $X=73550 $Y=11370
X1406 33 M1M2_PR $T=73710 13230 0 0 $X=73550 $Y=13070
X1407 33 M1M2_PR $T=73710 15950 0 0 $X=73550 $Y=15790
X1408 5 M1M2_PR $T=73710 16630 0 0 $X=73550 $Y=16470
X1409 41 M1M2_PR $T=73710 17650 0 0 $X=73550 $Y=17490
X1410 41 M1M2_PR $T=73710 18670 0 0 $X=73550 $Y=18510
X1411 11 M1M2_PR $T=73710 19350 0 0 $X=73550 $Y=19190
X1412 11 M1M2_PR $T=73710 25130 0 0 $X=73550 $Y=24970
X1413 5 M1M2_PR $T=73710 27170 0 0 $X=73550 $Y=27010
X1414 7 M1M2_PR $T=73710 27850 0 0 $X=73550 $Y=27690
X1415 37 M1M2_PR $T=73710 28530 0 0 $X=73550 $Y=28370
X1416 37 M1M2_PR $T=73710 29550 0 0 $X=73550 $Y=29390
X1417 7 M1M2_PR $T=73710 30230 0 0 $X=73550 $Y=30070
X1418 5 M1M2_PR $T=73710 30910 0 0 $X=73550 $Y=30750
X1419 5 M1M2_PR $T=73710 32270 0 0 $X=73550 $Y=32110
X1420 40 M1M2_PR $T=76470 16630 0 0 $X=76310 $Y=16470
X1421 39 M1M2_PR $T=76470 23090 0 0 $X=76310 $Y=22930
X1422 39 M1M2_PR $T=76470 29550 0 0 $X=76310 $Y=29390
X1423 109 M1M2_PR $T=76470 30230 0 0 $X=76310 $Y=30070
X1424 109 M1M2_PR $T=76470 31250 0 0 $X=76310 $Y=31090
X1425 109 M1M2_PR $T=76470 32610 0 0 $X=76310 $Y=32450
X1426 38 M1M2_PR $T=79230 11190 0 0 $X=79070 $Y=11030
X1427 5 M1M2_PR $T=79230 16970 0 0 $X=79070 $Y=16810
X1428 89 M1M2_PR $T=79230 17650 0 0 $X=79070 $Y=17490
X1429 89 M1M2_PR $T=79230 19010 0 0 $X=79070 $Y=18850
X1430 5 M1M2_PR $T=79230 20370 0 0 $X=79070 $Y=20210
X1431 10 M1M2_PR $T=79230 22410 0 0 $X=79070 $Y=22250
X1432 90 M1M2_PR $T=79230 24450 0 0 $X=79070 $Y=24290
X1433 90 M1M2_PR $T=79230 29550 0 0 $X=79070 $Y=29390
X1434 7 M1M2_PR $T=79230 30230 0 0 $X=79070 $Y=30070
X1435 43 M1M2_PR $T=81990 11530 0 0 $X=81830 $Y=11370
X1436 43 M1M2_PR $T=81990 16290 0 0 $X=81830 $Y=16130
X1437 41 M1M2_PR $T=81990 17650 0 0 $X=81830 $Y=17490
X1438 41 M1M2_PR $T=81990 19010 0 0 $X=81830 $Y=18850
X1439 7 M1M2_PR $T=81990 19690 0 0 $X=81830 $Y=19530
X1440 11 M1M2_PR $T=81990 23090 0 0 $X=81830 $Y=22930
X1441 5 M1M2_PR $T=81990 30910 0 0 $X=81830 $Y=30750
X1442 5 M1M2_PR $T=81990 32270 0 0 $X=81830 $Y=32110
X1443 7 M1M2_PR $T=82375 13910 0 0 $X=82215 $Y=13750
X1444 5 M1M2_PR $T=84750 16290 0 0 $X=84590 $Y=16130
X1445 35 M1M2_PR $T=84750 18670 0 0 $X=84590 $Y=18510
X1446 88 M1M2_PR $T=84750 20370 0 0 $X=84590 $Y=20210
X1447 88 M1M2_PR $T=84750 21390 0 0 $X=84590 $Y=21230
X1448 35 M1M2_PR $T=84750 24110 0 0 $X=84590 $Y=23950
X1449 91 M1M2_PR $T=84750 27510 0 0 $X=84590 $Y=27350
X1450 91 M1M2_PR $T=84750 29550 0 0 $X=84590 $Y=29390
X1451 5 M1M2_PR $T=84750 30570 0 0 $X=84590 $Y=30410
X1452 5 M1M2_PR $T=84750 32270 0 0 $X=84590 $Y=32110
X1453 44 M1M2_PR $T=86130 650 0 0 $X=85970 $Y=490
X1454 42 M1M2_PR $T=87510 10510 0 0 $X=87350 $Y=10350
X1455 43 M1M2_PR $T=87510 11870 0 0 $X=87350 $Y=11710
X1456 7 M1M2_PR $T=87510 14930 0 0 $X=87350 $Y=14770
X1457 7 M1M2_PR $T=87510 15950 0 0 $X=87350 $Y=15790
X1458 7 M1M2_PR $T=87510 16970 0 0 $X=87350 $Y=16810
X1459 43 M1M2_PR $T=87510 18670 0 0 $X=87350 $Y=18510
X1460 109 M1M2_PR $T=87510 19690 0 0 $X=87350 $Y=19530
X1461 109 M1M2_PR $T=87510 31250 0 0 $X=87350 $Y=31090
X1462 45 M1M2_PR $T=90270 11530 0 0 $X=90110 $Y=11370
X1463 45 M1M2_PR $T=90270 14590 0 0 $X=90110 $Y=14430
X1464 45 M1M2_PR $T=90270 19010 0 0 $X=90110 $Y=18850
X1465 45 M1M2_PR $T=90270 21390 0 0 $X=90110 $Y=21230
X1466 11 M1M2_PR $T=90270 22410 0 0 $X=90110 $Y=22250
X1467 11 M1M2_PR $T=90270 24790 0 0 $X=90110 $Y=24630
X1468 47 M1M2_PR $T=90270 28530 0 0 $X=90110 $Y=28370
X1469 47 M1M2_PR $T=90270 29890 0 0 $X=90110 $Y=29730
X1470 44 M1M2_PR $T=93030 650 0 0 $X=92870 $Y=490
X1471 44 M1M2_PR $T=93030 11190 0 0 $X=92870 $Y=11030
X1472 5 M1M2_PR $T=93030 13230 0 0 $X=92870 $Y=13070
X1473 5 M1M2_PR $T=93030 16630 0 0 $X=92870 $Y=16470
X1474 93 M1M2_PR $T=93030 17650 0 0 $X=92870 $Y=17490
X1475 93 M1M2_PR $T=93030 19010 0 0 $X=92870 $Y=18850
X1476 11 M1M2_PR $T=93030 19690 0 0 $X=92870 $Y=19530
X1477 11 M1M2_PR $T=93030 22410 0 0 $X=92870 $Y=22250
X1478 91 M1M2_PR $T=93030 23090 0 0 $X=92870 $Y=22930
X1479 91 M1M2_PR $T=93030 27170 0 0 $X=92870 $Y=27010
X1480 7 M1M2_PR $T=93030 27850 0 0 $X=92870 $Y=27690
X1481 7 M1M2_PR $T=93030 29890 0 0 $X=92870 $Y=29730
X1482 46 M1M2_PR $T=95790 11190 0 0 $X=95630 $Y=11030
X1483 92 M1M2_PR $T=95790 13230 0 0 $X=95630 $Y=13070
X1484 109 M1M2_PR $T=95790 13910 0 0 $X=95630 $Y=13750
X1485 109 M1M2_PR $T=95790 16970 0 0 $X=95630 $Y=16810
X1486 109 M1M2_PR $T=95790 19010 0 0 $X=95630 $Y=18850
X1487 43 M1M2_PR $T=95790 20370 0 0 $X=95630 $Y=20210
X1488 92 M1M2_PR $T=95790 24110 0 0 $X=95630 $Y=23950
X1489 43 M1M2_PR $T=95790 29550 0 0 $X=95630 $Y=29390
X1490 53 M1M2_PR $T=95790 30230 0 0 $X=95630 $Y=30070
X1491 47 M1M2_PR $T=98550 11530 0 0 $X=98390 $Y=11370
X1492 47 M1M2_PR $T=98550 13230 0 0 $X=98390 $Y=13070
X1493 47 M1M2_PR $T=98550 24110 0 0 $X=98390 $Y=23950
X1494 47 M1M2_PR $T=98550 28190 0 0 $X=98390 $Y=28030
X1495 50 M1M2_PR $T=101310 16290 0 0 $X=101150 $Y=16130
X1496 51 M1M2_PR $T=101310 16970 0 0 $X=101150 $Y=16810
X1497 51 M1M2_PR $T=101310 21390 0 0 $X=101150 $Y=21230
X1498 94 M1M2_PR $T=101310 22750 0 0 $X=101150 $Y=22590
X1499 94 M1M2_PR $T=101310 29550 0 0 $X=101150 $Y=29390
X1500 48 M1M2_PR $T=104070 14250 0 0 $X=103910 $Y=14090
X1501 7 M1M2_PR $T=104070 15950 0 0 $X=103910 $Y=15790
X1502 7 M1M2_PR $T=104070 17650 0 0 $X=103910 $Y=17490
X1503 52 M1M2_PR $T=106830 19010 0 0 $X=106670 $Y=18850
X1504 5 M1M2_PR $T=109590 15950 0 0 $X=109430 $Y=15790
X1505 7 M1M2_PR $T=109590 17650 0 0 $X=109430 $Y=17490
X1506 7 M1M2_PR $T=109590 24790 0 0 $X=109430 $Y=24630
X1507 7 M1M2_PR $T=109590 27850 0 0 $X=109430 $Y=27690
X1508 53 M1M2_PR $T=109590 29550 0 0 $X=109430 $Y=29390
X1509 49 M1M2_PR $T=112350 13910 0 0 $X=112190 $Y=13750
X1510 5 M1M2_PR $T=112350 15950 0 0 $X=112190 $Y=15790
X1511 5 M1M2_PR $T=112350 16970 0 0 $X=112190 $Y=16810
X1512 95 M1M2_PR $T=112350 17650 0 0 $X=112190 $Y=17490
X1513 95 M1M2_PR $T=112350 22750 0 0 $X=112190 $Y=22590
X1514 5 M1M2_PR $T=112350 24110 0 0 $X=112190 $Y=23950
X1515 109 M1M2_PR $T=112350 25810 0 0 $X=112190 $Y=25650
X1516 7 M1M2_PR $T=112350 27850 0 0 $X=112190 $Y=27690
X1517 7 M1M2_PR $T=112350 30230 0 0 $X=112190 $Y=30070
X1518 109 M1M2_PR $T=112350 30910 0 0 $X=112190 $Y=30750
X1519 109 M1M2_PR $T=112350 32270 0 0 $X=112190 $Y=32110
X1520 54 M1M2_PR $T=115110 14250 0 0 $X=114950 $Y=14090
X1521 49 M1M2_PR $T=115110 18670 0 0 $X=114950 $Y=18510
X1522 53 M1M2_PR $T=115110 19350 0 0 $X=114950 $Y=19190
X1523 53 M1M2_PR $T=115110 21390 0 0 $X=114950 $Y=21230
X1524 53 M1M2_PR $T=115110 29550 0 0 $X=114950 $Y=29390
X1525 55 M1M2_PR $T=117870 12210 0 0 $X=117710 $Y=12050
X1526 55 M1M2_PR $T=117870 13910 0 0 $X=117710 $Y=13750
X1527 109 M1M2_PR $T=117870 16970 0 0 $X=117710 $Y=16810
X1528 109 M1M2_PR $T=117870 19010 0 0 $X=117710 $Y=18850
X1529 12 M1M2_PR $T=117870 19690 0 0 $X=117710 $Y=19530
X1530 12 M1M2_PR $T=117870 22410 0 0 $X=117710 $Y=22250
X1531 12 M1M2_PR $T=117870 24790 0 0 $X=117710 $Y=24630
X1532 17 M1M2_PR $T=117870 25810 0 0 $X=117710 $Y=25650
X1533 17 M1M2_PR $T=117870 28190 0 0 $X=117710 $Y=28030
X1534 17 M1M2_PR $T=117870 38390 0 0 $X=117710 $Y=38230
X1535 7 M1M2_PR $T=118270 14590 0 0 $X=118110 $Y=14430
X1536 7 M1M2_PR $T=118270 16290 0 0 $X=118110 $Y=16130
X1537 96 M1M2_PR $T=120630 13230 0 0 $X=120470 $Y=13070
X1538 58 M1M2_PR $T=120630 16630 0 0 $X=120470 $Y=16470
X1539 96 M1M2_PR $T=120630 19010 0 0 $X=120470 $Y=18850
X1540 5 M1M2_PR $T=120630 27170 0 0 $X=120470 $Y=27010
X1541 5 M1M2_PR $T=120630 27850 0 0 $X=120470 $Y=27690
X1542 5 M1M2_PR $T=120630 30230 0 0 $X=120470 $Y=30070
X1543 56 M1M2_PR $T=123390 11190 0 0 $X=123230 $Y=11030
X1544 55 M1M2_PR $T=123390 12210 0 0 $X=123230 $Y=12050
X1545 55 M1M2_PR $T=123390 13570 0 0 $X=123230 $Y=13410
X1546 7 M1M2_PR $T=123390 14930 0 0 $X=123230 $Y=14770
X1547 7 M1M2_PR $T=123390 16290 0 0 $X=123230 $Y=16130
X1548 49 M1M2_PR $T=123390 17310 0 0 $X=123230 $Y=17150
X1549 49 M1M2_PR $T=123390 18670 0 0 $X=123230 $Y=18510
X1550 109 M1M2_PR $T=123390 19350 0 0 $X=123230 $Y=19190
X1551 12 M1M2_PR $T=123390 22410 0 0 $X=123230 $Y=22250
X1552 12 M1M2_PR $T=123390 27510 0 0 $X=123230 $Y=27350
X1553 109 M1M2_PR $T=123390 28190 0 0 $X=123230 $Y=28030
X1554 109 M1M2_PR $T=123390 30230 0 0 $X=123230 $Y=30070
X1555 109 M1M2_PR $T=123390 32270 0 0 $X=123230 $Y=32110
X1556 57 M1M2_PR $T=126150 11530 0 0 $X=125990 $Y=11370
X1557 57 M1M2_PR $T=126150 16290 0 0 $X=125990 $Y=16130
X1558 5 M1M2_PR $T=126150 16970 0 0 $X=125990 $Y=16810
X1559 59 M1M2_PR $T=126150 17650 0 0 $X=125990 $Y=17490
X1560 59 M1M2_PR $T=126150 21390 0 0 $X=125990 $Y=21230
X1561 98 M1M2_PR $T=126150 22750 0 0 $X=125990 $Y=22590
X1562 77 M1M2_PR $T=126150 24790 0 0 $X=125990 $Y=24630
X1563 77 M1M2_PR $T=126150 26830 0 0 $X=125990 $Y=26670
X1564 98 M1M2_PR $T=126150 29550 0 0 $X=125990 $Y=29390
X1565 5 M1M2_PR $T=126150 30570 0 0 $X=125990 $Y=30410
X1566 109 M1M2_PR $T=128910 13910 0 0 $X=128750 $Y=13750
X1567 7 M1M2_PR $T=128910 14590 0 0 $X=128750 $Y=14430
X1568 109 M1M2_PR $T=128910 16970 0 0 $X=128750 $Y=16810
X1569 7 M1M2_PR $T=128910 18670 0 0 $X=128750 $Y=18510
X1570 109 M1M2_PR $T=128910 19350 0 0 $X=128750 $Y=19190
X1571 12 M1M2_PR $T=128910 20030 0 0 $X=128750 $Y=19870
X1572 12 M1M2_PR $T=128910 22410 0 0 $X=128750 $Y=22250
X1573 109 M1M2_PR $T=128910 24110 0 0 $X=128750 $Y=23950
X1574 5 M1M2_PR $T=131670 14250 0 0 $X=131510 $Y=14090
X1575 5 M1M2_PR $T=131670 16970 0 0 $X=131510 $Y=16810
X1576 100 M1M2_PR $T=131670 17650 0 0 $X=131510 $Y=17490
X1577 100 M1M2_PR $T=131670 19010 0 0 $X=131510 $Y=18850
X1578 59 M1M2_PR $T=131670 21390 0 0 $X=131510 $Y=21230
X1579 10 M1M2_PR $T=131670 22410 0 0 $X=131510 $Y=22250
X1580 59 M1M2_PR $T=131670 25130 0 0 $X=131510 $Y=24970
X1581 75 M1M2_PR $T=131670 27850 0 0 $X=131510 $Y=27690
X1582 60 M1M2_PR $T=134430 14250 0 0 $X=134270 $Y=14090
X1583 61 M1M2_PR $T=134430 14930 0 0 $X=134270 $Y=14770
X1584 61 M1M2_PR $T=134430 16630 0 0 $X=134270 $Y=16470
X1585 61 M1M2_PR $T=134430 20370 0 0 $X=134270 $Y=20210
X1586 12 M1M2_PR $T=134430 23090 0 0 $X=134270 $Y=22930
X1587 12 M1M2_PR $T=134430 27510 0 0 $X=134270 $Y=27350
X1588 62 M1M2_PR $T=137190 11190 0 0 $X=137030 $Y=11030
X1589 55 M1M2_PR $T=137190 13570 0 0 $X=137030 $Y=13410
X1590 55 M1M2_PR $T=137190 17650 0 0 $X=137030 $Y=17490
X1591 55 M1M2_PR $T=137190 18670 0 0 $X=137030 $Y=18510
X1592 101 M1M2_PR $T=137190 22750 0 0 $X=137030 $Y=22590
X1593 101 M1M2_PR $T=137190 24110 0 0 $X=137030 $Y=23950
X1594 109 M1M2_PR $T=137190 24790 0 0 $X=137030 $Y=24630
X1595 102 M1M2_PR $T=137190 28190 0 0 $X=137030 $Y=28030
X1596 102 M1M2_PR $T=137190 29550 0 0 $X=137030 $Y=29390
X1597 109 M1M2_PR $T=137190 30230 0 0 $X=137030 $Y=30070
X1598 63 M1M2_PR $T=139950 11530 0 0 $X=139790 $Y=11370
X1599 104 M1M2_PR $T=139950 17650 0 0 $X=139790 $Y=17490
X1600 63 M1M2_PR $T=139950 23090 0 0 $X=139790 $Y=22930
X1601 63 M1M2_PR $T=139950 29890 0 0 $X=139790 $Y=29730
X1602 64 M1M2_PR $T=142710 14250 0 0 $X=142550 $Y=14090
X1603 5 M1M2_PR $T=142710 16290 0 0 $X=142550 $Y=16130
X1604 7 M1M2_PR $T=142710 16970 0 0 $X=142550 $Y=16810
X1605 109 M1M2_PR $T=142710 17650 0 0 $X=142550 $Y=17490
X1606 109 M1M2_PR $T=142710 18670 0 0 $X=142550 $Y=18510
X1607 7 M1M2_PR $T=142710 19350 0 0 $X=142550 $Y=19190
X1608 5 M1M2_PR $T=142710 20030 0 0 $X=142550 $Y=19870
X1609 7 M1M2_PR $T=142710 24790 0 0 $X=142550 $Y=24630
X1610 5 M1M2_PR $T=142710 25470 0 0 $X=142550 $Y=25310
X1611 5 M1M2_PR $T=142710 27170 0 0 $X=142550 $Y=27010
X1612 5 M1M2_PR $T=142710 29550 0 0 $X=142550 $Y=29390
X1613 5 M1M2_PR $T=142710 31250 0 0 $X=142550 $Y=31090
X1614 65 M1M2_PR $T=145470 13910 0 0 $X=145310 $Y=13750
X1615 65 M1M2_PR $T=145470 16290 0 0 $X=145310 $Y=16130
X1616 107 M1M2_PR $T=145470 17650 0 0 $X=145310 $Y=17490
X1617 107 M1M2_PR $T=145470 18670 0 0 $X=145310 $Y=18510
X1618 67 M1M2_PR $T=145470 24450 0 0 $X=145310 $Y=24290
X1619 67 M1M2_PR $T=145470 26830 0 0 $X=145310 $Y=26670
X1620 69 M1M2_PR $T=148230 11530 0 0 $X=148070 $Y=11370
X1621 103 M1M2_PR $T=148230 17650 0 0 $X=148070 $Y=17490
X1622 103 M1M2_PR $T=148230 19010 0 0 $X=148070 $Y=18850
X1623 69 M1M2_PR $T=148230 19690 0 0 $X=148070 $Y=19530
X1624 109 M1M2_PR $T=148230 22410 0 0 $X=148070 $Y=22250
X1625 109 M1M2_PR $T=148230 24110 0 0 $X=148070 $Y=23950
X1626 104 M1M2_PR $T=150990 16630 0 0 $X=150830 $Y=16470
X1627 66 M1M2_PR $T=150990 25130 0 0 $X=150830 $Y=24970
X1628 7 M1M2_PR $T=150990 25810 0 0 $X=150830 $Y=25650
X1629 7 M1M2_PR $T=150990 27850 0 0 $X=150830 $Y=27690
X1630 7 M1M2_PR $T=150990 29890 0 0 $X=150830 $Y=29730
X1631 68 M1M2_PR $T=153750 11190 0 0 $X=153590 $Y=11030
X1632 13 M1M2_PR $T=153750 16970 0 0 $X=153590 $Y=16810
X1633 13 M1M2_PR $T=153750 19350 0 0 $X=153590 $Y=19190
X1634 13 M1M2_PR $T=153750 22070 0 0 $X=153590 $Y=21910
X1635 105 M1M2_PR $T=153750 22750 0 0 $X=153590 $Y=22590
X1636 105 M1M2_PR $T=153750 24110 0 0 $X=153590 $Y=23950
X1637 5 M1M2_PR $T=153750 25470 0 0 $X=153590 $Y=25310
X1638 5 M1M2_PR $T=153750 26830 0 0 $X=153590 $Y=26670
X1639 71 M1M2_PR $T=156510 16970 0 0 $X=156350 $Y=16810
X1640 71 M1M2_PR $T=156510 23090 0 0 $X=156350 $Y=22930
X1641 71 M1M2_PR $T=156510 28190 0 0 $X=156350 $Y=28030
X1642 71 M1M2_PR $T=156510 30230 0 0 $X=156350 $Y=30070
X1643 109 M1M2_PR $T=159270 13910 0 0 $X=159110 $Y=13750
X1644 109 M1M2_PR $T=159270 22410 0 0 $X=159110 $Y=22250
X1645 109 M1M2_PR $T=159270 27850 0 0 $X=159110 $Y=27690
X1646 72 M1M2_PR $T=162030 11190 0 0 $X=161870 $Y=11030
X1647 13 M1M2_PR $T=162030 22410 0 0 $X=161870 $Y=22250
X1648 106 M1M2_PR $T=162030 23090 0 0 $X=161870 $Y=22930
X1649 106 M1M2_PR $T=162030 26830 0 0 $X=161870 $Y=26670
X1650 70 M1M2_PR $T=164790 16630 0 0 $X=164630 $Y=16470
X1651 13 M1M2_PR $T=164790 19350 0 0 $X=164630 $Y=19190
X1652 75 M1M2_PR $T=164790 23090 0 0 $X=164630 $Y=22930
X1653 75 M1M2_PR $T=164790 24110 0 0 $X=164630 $Y=23950
X1654 73 M1M2_PR $T=167550 12210 0 0 $X=167390 $Y=12050
X1655 73 M1M2_PR $T=167550 13570 0 0 $X=167390 $Y=13410
X1656 4 M1M2_PR $T=167550 14930 0 0 $X=167390 $Y=14770
X1657 4 M1M2_PR $T=167550 18670 0 0 $X=167390 $Y=18510
X1658 7 M1M2_PR $T=167550 20370 0 0 $X=167390 $Y=20210
X1659 7 M1M2_PR $T=167550 24450 0 0 $X=167390 $Y=24290
X1660 5 M1M2_PR $T=167550 25470 0 0 $X=167390 $Y=25310
X1661 5 M1M2_PR $T=167550 26830 0 0 $X=167390 $Y=26670
X1662 6 M1M2_PR $T=170310 13910 0 0 $X=170150 $Y=13750
X1663 13 M1M2_PR $T=170310 17310 0 0 $X=170150 $Y=17150
X1664 13 M1M2_PR $T=170310 21730 0 0 $X=170150 $Y=21570
X1665 10 M1M2_PR $T=170310 22410 0 0 $X=170150 $Y=22250
X1666 6 M1M2_PR $T=170310 23090 0 0 $X=170150 $Y=22930
X1667 6 M1M2_PR $T=170310 32950 0 0 $X=170150 $Y=32790
X1668 69 M1M2_PR $T=173070 10510 0 0 $X=172910 $Y=10350
X1669 8 M1M2_PR $T=173070 13910 0 0 $X=172910 $Y=13750
X1670 8 M1M2_PR $T=173070 19350 0 0 $X=172910 $Y=19190
X1671 69 M1M2_PR $T=173070 20030 0 0 $X=172910 $Y=19870
X1672 5 M1M2_PR $T=173070 22750 0 0 $X=172910 $Y=22590
X1673 69 M1M2_PR $T=173070 24110 0 0 $X=172910 $Y=23950
X1674 5 M1M2_PR $T=173070 24790 0 0 $X=172910 $Y=24630
X1675 8 M1M2_PR $T=173530 9490 0 0 $X=173370 $Y=9330
X1676 65 M1M2_PR $T=175830 14590 0 0 $X=175670 $Y=14430
X1677 65 M1M2_PR $T=175830 15950 0 0 $X=175670 $Y=15790
X1678 75 M1M2_PR $T=175830 16970 0 0 $X=175670 $Y=16810
X1679 75 M1M2_PR $T=175830 21390 0 0 $X=175670 $Y=21230
X1680 108 M1M2_PR $T=175830 22750 0 0 $X=175670 $Y=22590
X1681 108 M1M2_PR $T=175830 24110 0 0 $X=175670 $Y=23950
X1682 74 M1M2_PR $T=178590 16630 0 0 $X=178430 $Y=16470
X1683 8 M1M2_PR $T=180430 9490 0 0 $X=180270 $Y=9330
X1684 77 M1M2_PR $T=181350 24790 0 0 $X=181190 $Y=24630
X1685 77 M1M2_PR $T=181350 28190 0 0 $X=181190 $Y=28030
X1686 73 M1M2_PR $T=184110 13570 0 0 $X=183950 $Y=13410
X1687 73 M1M2_PR $T=184110 21390 0 0 $X=183950 $Y=21230
X1688 76 M1M2_PR $T=186870 24450 0 0 $X=186710 $Y=24290
X1689 14 M2M3_PR $T=15750 1630 0 0 $X=15585 $Y=1445
X1690 20 M2M3_PR $T=26790 1020 0 0 $X=26625 $Y=835
X1691 24 M2M3_PR $T=35070 1020 0 0 $X=34905 $Y=835
X1692 7 M2M3_PR $T=43350 15050 0 0 $X=43185 $Y=14865
X1693 25 M2M3_PR $T=46570 8950 0 0 $X=46405 $Y=8765
X1694 30 M2M3_PR $T=48870 10170 0 0 $X=48705 $Y=9985
X1695 9 M2M3_PR $T=48870 22980 0 0 $X=48705 $Y=22795
X1696 7 M2M3_PR $T=51630 14440 0 0 $X=51465 $Y=14255
X1697 109 M2M3_PR $T=54390 27250 0 0 $X=54225 $Y=27065
X1698 5 M2M3_PR $T=59910 15050 0 0 $X=59745 $Y=14865
X1699 9 M2M3_PR $T=59910 22980 0 0 $X=59745 $Y=22795
X1700 25 M2M3_PR $T=62670 13830 0 0 $X=62505 $Y=13645
X1701 32 M2M3_PR $T=65430 1020 0 0 $X=65265 $Y=835
X1702 11 M2M3_PR $T=65430 26030 0 0 $X=65265 $Y=25845
X1703 109 M2M3_PR $T=65430 27250 0 0 $X=65265 $Y=27065
X1704 39 M2M3_PR $T=73710 10780 0 0 $X=73545 $Y=10595
X1705 11 M2M3_PR $T=73710 26030 0 0 $X=73545 $Y=25845
X1706 7 M2M3_PR $T=73710 30300 0 0 $X=73545 $Y=30115
X1707 40 M2M3_PR $T=76470 3460 0 0 $X=76305 $Y=3275
X1708 39 M2M3_PR $T=76470 18100 0 0 $X=76305 $Y=17915
X1709 5 M2M3_PR $T=79230 15050 0 0 $X=79065 $Y=14865
X1710 10 M2M3_PR $T=79230 22370 0 0 $X=79065 $Y=22185
X1711 7 M2M3_PR $T=79230 30300 0 0 $X=79065 $Y=30115
X1712 11 M2M3_PR $T=81990 26030 0 0 $X=81825 $Y=25845
X1713 5 M2M3_PR $T=84750 15050 0 0 $X=84585 $Y=14865
X1714 42 M2M3_PR $T=87510 10170 0 0 $X=87345 $Y=9985
X1715 5 M2M3_PR $T=93030 15050 0 0 $X=92865 $Y=14865
X1716 7 M2M3_PR $T=93030 30910 0 0 $X=92865 $Y=30725
X1717 53 M2M3_PR $T=95790 30300 0 0 $X=95625 $Y=30115
X1718 50 M2M3_PR $T=101310 2850 0 0 $X=101145 $Y=2665
X1719 52 M2M3_PR $T=107290 8950 0 0 $X=107125 $Y=8765
X1720 5 M2M3_PR $T=109590 15050 0 0 $X=109425 $Y=14865
X1721 53 M2M3_PR $T=109590 30300 0 0 $X=109425 $Y=30115
X1722 49 M2M3_PR $T=112350 15050 0 0 $X=112185 $Y=14865
X1723 49 M2M3_PR $T=115110 15050 0 0 $X=114945 $Y=14865
X1724 58 M2M3_PR $T=120630 14440 0 0 $X=120465 $Y=14255
X1725 109 M2M3_PR $T=128910 18100 0 0 $X=128745 $Y=17915
X1726 5 M2M3_PR $T=131670 15050 0 0 $X=131505 $Y=14865
X1727 10 M2M3_PR $T=131670 22370 0 0 $X=131505 $Y=22185
X1728 75 M2M3_PR $T=131670 26030 0 0 $X=131505 $Y=25845
X1729 62 M2M3_PR $T=137190 1020 0 0 $X=137025 $Y=835
X1730 104 M2M3_PR $T=140410 9560 0 0 $X=140245 $Y=9375
X1731 5 M2M3_PR $T=142710 15050 0 0 $X=142545 $Y=14865
X1732 109 M2M3_PR $T=142710 18710 0 0 $X=142545 $Y=18525
X1733 104 M2M3_PR $T=150530 9560 0 0 $X=150365 $Y=9375
X1734 66 M2M3_PR $T=151450 8950 0 0 $X=151285 $Y=8765
X1735 13 M2M3_PR $T=153750 18710 0 0 $X=153585 $Y=18525
X1736 13 M2M3_PR $T=162030 18710 0 0 $X=161865 $Y=18525
X1737 70 M2M3_PR $T=164790 3460 0 0 $X=164625 $Y=3275
X1738 13 M2M3_PR $T=164790 18710 0 0 $X=164625 $Y=18525
X1739 75 M2M3_PR $T=164790 26030 0 0 $X=164625 $Y=25845
X1740 13 M2M3_PR $T=170310 18710 0 0 $X=170145 $Y=18525
X1741 10 M2M3_PR $T=170310 22370 0 0 $X=170145 $Y=22185
X1742 74 M2M3_PR $T=178590 4070 0 0 $X=178425 $Y=3885
X1743 76 M2M3_PR $T=186870 5290 0 0 $X=186705 $Y=5105
X1744 10 M2M3_PR $T=189630 1020 0 0 $X=189465 $Y=835
X1745 14 M3M4_PR $T=10230 1630 0 0 $X=10040 $Y=1465
X1746 20 M3M4_PR $T=23340 1020 0 0 $X=23150 $Y=855
X1747 24 M3M4_PR $T=36450 1020 0 0 $X=36260 $Y=855
X1748 30 M3M4_PR $T=48870 10170 0 0 $X=48680 $Y=10005
X1749 25 M3M4_PR $T=60600 8950 0 0 $X=60410 $Y=8785
X1750 25 M3M4_PR $T=60600 13830 0 0 $X=60410 $Y=13665
X1751 32 M3M4_PR $T=61980 1020 0 0 $X=61790 $Y=855
X1752 40 M3M4_PR $T=74400 3460 0 0 $X=74210 $Y=3295
X1753 39 M3M4_PR $T=76470 10780 0 0 $X=76280 $Y=10615
X1754 39 M3M4_PR $T=76470 18100 0 0 $X=76280 $Y=17935
X1755 42 M3M4_PR $T=87510 10170 0 0 $X=87320 $Y=10005
X1756 50 M3M4_PR $T=99930 2850 0 0 $X=99740 $Y=2685
X1757 52 M3M4_PR $T=113040 8950 0 0 $X=112850 $Y=8785
X1758 58 M3M4_PR $T=126150 14440 0 0 $X=125960 $Y=14275
X1759 62 M3M4_PR $T=138570 1020 0 0 $X=138380 $Y=855
X1760 66 M3M4_PR $T=151680 8950 0 0 $X=151490 $Y=8785
X1761 70 M3M4_PR $T=164100 3460 0 0 $X=163910 $Y=3295
X1762 10 M3M4_PR $T=171000 1020 0 0 $X=170810 $Y=855
X1763 10 M3M4_PR $T=171000 22370 0 0 $X=170810 $Y=22205
X1764 74 M3M4_PR $T=177210 4070 0 0 $X=177020 $Y=3905
X1765 76 M3M4_PR $T=189630 5290 0 0 $X=189440 $Y=5125
X1766 3 DigitalLDOLogic_VIA0 $T=11150 12720 0 0 $X=10900 $Y=12480
X1767 3 DigitalLDOLogic_VIA0 $T=11150 18160 0 0 $X=10900 $Y=17920
X1768 3 DigitalLDOLogic_VIA0 $T=11150 23600 0 0 $X=10900 $Y=23360
X1769 3 DigitalLDOLogic_VIA0 $T=11150 29040 0 0 $X=10900 $Y=28800
X1770 3 DigitalLDOLogic_VIA0 $T=11150 34480 0 0 $X=10900 $Y=34240
X1771 3 DigitalLDOLogic_VIA0 $T=11150 39920 0 0 $X=10900 $Y=39680
X1772 3 DigitalLDOLogic_VIA0 $T=11150 45360 0 0 $X=10900 $Y=45120
X1773 3 DigitalLDOLogic_VIA0 $T=11150 50800 0 0 $X=10900 $Y=50560
X1774 3 DigitalLDOLogic_VIA0 $T=11150 56240 0 0 $X=10900 $Y=56000
X1775 1 DigitalLDOLogic_VIA0 $T=12070 15440 0 0 $X=11820 $Y=15200
X1776 1 DigitalLDOLogic_VIA0 $T=12070 20880 0 0 $X=11820 $Y=20640
X1777 1 DigitalLDOLogic_VIA0 $T=12070 26320 0 0 $X=11820 $Y=26080
X1778 1 DigitalLDOLogic_VIA0 $T=12070 31760 0 0 $X=11820 $Y=31520
X1779 1 DigitalLDOLogic_VIA0 $T=12070 37200 0 0 $X=11820 $Y=36960
X1780 1 DigitalLDOLogic_VIA0 $T=12070 42640 0 0 $X=11820 $Y=42400
X1781 1 DigitalLDOLogic_VIA0 $T=12070 48080 0 0 $X=11820 $Y=47840
X1782 1 DigitalLDOLogic_VIA0 $T=12070 53520 0 0 $X=11820 $Y=53280
X1783 1 DigitalLDOLogic_VIA0 $T=12070 58960 0 0 $X=11820 $Y=58720
X1784 3 DigitalLDOLogic_VIA0 $T=13910 12720 0 0 $X=13660 $Y=12480
X1785 3 DigitalLDOLogic_VIA0 $T=13910 18160 0 0 $X=13660 $Y=17920
X1786 3 DigitalLDOLogic_VIA0 $T=13910 23600 0 0 $X=13660 $Y=23360
X1787 3 DigitalLDOLogic_VIA0 $T=13910 29040 0 0 $X=13660 $Y=28800
X1788 3 DigitalLDOLogic_VIA0 $T=13910 34480 0 0 $X=13660 $Y=34240
X1789 3 DigitalLDOLogic_VIA0 $T=13910 39920 0 0 $X=13660 $Y=39680
X1790 3 DigitalLDOLogic_VIA0 $T=13910 45360 0 0 $X=13660 $Y=45120
X1791 3 DigitalLDOLogic_VIA0 $T=13910 50800 0 0 $X=13660 $Y=50560
X1792 3 DigitalLDOLogic_VIA0 $T=13910 56240 0 0 $X=13660 $Y=56000
X1793 1 DigitalLDOLogic_VIA0 $T=14830 15440 0 0 $X=14580 $Y=15200
X1794 1 DigitalLDOLogic_VIA0 $T=14830 20880 0 0 $X=14580 $Y=20640
X1795 1 DigitalLDOLogic_VIA0 $T=14830 26320 0 0 $X=14580 $Y=26080
X1796 1 DigitalLDOLogic_VIA0 $T=14830 31760 0 0 $X=14580 $Y=31520
X1797 1 DigitalLDOLogic_VIA0 $T=14830 37200 0 0 $X=14580 $Y=36960
X1798 1 DigitalLDOLogic_VIA0 $T=14830 42640 0 0 $X=14580 $Y=42400
X1799 1 DigitalLDOLogic_VIA0 $T=14830 48080 0 0 $X=14580 $Y=47840
X1800 1 DigitalLDOLogic_VIA0 $T=14830 53520 0 0 $X=14580 $Y=53280
X1801 1 DigitalLDOLogic_VIA0 $T=14830 58960 0 0 $X=14580 $Y=58720
X1802 3 DigitalLDOLogic_VIA0 $T=16670 12720 0 0 $X=16420 $Y=12480
X1803 3 DigitalLDOLogic_VIA0 $T=16670 18160 0 0 $X=16420 $Y=17920
X1804 3 DigitalLDOLogic_VIA0 $T=16670 23600 0 0 $X=16420 $Y=23360
X1805 3 DigitalLDOLogic_VIA0 $T=16670 29040 0 0 $X=16420 $Y=28800
X1806 3 DigitalLDOLogic_VIA0 $T=16670 34480 0 0 $X=16420 $Y=34240
X1807 3 DigitalLDOLogic_VIA0 $T=16670 39920 0 0 $X=16420 $Y=39680
X1808 3 DigitalLDOLogic_VIA0 $T=16670 45360 0 0 $X=16420 $Y=45120
X1809 3 DigitalLDOLogic_VIA0 $T=16670 50800 0 0 $X=16420 $Y=50560
X1810 3 DigitalLDOLogic_VIA0 $T=16670 56240 0 0 $X=16420 $Y=56000
X1811 1 DigitalLDOLogic_VIA0 $T=17590 15440 0 0 $X=17340 $Y=15200
X1812 1 DigitalLDOLogic_VIA0 $T=17590 20880 0 0 $X=17340 $Y=20640
X1813 1 DigitalLDOLogic_VIA0 $T=17590 26320 0 0 $X=17340 $Y=26080
X1814 1 DigitalLDOLogic_VIA0 $T=17590 31760 0 0 $X=17340 $Y=31520
X1815 1 DigitalLDOLogic_VIA0 $T=17590 37200 0 0 $X=17340 $Y=36960
X1816 1 DigitalLDOLogic_VIA0 $T=17590 42640 0 0 $X=17340 $Y=42400
X1817 1 DigitalLDOLogic_VIA0 $T=17590 48080 0 0 $X=17340 $Y=47840
X1818 1 DigitalLDOLogic_VIA0 $T=17590 53520 0 0 $X=17340 $Y=53280
X1819 1 DigitalLDOLogic_VIA0 $T=17590 58960 0 0 $X=17340 $Y=58720
X1820 3 DigitalLDOLogic_VIA0 $T=19430 12720 0 0 $X=19180 $Y=12480
X1821 3 DigitalLDOLogic_VIA0 $T=19430 18160 0 0 $X=19180 $Y=17920
X1822 3 DigitalLDOLogic_VIA0 $T=19430 23600 0 0 $X=19180 $Y=23360
X1823 3 DigitalLDOLogic_VIA0 $T=19430 29040 0 0 $X=19180 $Y=28800
X1824 3 DigitalLDOLogic_VIA0 $T=19430 34480 0 0 $X=19180 $Y=34240
X1825 3 DigitalLDOLogic_VIA0 $T=19430 39920 0 0 $X=19180 $Y=39680
X1826 3 DigitalLDOLogic_VIA0 $T=19430 45360 0 0 $X=19180 $Y=45120
X1827 3 DigitalLDOLogic_VIA0 $T=19430 50800 0 0 $X=19180 $Y=50560
X1828 3 DigitalLDOLogic_VIA0 $T=19430 56240 0 0 $X=19180 $Y=56000
X1829 1 DigitalLDOLogic_VIA0 $T=20350 15440 0 0 $X=20100 $Y=15200
X1830 1 DigitalLDOLogic_VIA0 $T=20350 20880 0 0 $X=20100 $Y=20640
X1831 1 DigitalLDOLogic_VIA0 $T=20350 26320 0 0 $X=20100 $Y=26080
X1832 1 DigitalLDOLogic_VIA0 $T=20350 31760 0 0 $X=20100 $Y=31520
X1833 1 DigitalLDOLogic_VIA0 $T=20350 37200 0 0 $X=20100 $Y=36960
X1834 1 DigitalLDOLogic_VIA0 $T=20350 42640 0 0 $X=20100 $Y=42400
X1835 1 DigitalLDOLogic_VIA0 $T=20350 48080 0 0 $X=20100 $Y=47840
X1836 1 DigitalLDOLogic_VIA0 $T=20350 53520 0 0 $X=20100 $Y=53280
X1837 1 DigitalLDOLogic_VIA0 $T=20350 58960 0 0 $X=20100 $Y=58720
X1838 3 DigitalLDOLogic_VIA0 $T=22190 12720 0 0 $X=21940 $Y=12480
X1839 3 DigitalLDOLogic_VIA0 $T=22190 18160 0 0 $X=21940 $Y=17920
X1840 3 DigitalLDOLogic_VIA0 $T=22190 23600 0 0 $X=21940 $Y=23360
X1841 3 DigitalLDOLogic_VIA0 $T=22190 29040 0 0 $X=21940 $Y=28800
X1842 3 DigitalLDOLogic_VIA0 $T=22190 34480 0 0 $X=21940 $Y=34240
X1843 3 DigitalLDOLogic_VIA0 $T=22190 39920 0 0 $X=21940 $Y=39680
X1844 3 DigitalLDOLogic_VIA0 $T=22190 45360 0 0 $X=21940 $Y=45120
X1845 3 DigitalLDOLogic_VIA0 $T=22190 50800 0 0 $X=21940 $Y=50560
X1846 3 DigitalLDOLogic_VIA0 $T=22190 56240 0 0 $X=21940 $Y=56000
X1847 1 DigitalLDOLogic_VIA0 $T=23110 15440 0 0 $X=22860 $Y=15200
X1848 1 DigitalLDOLogic_VIA0 $T=23110 20880 0 0 $X=22860 $Y=20640
X1849 1 DigitalLDOLogic_VIA0 $T=23110 26320 0 0 $X=22860 $Y=26080
X1850 1 DigitalLDOLogic_VIA0 $T=23110 31760 0 0 $X=22860 $Y=31520
X1851 1 DigitalLDOLogic_VIA0 $T=23110 37200 0 0 $X=22860 $Y=36960
X1852 1 DigitalLDOLogic_VIA0 $T=23110 42640 0 0 $X=22860 $Y=42400
X1853 1 DigitalLDOLogic_VIA0 $T=23110 48080 0 0 $X=22860 $Y=47840
X1854 1 DigitalLDOLogic_VIA0 $T=23110 53520 0 0 $X=22860 $Y=53280
X1855 1 DigitalLDOLogic_VIA0 $T=23110 58960 0 0 $X=22860 $Y=58720
X1856 3 DigitalLDOLogic_VIA0 $T=24950 12720 0 0 $X=24700 $Y=12480
X1857 3 DigitalLDOLogic_VIA0 $T=24950 18160 0 0 $X=24700 $Y=17920
X1858 3 DigitalLDOLogic_VIA0 $T=24950 23600 0 0 $X=24700 $Y=23360
X1859 3 DigitalLDOLogic_VIA0 $T=24950 29040 0 0 $X=24700 $Y=28800
X1860 3 DigitalLDOLogic_VIA0 $T=24950 34480 0 0 $X=24700 $Y=34240
X1861 3 DigitalLDOLogic_VIA0 $T=24950 39920 0 0 $X=24700 $Y=39680
X1862 3 DigitalLDOLogic_VIA0 $T=24950 45360 0 0 $X=24700 $Y=45120
X1863 3 DigitalLDOLogic_VIA0 $T=24950 50800 0 0 $X=24700 $Y=50560
X1864 3 DigitalLDOLogic_VIA0 $T=24950 56240 0 0 $X=24700 $Y=56000
X1865 1 DigitalLDOLogic_VIA0 $T=25870 15440 0 0 $X=25620 $Y=15200
X1866 1 DigitalLDOLogic_VIA0 $T=25870 20880 0 0 $X=25620 $Y=20640
X1867 1 DigitalLDOLogic_VIA0 $T=25870 26320 0 0 $X=25620 $Y=26080
X1868 1 DigitalLDOLogic_VIA0 $T=25870 31760 0 0 $X=25620 $Y=31520
X1869 1 DigitalLDOLogic_VIA0 $T=25870 37200 0 0 $X=25620 $Y=36960
X1870 1 DigitalLDOLogic_VIA0 $T=25870 42640 0 0 $X=25620 $Y=42400
X1871 1 DigitalLDOLogic_VIA0 $T=25870 48080 0 0 $X=25620 $Y=47840
X1872 1 DigitalLDOLogic_VIA0 $T=25870 53520 0 0 $X=25620 $Y=53280
X1873 1 DigitalLDOLogic_VIA0 $T=25870 58960 0 0 $X=25620 $Y=58720
X1874 3 DigitalLDOLogic_VIA0 $T=27710 12720 0 0 $X=27460 $Y=12480
X1875 3 DigitalLDOLogic_VIA0 $T=27710 18160 0 0 $X=27460 $Y=17920
X1876 3 DigitalLDOLogic_VIA0 $T=27710 23600 0 0 $X=27460 $Y=23360
X1877 3 DigitalLDOLogic_VIA0 $T=27710 29040 0 0 $X=27460 $Y=28800
X1878 3 DigitalLDOLogic_VIA0 $T=27710 34480 0 0 $X=27460 $Y=34240
X1879 3 DigitalLDOLogic_VIA0 $T=27710 39920 0 0 $X=27460 $Y=39680
X1880 3 DigitalLDOLogic_VIA0 $T=27710 45360 0 0 $X=27460 $Y=45120
X1881 3 DigitalLDOLogic_VIA0 $T=27710 50800 0 0 $X=27460 $Y=50560
X1882 3 DigitalLDOLogic_VIA0 $T=27710 56240 0 0 $X=27460 $Y=56000
X1883 1 DigitalLDOLogic_VIA0 $T=28630 15440 0 0 $X=28380 $Y=15200
X1884 1 DigitalLDOLogic_VIA0 $T=28630 20880 0 0 $X=28380 $Y=20640
X1885 1 DigitalLDOLogic_VIA0 $T=28630 26320 0 0 $X=28380 $Y=26080
X1886 1 DigitalLDOLogic_VIA0 $T=28630 31760 0 0 $X=28380 $Y=31520
X1887 1 DigitalLDOLogic_VIA0 $T=28630 37200 0 0 $X=28380 $Y=36960
X1888 1 DigitalLDOLogic_VIA0 $T=28630 42640 0 0 $X=28380 $Y=42400
X1889 1 DigitalLDOLogic_VIA0 $T=28630 48080 0 0 $X=28380 $Y=47840
X1890 1 DigitalLDOLogic_VIA0 $T=28630 53520 0 0 $X=28380 $Y=53280
X1891 1 DigitalLDOLogic_VIA0 $T=28630 58960 0 0 $X=28380 $Y=58720
X1892 3 DigitalLDOLogic_VIA0 $T=30470 12720 0 0 $X=30220 $Y=12480
X1893 3 DigitalLDOLogic_VIA0 $T=30470 18160 0 0 $X=30220 $Y=17920
X1894 3 DigitalLDOLogic_VIA0 $T=30470 23600 0 0 $X=30220 $Y=23360
X1895 3 DigitalLDOLogic_VIA0 $T=30470 29040 0 0 $X=30220 $Y=28800
X1896 3 DigitalLDOLogic_VIA0 $T=30470 34480 0 0 $X=30220 $Y=34240
X1897 3 DigitalLDOLogic_VIA0 $T=30470 39920 0 0 $X=30220 $Y=39680
X1898 3 DigitalLDOLogic_VIA0 $T=30470 45360 0 0 $X=30220 $Y=45120
X1899 3 DigitalLDOLogic_VIA0 $T=30470 50800 0 0 $X=30220 $Y=50560
X1900 3 DigitalLDOLogic_VIA0 $T=30470 56240 0 0 $X=30220 $Y=56000
X1901 1 DigitalLDOLogic_VIA0 $T=31390 15440 0 0 $X=31140 $Y=15200
X1902 1 DigitalLDOLogic_VIA0 $T=31390 20880 0 0 $X=31140 $Y=20640
X1903 1 DigitalLDOLogic_VIA0 $T=31390 26320 0 0 $X=31140 $Y=26080
X1904 1 DigitalLDOLogic_VIA0 $T=31390 31760 0 0 $X=31140 $Y=31520
X1905 1 DigitalLDOLogic_VIA0 $T=31390 37200 0 0 $X=31140 $Y=36960
X1906 1 DigitalLDOLogic_VIA0 $T=31390 42640 0 0 $X=31140 $Y=42400
X1907 1 DigitalLDOLogic_VIA0 $T=31390 48080 0 0 $X=31140 $Y=47840
X1908 1 DigitalLDOLogic_VIA0 $T=31390 53520 0 0 $X=31140 $Y=53280
X1909 1 DigitalLDOLogic_VIA0 $T=31390 58960 0 0 $X=31140 $Y=58720
X1910 3 DigitalLDOLogic_VIA0 $T=33230 12720 0 0 $X=32980 $Y=12480
X1911 3 DigitalLDOLogic_VIA0 $T=33230 18160 0 0 $X=32980 $Y=17920
X1912 3 DigitalLDOLogic_VIA0 $T=33230 23600 0 0 $X=32980 $Y=23360
X1913 3 DigitalLDOLogic_VIA0 $T=33230 29040 0 0 $X=32980 $Y=28800
X1914 3 DigitalLDOLogic_VIA0 $T=33230 34480 0 0 $X=32980 $Y=34240
X1915 3 DigitalLDOLogic_VIA0 $T=33230 39920 0 0 $X=32980 $Y=39680
X1916 3 DigitalLDOLogic_VIA0 $T=33230 45360 0 0 $X=32980 $Y=45120
X1917 3 DigitalLDOLogic_VIA0 $T=33230 50800 0 0 $X=32980 $Y=50560
X1918 3 DigitalLDOLogic_VIA0 $T=33230 56240 0 0 $X=32980 $Y=56000
X1919 1 DigitalLDOLogic_VIA0 $T=34150 15440 0 0 $X=33900 $Y=15200
X1920 1 DigitalLDOLogic_VIA0 $T=34150 20880 0 0 $X=33900 $Y=20640
X1921 1 DigitalLDOLogic_VIA0 $T=34150 26320 0 0 $X=33900 $Y=26080
X1922 1 DigitalLDOLogic_VIA0 $T=34150 31760 0 0 $X=33900 $Y=31520
X1923 1 DigitalLDOLogic_VIA0 $T=34150 37200 0 0 $X=33900 $Y=36960
X1924 1 DigitalLDOLogic_VIA0 $T=34150 42640 0 0 $X=33900 $Y=42400
X1925 1 DigitalLDOLogic_VIA0 $T=34150 48080 0 0 $X=33900 $Y=47840
X1926 1 DigitalLDOLogic_VIA0 $T=34150 53520 0 0 $X=33900 $Y=53280
X1927 1 DigitalLDOLogic_VIA0 $T=34150 58960 0 0 $X=33900 $Y=58720
X1928 3 DigitalLDOLogic_VIA0 $T=35990 12720 0 0 $X=35740 $Y=12480
X1929 3 DigitalLDOLogic_VIA0 $T=35990 18160 0 0 $X=35740 $Y=17920
X1930 3 DigitalLDOLogic_VIA0 $T=35990 23600 0 0 $X=35740 $Y=23360
X1931 3 DigitalLDOLogic_VIA0 $T=35990 29040 0 0 $X=35740 $Y=28800
X1932 3 DigitalLDOLogic_VIA0 $T=35990 34480 0 0 $X=35740 $Y=34240
X1933 3 DigitalLDOLogic_VIA0 $T=35990 39920 0 0 $X=35740 $Y=39680
X1934 3 DigitalLDOLogic_VIA0 $T=35990 45360 0 0 $X=35740 $Y=45120
X1935 3 DigitalLDOLogic_VIA0 $T=35990 50800 0 0 $X=35740 $Y=50560
X1936 3 DigitalLDOLogic_VIA0 $T=35990 56240 0 0 $X=35740 $Y=56000
X1937 1 DigitalLDOLogic_VIA0 $T=36910 15440 0 0 $X=36660 $Y=15200
X1938 1 DigitalLDOLogic_VIA0 $T=36910 20880 0 0 $X=36660 $Y=20640
X1939 1 DigitalLDOLogic_VIA0 $T=36910 26320 0 0 $X=36660 $Y=26080
X1940 1 DigitalLDOLogic_VIA0 $T=36910 31760 0 0 $X=36660 $Y=31520
X1941 1 DigitalLDOLogic_VIA0 $T=36910 37200 0 0 $X=36660 $Y=36960
X1942 1 DigitalLDOLogic_VIA0 $T=36910 42640 0 0 $X=36660 $Y=42400
X1943 1 DigitalLDOLogic_VIA0 $T=36910 48080 0 0 $X=36660 $Y=47840
X1944 1 DigitalLDOLogic_VIA0 $T=36910 53520 0 0 $X=36660 $Y=53280
X1945 1 DigitalLDOLogic_VIA0 $T=36910 58960 0 0 $X=36660 $Y=58720
X1946 3 DigitalLDOLogic_VIA0 $T=38750 12720 0 0 $X=38500 $Y=12480
X1947 3 DigitalLDOLogic_VIA0 $T=38750 18160 0 0 $X=38500 $Y=17920
X1948 3 DigitalLDOLogic_VIA0 $T=38750 23600 0 0 $X=38500 $Y=23360
X1949 3 DigitalLDOLogic_VIA0 $T=38750 29040 0 0 $X=38500 $Y=28800
X1950 3 DigitalLDOLogic_VIA0 $T=38750 34480 0 0 $X=38500 $Y=34240
X1951 3 DigitalLDOLogic_VIA0 $T=38750 39920 0 0 $X=38500 $Y=39680
X1952 3 DigitalLDOLogic_VIA0 $T=38750 45360 0 0 $X=38500 $Y=45120
X1953 3 DigitalLDOLogic_VIA0 $T=38750 50800 0 0 $X=38500 $Y=50560
X1954 3 DigitalLDOLogic_VIA0 $T=38750 56240 0 0 $X=38500 $Y=56000
X1955 1 DigitalLDOLogic_VIA0 $T=39670 15440 0 0 $X=39420 $Y=15200
X1956 1 DigitalLDOLogic_VIA0 $T=39670 20880 0 0 $X=39420 $Y=20640
X1957 1 DigitalLDOLogic_VIA0 $T=39670 26320 0 0 $X=39420 $Y=26080
X1958 1 DigitalLDOLogic_VIA0 $T=39670 31760 0 0 $X=39420 $Y=31520
X1959 1 DigitalLDOLogic_VIA0 $T=39670 37200 0 0 $X=39420 $Y=36960
X1960 1 DigitalLDOLogic_VIA0 $T=39670 42640 0 0 $X=39420 $Y=42400
X1961 1 DigitalLDOLogic_VIA0 $T=39670 48080 0 0 $X=39420 $Y=47840
X1962 1 DigitalLDOLogic_VIA0 $T=39670 53520 0 0 $X=39420 $Y=53280
X1963 1 DigitalLDOLogic_VIA0 $T=39670 58960 0 0 $X=39420 $Y=58720
X1964 3 DigitalLDOLogic_VIA0 $T=41510 12720 0 0 $X=41260 $Y=12480
X1965 3 DigitalLDOLogic_VIA0 $T=41510 18160 0 0 $X=41260 $Y=17920
X1966 3 DigitalLDOLogic_VIA0 $T=41510 23600 0 0 $X=41260 $Y=23360
X1967 3 DigitalLDOLogic_VIA0 $T=41510 29040 0 0 $X=41260 $Y=28800
X1968 3 DigitalLDOLogic_VIA0 $T=41510 34480 0 0 $X=41260 $Y=34240
X1969 3 DigitalLDOLogic_VIA0 $T=41510 39920 0 0 $X=41260 $Y=39680
X1970 3 DigitalLDOLogic_VIA0 $T=41510 45360 0 0 $X=41260 $Y=45120
X1971 3 DigitalLDOLogic_VIA0 $T=41510 50800 0 0 $X=41260 $Y=50560
X1972 3 DigitalLDOLogic_VIA0 $T=41510 56240 0 0 $X=41260 $Y=56000
X1973 1 DigitalLDOLogic_VIA0 $T=42430 15440 0 0 $X=42180 $Y=15200
X1974 1 DigitalLDOLogic_VIA0 $T=42430 20880 0 0 $X=42180 $Y=20640
X1975 1 DigitalLDOLogic_VIA0 $T=42430 26320 0 0 $X=42180 $Y=26080
X1976 1 DigitalLDOLogic_VIA0 $T=42430 31760 0 0 $X=42180 $Y=31520
X1977 1 DigitalLDOLogic_VIA0 $T=42430 37200 0 0 $X=42180 $Y=36960
X1978 1 DigitalLDOLogic_VIA0 $T=42430 42640 0 0 $X=42180 $Y=42400
X1979 1 DigitalLDOLogic_VIA0 $T=42430 48080 0 0 $X=42180 $Y=47840
X1980 1 DigitalLDOLogic_VIA0 $T=42430 53520 0 0 $X=42180 $Y=53280
X1981 1 DigitalLDOLogic_VIA0 $T=42430 58960 0 0 $X=42180 $Y=58720
X1982 3 DigitalLDOLogic_VIA0 $T=44270 12720 0 0 $X=44020 $Y=12480
X1983 3 DigitalLDOLogic_VIA0 $T=44270 18160 0 0 $X=44020 $Y=17920
X1984 3 DigitalLDOLogic_VIA0 $T=44270 23600 0 0 $X=44020 $Y=23360
X1985 3 DigitalLDOLogic_VIA0 $T=44270 29040 0 0 $X=44020 $Y=28800
X1986 3 DigitalLDOLogic_VIA0 $T=44270 34480 0 0 $X=44020 $Y=34240
X1987 3 DigitalLDOLogic_VIA0 $T=44270 39920 0 0 $X=44020 $Y=39680
X1988 3 DigitalLDOLogic_VIA0 $T=44270 45360 0 0 $X=44020 $Y=45120
X1989 3 DigitalLDOLogic_VIA0 $T=44270 50800 0 0 $X=44020 $Y=50560
X1990 3 DigitalLDOLogic_VIA0 $T=44270 56240 0 0 $X=44020 $Y=56000
X1991 1 DigitalLDOLogic_VIA0 $T=45190 15440 0 0 $X=44940 $Y=15200
X1992 1 DigitalLDOLogic_VIA0 $T=45190 20880 0 0 $X=44940 $Y=20640
X1993 1 DigitalLDOLogic_VIA0 $T=45190 26320 0 0 $X=44940 $Y=26080
X1994 1 DigitalLDOLogic_VIA0 $T=45190 31760 0 0 $X=44940 $Y=31520
X1995 1 DigitalLDOLogic_VIA0 $T=45190 37200 0 0 $X=44940 $Y=36960
X1996 1 DigitalLDOLogic_VIA0 $T=45190 42640 0 0 $X=44940 $Y=42400
X1997 1 DigitalLDOLogic_VIA0 $T=45190 48080 0 0 $X=44940 $Y=47840
X1998 1 DigitalLDOLogic_VIA0 $T=45190 53520 0 0 $X=44940 $Y=53280
X1999 1 DigitalLDOLogic_VIA0 $T=45190 58960 0 0 $X=44940 $Y=58720
X2000 3 DigitalLDOLogic_VIA0 $T=47030 12720 0 0 $X=46780 $Y=12480
X2001 3 DigitalLDOLogic_VIA0 $T=47030 18160 0 0 $X=46780 $Y=17920
X2002 3 DigitalLDOLogic_VIA0 $T=47030 23600 0 0 $X=46780 $Y=23360
X2003 3 DigitalLDOLogic_VIA0 $T=47030 29040 0 0 $X=46780 $Y=28800
X2004 3 DigitalLDOLogic_VIA0 $T=47030 34480 0 0 $X=46780 $Y=34240
X2005 3 DigitalLDOLogic_VIA0 $T=47030 39920 0 0 $X=46780 $Y=39680
X2006 3 DigitalLDOLogic_VIA0 $T=47030 45360 0 0 $X=46780 $Y=45120
X2007 3 DigitalLDOLogic_VIA0 $T=47030 50800 0 0 $X=46780 $Y=50560
X2008 3 DigitalLDOLogic_VIA0 $T=47030 56240 0 0 $X=46780 $Y=56000
X2009 1 DigitalLDOLogic_VIA0 $T=47950 15440 0 0 $X=47700 $Y=15200
X2010 1 DigitalLDOLogic_VIA0 $T=47950 20880 0 0 $X=47700 $Y=20640
X2011 1 DigitalLDOLogic_VIA0 $T=47950 26320 0 0 $X=47700 $Y=26080
X2012 1 DigitalLDOLogic_VIA0 $T=47950 31760 0 0 $X=47700 $Y=31520
X2013 1 DigitalLDOLogic_VIA0 $T=47950 37200 0 0 $X=47700 $Y=36960
X2014 1 DigitalLDOLogic_VIA0 $T=47950 42640 0 0 $X=47700 $Y=42400
X2015 1 DigitalLDOLogic_VIA0 $T=47950 48080 0 0 $X=47700 $Y=47840
X2016 1 DigitalLDOLogic_VIA0 $T=47950 53520 0 0 $X=47700 $Y=53280
X2017 1 DigitalLDOLogic_VIA0 $T=47950 58960 0 0 $X=47700 $Y=58720
X2018 3 DigitalLDOLogic_VIA0 $T=49790 12720 0 0 $X=49540 $Y=12480
X2019 3 DigitalLDOLogic_VIA0 $T=49790 18160 0 0 $X=49540 $Y=17920
X2020 3 DigitalLDOLogic_VIA0 $T=49790 23600 0 0 $X=49540 $Y=23360
X2021 3 DigitalLDOLogic_VIA0 $T=49790 29040 0 0 $X=49540 $Y=28800
X2022 3 DigitalLDOLogic_VIA0 $T=49790 34480 0 0 $X=49540 $Y=34240
X2023 3 DigitalLDOLogic_VIA0 $T=49790 39920 0 0 $X=49540 $Y=39680
X2024 3 DigitalLDOLogic_VIA0 $T=49790 45360 0 0 $X=49540 $Y=45120
X2025 3 DigitalLDOLogic_VIA0 $T=49790 50800 0 0 $X=49540 $Y=50560
X2026 3 DigitalLDOLogic_VIA0 $T=49790 56240 0 0 $X=49540 $Y=56000
X2027 1 DigitalLDOLogic_VIA0 $T=50710 15440 0 0 $X=50460 $Y=15200
X2028 1 DigitalLDOLogic_VIA0 $T=50710 20880 0 0 $X=50460 $Y=20640
X2029 1 DigitalLDOLogic_VIA0 $T=50710 26320 0 0 $X=50460 $Y=26080
X2030 1 DigitalLDOLogic_VIA0 $T=50710 31760 0 0 $X=50460 $Y=31520
X2031 1 DigitalLDOLogic_VIA0 $T=50710 37200 0 0 $X=50460 $Y=36960
X2032 1 DigitalLDOLogic_VIA0 $T=50710 42640 0 0 $X=50460 $Y=42400
X2033 1 DigitalLDOLogic_VIA0 $T=50710 48080 0 0 $X=50460 $Y=47840
X2034 1 DigitalLDOLogic_VIA0 $T=50710 53520 0 0 $X=50460 $Y=53280
X2035 1 DigitalLDOLogic_VIA0 $T=50710 58960 0 0 $X=50460 $Y=58720
X2036 3 DigitalLDOLogic_VIA0 $T=52550 12720 0 0 $X=52300 $Y=12480
X2037 3 DigitalLDOLogic_VIA0 $T=52550 18160 0 0 $X=52300 $Y=17920
X2038 3 DigitalLDOLogic_VIA0 $T=52550 23600 0 0 $X=52300 $Y=23360
X2039 3 DigitalLDOLogic_VIA0 $T=52550 29040 0 0 $X=52300 $Y=28800
X2040 3 DigitalLDOLogic_VIA0 $T=52550 34480 0 0 $X=52300 $Y=34240
X2041 3 DigitalLDOLogic_VIA0 $T=52550 39920 0 0 $X=52300 $Y=39680
X2042 3 DigitalLDOLogic_VIA0 $T=52550 45360 0 0 $X=52300 $Y=45120
X2043 3 DigitalLDOLogic_VIA0 $T=52550 50800 0 0 $X=52300 $Y=50560
X2044 3 DigitalLDOLogic_VIA0 $T=52550 56240 0 0 $X=52300 $Y=56000
X2045 1 DigitalLDOLogic_VIA0 $T=53470 15440 0 0 $X=53220 $Y=15200
X2046 1 DigitalLDOLogic_VIA0 $T=53470 20880 0 0 $X=53220 $Y=20640
X2047 1 DigitalLDOLogic_VIA0 $T=53470 26320 0 0 $X=53220 $Y=26080
X2048 1 DigitalLDOLogic_VIA0 $T=53470 31760 0 0 $X=53220 $Y=31520
X2049 1 DigitalLDOLogic_VIA0 $T=53470 37200 0 0 $X=53220 $Y=36960
X2050 1 DigitalLDOLogic_VIA0 $T=53470 42640 0 0 $X=53220 $Y=42400
X2051 1 DigitalLDOLogic_VIA0 $T=53470 48080 0 0 $X=53220 $Y=47840
X2052 1 DigitalLDOLogic_VIA0 $T=53470 53520 0 0 $X=53220 $Y=53280
X2053 1 DigitalLDOLogic_VIA0 $T=53470 58960 0 0 $X=53220 $Y=58720
X2054 3 DigitalLDOLogic_VIA0 $T=55310 12720 0 0 $X=55060 $Y=12480
X2055 3 DigitalLDOLogic_VIA0 $T=55310 18160 0 0 $X=55060 $Y=17920
X2056 3 DigitalLDOLogic_VIA0 $T=55310 23600 0 0 $X=55060 $Y=23360
X2057 3 DigitalLDOLogic_VIA0 $T=55310 29040 0 0 $X=55060 $Y=28800
X2058 3 DigitalLDOLogic_VIA0 $T=55310 34480 0 0 $X=55060 $Y=34240
X2059 3 DigitalLDOLogic_VIA0 $T=55310 39920 0 0 $X=55060 $Y=39680
X2060 3 DigitalLDOLogic_VIA0 $T=55310 45360 0 0 $X=55060 $Y=45120
X2061 3 DigitalLDOLogic_VIA0 $T=55310 50800 0 0 $X=55060 $Y=50560
X2062 3 DigitalLDOLogic_VIA0 $T=55310 56240 0 0 $X=55060 $Y=56000
X2063 1 DigitalLDOLogic_VIA0 $T=56230 15440 0 0 $X=55980 $Y=15200
X2064 1 DigitalLDOLogic_VIA0 $T=56230 20880 0 0 $X=55980 $Y=20640
X2065 1 DigitalLDOLogic_VIA0 $T=56230 26320 0 0 $X=55980 $Y=26080
X2066 1 DigitalLDOLogic_VIA0 $T=56230 31760 0 0 $X=55980 $Y=31520
X2067 1 DigitalLDOLogic_VIA0 $T=56230 37200 0 0 $X=55980 $Y=36960
X2068 1 DigitalLDOLogic_VIA0 $T=56230 42640 0 0 $X=55980 $Y=42400
X2069 1 DigitalLDOLogic_VIA0 $T=56230 48080 0 0 $X=55980 $Y=47840
X2070 1 DigitalLDOLogic_VIA0 $T=56230 53520 0 0 $X=55980 $Y=53280
X2071 1 DigitalLDOLogic_VIA0 $T=56230 58960 0 0 $X=55980 $Y=58720
X2072 3 DigitalLDOLogic_VIA0 $T=58070 12720 0 0 $X=57820 $Y=12480
X2073 3 DigitalLDOLogic_VIA0 $T=58070 18160 0 0 $X=57820 $Y=17920
X2074 3 DigitalLDOLogic_VIA0 $T=58070 23600 0 0 $X=57820 $Y=23360
X2075 3 DigitalLDOLogic_VIA0 $T=58070 29040 0 0 $X=57820 $Y=28800
X2076 3 DigitalLDOLogic_VIA0 $T=58070 34480 0 0 $X=57820 $Y=34240
X2077 3 DigitalLDOLogic_VIA0 $T=58070 39920 0 0 $X=57820 $Y=39680
X2078 3 DigitalLDOLogic_VIA0 $T=58070 45360 0 0 $X=57820 $Y=45120
X2079 3 DigitalLDOLogic_VIA0 $T=58070 50800 0 0 $X=57820 $Y=50560
X2080 3 DigitalLDOLogic_VIA0 $T=58070 56240 0 0 $X=57820 $Y=56000
X2081 1 DigitalLDOLogic_VIA0 $T=58990 15440 0 0 $X=58740 $Y=15200
X2082 1 DigitalLDOLogic_VIA0 $T=58990 20880 0 0 $X=58740 $Y=20640
X2083 1 DigitalLDOLogic_VIA0 $T=58990 26320 0 0 $X=58740 $Y=26080
X2084 1 DigitalLDOLogic_VIA0 $T=58990 31760 0 0 $X=58740 $Y=31520
X2085 1 DigitalLDOLogic_VIA0 $T=58990 37200 0 0 $X=58740 $Y=36960
X2086 1 DigitalLDOLogic_VIA0 $T=58990 42640 0 0 $X=58740 $Y=42400
X2087 1 DigitalLDOLogic_VIA0 $T=58990 48080 0 0 $X=58740 $Y=47840
X2088 1 DigitalLDOLogic_VIA0 $T=58990 53520 0 0 $X=58740 $Y=53280
X2089 1 DigitalLDOLogic_VIA0 $T=58990 58960 0 0 $X=58740 $Y=58720
X2090 3 DigitalLDOLogic_VIA0 $T=60830 12720 0 0 $X=60580 $Y=12480
X2091 3 DigitalLDOLogic_VIA0 $T=60830 18160 0 0 $X=60580 $Y=17920
X2092 3 DigitalLDOLogic_VIA0 $T=60830 23600 0 0 $X=60580 $Y=23360
X2093 3 DigitalLDOLogic_VIA0 $T=60830 29040 0 0 $X=60580 $Y=28800
X2094 3 DigitalLDOLogic_VIA0 $T=60830 34480 0 0 $X=60580 $Y=34240
X2095 3 DigitalLDOLogic_VIA0 $T=60830 39920 0 0 $X=60580 $Y=39680
X2096 3 DigitalLDOLogic_VIA0 $T=60830 45360 0 0 $X=60580 $Y=45120
X2097 3 DigitalLDOLogic_VIA0 $T=60830 50800 0 0 $X=60580 $Y=50560
X2098 3 DigitalLDOLogic_VIA0 $T=60830 56240 0 0 $X=60580 $Y=56000
X2099 1 DigitalLDOLogic_VIA0 $T=61750 15440 0 0 $X=61500 $Y=15200
X2100 1 DigitalLDOLogic_VIA0 $T=61750 20880 0 0 $X=61500 $Y=20640
X2101 1 DigitalLDOLogic_VIA0 $T=61750 26320 0 0 $X=61500 $Y=26080
X2102 1 DigitalLDOLogic_VIA0 $T=61750 31760 0 0 $X=61500 $Y=31520
X2103 1 DigitalLDOLogic_VIA0 $T=61750 37200 0 0 $X=61500 $Y=36960
X2104 1 DigitalLDOLogic_VIA0 $T=61750 42640 0 0 $X=61500 $Y=42400
X2105 1 DigitalLDOLogic_VIA0 $T=61750 48080 0 0 $X=61500 $Y=47840
X2106 1 DigitalLDOLogic_VIA0 $T=61750 53520 0 0 $X=61500 $Y=53280
X2107 1 DigitalLDOLogic_VIA0 $T=61750 58960 0 0 $X=61500 $Y=58720
X2108 3 DigitalLDOLogic_VIA0 $T=63590 12720 0 0 $X=63340 $Y=12480
X2109 3 DigitalLDOLogic_VIA0 $T=63590 18160 0 0 $X=63340 $Y=17920
X2110 3 DigitalLDOLogic_VIA0 $T=63590 23600 0 0 $X=63340 $Y=23360
X2111 3 DigitalLDOLogic_VIA0 $T=63590 29040 0 0 $X=63340 $Y=28800
X2112 3 DigitalLDOLogic_VIA0 $T=63590 34480 0 0 $X=63340 $Y=34240
X2113 3 DigitalLDOLogic_VIA0 $T=63590 39920 0 0 $X=63340 $Y=39680
X2114 3 DigitalLDOLogic_VIA0 $T=63590 45360 0 0 $X=63340 $Y=45120
X2115 3 DigitalLDOLogic_VIA0 $T=63590 50800 0 0 $X=63340 $Y=50560
X2116 3 DigitalLDOLogic_VIA0 $T=63590 56240 0 0 $X=63340 $Y=56000
X2117 1 DigitalLDOLogic_VIA0 $T=64510 15440 0 0 $X=64260 $Y=15200
X2118 1 DigitalLDOLogic_VIA0 $T=64510 20880 0 0 $X=64260 $Y=20640
X2119 1 DigitalLDOLogic_VIA0 $T=64510 26320 0 0 $X=64260 $Y=26080
X2120 1 DigitalLDOLogic_VIA0 $T=64510 31760 0 0 $X=64260 $Y=31520
X2121 1 DigitalLDOLogic_VIA0 $T=64510 37200 0 0 $X=64260 $Y=36960
X2122 1 DigitalLDOLogic_VIA0 $T=64510 42640 0 0 $X=64260 $Y=42400
X2123 1 DigitalLDOLogic_VIA0 $T=64510 48080 0 0 $X=64260 $Y=47840
X2124 1 DigitalLDOLogic_VIA0 $T=64510 53520 0 0 $X=64260 $Y=53280
X2125 1 DigitalLDOLogic_VIA0 $T=64510 58960 0 0 $X=64260 $Y=58720
X2126 3 DigitalLDOLogic_VIA0 $T=66350 12720 0 0 $X=66100 $Y=12480
X2127 3 DigitalLDOLogic_VIA0 $T=66350 18160 0 0 $X=66100 $Y=17920
X2128 3 DigitalLDOLogic_VIA0 $T=66350 23600 0 0 $X=66100 $Y=23360
X2129 3 DigitalLDOLogic_VIA0 $T=66350 29040 0 0 $X=66100 $Y=28800
X2130 3 DigitalLDOLogic_VIA0 $T=66350 34480 0 0 $X=66100 $Y=34240
X2131 3 DigitalLDOLogic_VIA0 $T=66350 39920 0 0 $X=66100 $Y=39680
X2132 3 DigitalLDOLogic_VIA0 $T=66350 45360 0 0 $X=66100 $Y=45120
X2133 3 DigitalLDOLogic_VIA0 $T=66350 50800 0 0 $X=66100 $Y=50560
X2134 3 DigitalLDOLogic_VIA0 $T=66350 56240 0 0 $X=66100 $Y=56000
X2135 1 DigitalLDOLogic_VIA0 $T=67270 15440 0 0 $X=67020 $Y=15200
X2136 1 DigitalLDOLogic_VIA0 $T=67270 20880 0 0 $X=67020 $Y=20640
X2137 1 DigitalLDOLogic_VIA0 $T=67270 26320 0 0 $X=67020 $Y=26080
X2138 1 DigitalLDOLogic_VIA0 $T=67270 31760 0 0 $X=67020 $Y=31520
X2139 1 DigitalLDOLogic_VIA0 $T=67270 37200 0 0 $X=67020 $Y=36960
X2140 1 DigitalLDOLogic_VIA0 $T=67270 42640 0 0 $X=67020 $Y=42400
X2141 1 DigitalLDOLogic_VIA0 $T=67270 48080 0 0 $X=67020 $Y=47840
X2142 1 DigitalLDOLogic_VIA0 $T=67270 53520 0 0 $X=67020 $Y=53280
X2143 1 DigitalLDOLogic_VIA0 $T=67270 58960 0 0 $X=67020 $Y=58720
X2144 3 DigitalLDOLogic_VIA0 $T=69110 12720 0 0 $X=68860 $Y=12480
X2145 3 DigitalLDOLogic_VIA0 $T=69110 18160 0 0 $X=68860 $Y=17920
X2146 3 DigitalLDOLogic_VIA0 $T=69110 23600 0 0 $X=68860 $Y=23360
X2147 3 DigitalLDOLogic_VIA0 $T=69110 29040 0 0 $X=68860 $Y=28800
X2148 3 DigitalLDOLogic_VIA0 $T=69110 34480 0 0 $X=68860 $Y=34240
X2149 3 DigitalLDOLogic_VIA0 $T=69110 39920 0 0 $X=68860 $Y=39680
X2150 3 DigitalLDOLogic_VIA0 $T=69110 45360 0 0 $X=68860 $Y=45120
X2151 3 DigitalLDOLogic_VIA0 $T=69110 50800 0 0 $X=68860 $Y=50560
X2152 3 DigitalLDOLogic_VIA0 $T=69110 56240 0 0 $X=68860 $Y=56000
X2153 1 DigitalLDOLogic_VIA0 $T=70030 15440 0 0 $X=69780 $Y=15200
X2154 1 DigitalLDOLogic_VIA0 $T=70030 20880 0 0 $X=69780 $Y=20640
X2155 1 DigitalLDOLogic_VIA0 $T=70030 26320 0 0 $X=69780 $Y=26080
X2156 1 DigitalLDOLogic_VIA0 $T=70030 31760 0 0 $X=69780 $Y=31520
X2157 1 DigitalLDOLogic_VIA0 $T=70030 37200 0 0 $X=69780 $Y=36960
X2158 1 DigitalLDOLogic_VIA0 $T=70030 42640 0 0 $X=69780 $Y=42400
X2159 1 DigitalLDOLogic_VIA0 $T=70030 48080 0 0 $X=69780 $Y=47840
X2160 1 DigitalLDOLogic_VIA0 $T=70030 53520 0 0 $X=69780 $Y=53280
X2161 1 DigitalLDOLogic_VIA0 $T=70030 58960 0 0 $X=69780 $Y=58720
X2162 3 DigitalLDOLogic_VIA0 $T=71870 12720 0 0 $X=71620 $Y=12480
X2163 3 DigitalLDOLogic_VIA0 $T=71870 18160 0 0 $X=71620 $Y=17920
X2164 3 DigitalLDOLogic_VIA0 $T=71870 23600 0 0 $X=71620 $Y=23360
X2165 3 DigitalLDOLogic_VIA0 $T=71870 29040 0 0 $X=71620 $Y=28800
X2166 3 DigitalLDOLogic_VIA0 $T=71870 34480 0 0 $X=71620 $Y=34240
X2167 3 DigitalLDOLogic_VIA0 $T=71870 39920 0 0 $X=71620 $Y=39680
X2168 3 DigitalLDOLogic_VIA0 $T=71870 45360 0 0 $X=71620 $Y=45120
X2169 3 DigitalLDOLogic_VIA0 $T=71870 50800 0 0 $X=71620 $Y=50560
X2170 3 DigitalLDOLogic_VIA0 $T=71870 56240 0 0 $X=71620 $Y=56000
X2171 1 DigitalLDOLogic_VIA0 $T=72790 15440 0 0 $X=72540 $Y=15200
X2172 1 DigitalLDOLogic_VIA0 $T=72790 20880 0 0 $X=72540 $Y=20640
X2173 1 DigitalLDOLogic_VIA0 $T=72790 26320 0 0 $X=72540 $Y=26080
X2174 1 DigitalLDOLogic_VIA0 $T=72790 31760 0 0 $X=72540 $Y=31520
X2175 1 DigitalLDOLogic_VIA0 $T=72790 37200 0 0 $X=72540 $Y=36960
X2176 1 DigitalLDOLogic_VIA0 $T=72790 42640 0 0 $X=72540 $Y=42400
X2177 1 DigitalLDOLogic_VIA0 $T=72790 48080 0 0 $X=72540 $Y=47840
X2178 1 DigitalLDOLogic_VIA0 $T=72790 53520 0 0 $X=72540 $Y=53280
X2179 1 DigitalLDOLogic_VIA0 $T=72790 58960 0 0 $X=72540 $Y=58720
X2180 3 DigitalLDOLogic_VIA0 $T=74630 12720 0 0 $X=74380 $Y=12480
X2181 3 DigitalLDOLogic_VIA0 $T=74630 18160 0 0 $X=74380 $Y=17920
X2182 3 DigitalLDOLogic_VIA0 $T=74630 23600 0 0 $X=74380 $Y=23360
X2183 3 DigitalLDOLogic_VIA0 $T=74630 29040 0 0 $X=74380 $Y=28800
X2184 3 DigitalLDOLogic_VIA0 $T=74630 34480 0 0 $X=74380 $Y=34240
X2185 3 DigitalLDOLogic_VIA0 $T=74630 39920 0 0 $X=74380 $Y=39680
X2186 3 DigitalLDOLogic_VIA0 $T=74630 45360 0 0 $X=74380 $Y=45120
X2187 3 DigitalLDOLogic_VIA0 $T=74630 50800 0 0 $X=74380 $Y=50560
X2188 3 DigitalLDOLogic_VIA0 $T=74630 56240 0 0 $X=74380 $Y=56000
X2189 1 DigitalLDOLogic_VIA0 $T=75550 15440 0 0 $X=75300 $Y=15200
X2190 1 DigitalLDOLogic_VIA0 $T=75550 20880 0 0 $X=75300 $Y=20640
X2191 1 DigitalLDOLogic_VIA0 $T=75550 26320 0 0 $X=75300 $Y=26080
X2192 1 DigitalLDOLogic_VIA0 $T=75550 31760 0 0 $X=75300 $Y=31520
X2193 1 DigitalLDOLogic_VIA0 $T=75550 37200 0 0 $X=75300 $Y=36960
X2194 1 DigitalLDOLogic_VIA0 $T=75550 42640 0 0 $X=75300 $Y=42400
X2195 1 DigitalLDOLogic_VIA0 $T=75550 48080 0 0 $X=75300 $Y=47840
X2196 1 DigitalLDOLogic_VIA0 $T=75550 53520 0 0 $X=75300 $Y=53280
X2197 1 DigitalLDOLogic_VIA0 $T=75550 58960 0 0 $X=75300 $Y=58720
X2198 3 DigitalLDOLogic_VIA0 $T=77390 12720 0 0 $X=77140 $Y=12480
X2199 3 DigitalLDOLogic_VIA0 $T=77390 18160 0 0 $X=77140 $Y=17920
X2200 3 DigitalLDOLogic_VIA0 $T=77390 23600 0 0 $X=77140 $Y=23360
X2201 3 DigitalLDOLogic_VIA0 $T=77390 29040 0 0 $X=77140 $Y=28800
X2202 3 DigitalLDOLogic_VIA0 $T=77390 34480 0 0 $X=77140 $Y=34240
X2203 3 DigitalLDOLogic_VIA0 $T=77390 39920 0 0 $X=77140 $Y=39680
X2204 3 DigitalLDOLogic_VIA0 $T=77390 45360 0 0 $X=77140 $Y=45120
X2205 3 DigitalLDOLogic_VIA0 $T=77390 50800 0 0 $X=77140 $Y=50560
X2206 3 DigitalLDOLogic_VIA0 $T=77390 56240 0 0 $X=77140 $Y=56000
X2207 1 DigitalLDOLogic_VIA0 $T=78310 15440 0 0 $X=78060 $Y=15200
X2208 1 DigitalLDOLogic_VIA0 $T=78310 20880 0 0 $X=78060 $Y=20640
X2209 1 DigitalLDOLogic_VIA0 $T=78310 26320 0 0 $X=78060 $Y=26080
X2210 1 DigitalLDOLogic_VIA0 $T=78310 31760 0 0 $X=78060 $Y=31520
X2211 1 DigitalLDOLogic_VIA0 $T=78310 37200 0 0 $X=78060 $Y=36960
X2212 1 DigitalLDOLogic_VIA0 $T=78310 42640 0 0 $X=78060 $Y=42400
X2213 1 DigitalLDOLogic_VIA0 $T=78310 48080 0 0 $X=78060 $Y=47840
X2214 1 DigitalLDOLogic_VIA0 $T=78310 53520 0 0 $X=78060 $Y=53280
X2215 1 DigitalLDOLogic_VIA0 $T=78310 58960 0 0 $X=78060 $Y=58720
X2216 3 DigitalLDOLogic_VIA0 $T=80150 12720 0 0 $X=79900 $Y=12480
X2217 3 DigitalLDOLogic_VIA0 $T=80150 18160 0 0 $X=79900 $Y=17920
X2218 3 DigitalLDOLogic_VIA0 $T=80150 23600 0 0 $X=79900 $Y=23360
X2219 3 DigitalLDOLogic_VIA0 $T=80150 29040 0 0 $X=79900 $Y=28800
X2220 3 DigitalLDOLogic_VIA0 $T=80150 34480 0 0 $X=79900 $Y=34240
X2221 3 DigitalLDOLogic_VIA0 $T=80150 39920 0 0 $X=79900 $Y=39680
X2222 3 DigitalLDOLogic_VIA0 $T=80150 45360 0 0 $X=79900 $Y=45120
X2223 3 DigitalLDOLogic_VIA0 $T=80150 50800 0 0 $X=79900 $Y=50560
X2224 3 DigitalLDOLogic_VIA0 $T=80150 56240 0 0 $X=79900 $Y=56000
X2225 1 DigitalLDOLogic_VIA0 $T=81070 15440 0 0 $X=80820 $Y=15200
X2226 1 DigitalLDOLogic_VIA0 $T=81070 20880 0 0 $X=80820 $Y=20640
X2227 1 DigitalLDOLogic_VIA0 $T=81070 26320 0 0 $X=80820 $Y=26080
X2228 1 DigitalLDOLogic_VIA0 $T=81070 31760 0 0 $X=80820 $Y=31520
X2229 1 DigitalLDOLogic_VIA0 $T=81070 37200 0 0 $X=80820 $Y=36960
X2230 1 DigitalLDOLogic_VIA0 $T=81070 42640 0 0 $X=80820 $Y=42400
X2231 1 DigitalLDOLogic_VIA0 $T=81070 48080 0 0 $X=80820 $Y=47840
X2232 1 DigitalLDOLogic_VIA0 $T=81070 53520 0 0 $X=80820 $Y=53280
X2233 1 DigitalLDOLogic_VIA0 $T=81070 58960 0 0 $X=80820 $Y=58720
X2234 3 DigitalLDOLogic_VIA0 $T=82910 12720 0 0 $X=82660 $Y=12480
X2235 3 DigitalLDOLogic_VIA0 $T=82910 18160 0 0 $X=82660 $Y=17920
X2236 3 DigitalLDOLogic_VIA0 $T=82910 23600 0 0 $X=82660 $Y=23360
X2237 3 DigitalLDOLogic_VIA0 $T=82910 29040 0 0 $X=82660 $Y=28800
X2238 3 DigitalLDOLogic_VIA0 $T=82910 34480 0 0 $X=82660 $Y=34240
X2239 3 DigitalLDOLogic_VIA0 $T=82910 39920 0 0 $X=82660 $Y=39680
X2240 3 DigitalLDOLogic_VIA0 $T=82910 45360 0 0 $X=82660 $Y=45120
X2241 3 DigitalLDOLogic_VIA0 $T=82910 50800 0 0 $X=82660 $Y=50560
X2242 3 DigitalLDOLogic_VIA0 $T=82910 56240 0 0 $X=82660 $Y=56000
X2243 1 DigitalLDOLogic_VIA0 $T=83830 15440 0 0 $X=83580 $Y=15200
X2244 1 DigitalLDOLogic_VIA0 $T=83830 20880 0 0 $X=83580 $Y=20640
X2245 1 DigitalLDOLogic_VIA0 $T=83830 26320 0 0 $X=83580 $Y=26080
X2246 1 DigitalLDOLogic_VIA0 $T=83830 31760 0 0 $X=83580 $Y=31520
X2247 1 DigitalLDOLogic_VIA0 $T=83830 37200 0 0 $X=83580 $Y=36960
X2248 1 DigitalLDOLogic_VIA0 $T=83830 42640 0 0 $X=83580 $Y=42400
X2249 1 DigitalLDOLogic_VIA0 $T=83830 48080 0 0 $X=83580 $Y=47840
X2250 1 DigitalLDOLogic_VIA0 $T=83830 53520 0 0 $X=83580 $Y=53280
X2251 1 DigitalLDOLogic_VIA0 $T=83830 58960 0 0 $X=83580 $Y=58720
X2252 3 DigitalLDOLogic_VIA0 $T=85670 12720 0 0 $X=85420 $Y=12480
X2253 3 DigitalLDOLogic_VIA0 $T=85670 18160 0 0 $X=85420 $Y=17920
X2254 3 DigitalLDOLogic_VIA0 $T=85670 23600 0 0 $X=85420 $Y=23360
X2255 3 DigitalLDOLogic_VIA0 $T=85670 29040 0 0 $X=85420 $Y=28800
X2256 3 DigitalLDOLogic_VIA0 $T=85670 34480 0 0 $X=85420 $Y=34240
X2257 3 DigitalLDOLogic_VIA0 $T=85670 39920 0 0 $X=85420 $Y=39680
X2258 3 DigitalLDOLogic_VIA0 $T=85670 45360 0 0 $X=85420 $Y=45120
X2259 3 DigitalLDOLogic_VIA0 $T=85670 50800 0 0 $X=85420 $Y=50560
X2260 3 DigitalLDOLogic_VIA0 $T=85670 56240 0 0 $X=85420 $Y=56000
X2261 1 DigitalLDOLogic_VIA0 $T=86590 15440 0 0 $X=86340 $Y=15200
X2262 1 DigitalLDOLogic_VIA0 $T=86590 20880 0 0 $X=86340 $Y=20640
X2263 1 DigitalLDOLogic_VIA0 $T=86590 26320 0 0 $X=86340 $Y=26080
X2264 1 DigitalLDOLogic_VIA0 $T=86590 31760 0 0 $X=86340 $Y=31520
X2265 1 DigitalLDOLogic_VIA0 $T=86590 37200 0 0 $X=86340 $Y=36960
X2266 1 DigitalLDOLogic_VIA0 $T=86590 42640 0 0 $X=86340 $Y=42400
X2267 1 DigitalLDOLogic_VIA0 $T=86590 48080 0 0 $X=86340 $Y=47840
X2268 1 DigitalLDOLogic_VIA0 $T=86590 53520 0 0 $X=86340 $Y=53280
X2269 1 DigitalLDOLogic_VIA0 $T=86590 58960 0 0 $X=86340 $Y=58720
X2270 3 DigitalLDOLogic_VIA0 $T=88430 12720 0 0 $X=88180 $Y=12480
X2271 3 DigitalLDOLogic_VIA0 $T=88430 18160 0 0 $X=88180 $Y=17920
X2272 3 DigitalLDOLogic_VIA0 $T=88430 23600 0 0 $X=88180 $Y=23360
X2273 3 DigitalLDOLogic_VIA0 $T=88430 29040 0 0 $X=88180 $Y=28800
X2274 3 DigitalLDOLogic_VIA0 $T=88430 34480 0 0 $X=88180 $Y=34240
X2275 3 DigitalLDOLogic_VIA0 $T=88430 39920 0 0 $X=88180 $Y=39680
X2276 3 DigitalLDOLogic_VIA0 $T=88430 45360 0 0 $X=88180 $Y=45120
X2277 3 DigitalLDOLogic_VIA0 $T=88430 50800 0 0 $X=88180 $Y=50560
X2278 3 DigitalLDOLogic_VIA0 $T=88430 56240 0 0 $X=88180 $Y=56000
X2279 1 DigitalLDOLogic_VIA0 $T=89350 15440 0 0 $X=89100 $Y=15200
X2280 1 DigitalLDOLogic_VIA0 $T=89350 20880 0 0 $X=89100 $Y=20640
X2281 1 DigitalLDOLogic_VIA0 $T=89350 26320 0 0 $X=89100 $Y=26080
X2282 1 DigitalLDOLogic_VIA0 $T=89350 31760 0 0 $X=89100 $Y=31520
X2283 1 DigitalLDOLogic_VIA0 $T=89350 37200 0 0 $X=89100 $Y=36960
X2284 1 DigitalLDOLogic_VIA0 $T=89350 42640 0 0 $X=89100 $Y=42400
X2285 1 DigitalLDOLogic_VIA0 $T=89350 48080 0 0 $X=89100 $Y=47840
X2286 1 DigitalLDOLogic_VIA0 $T=89350 53520 0 0 $X=89100 $Y=53280
X2287 1 DigitalLDOLogic_VIA0 $T=89350 58960 0 0 $X=89100 $Y=58720
X2288 3 DigitalLDOLogic_VIA0 $T=91190 12720 0 0 $X=90940 $Y=12480
X2289 3 DigitalLDOLogic_VIA0 $T=91190 18160 0 0 $X=90940 $Y=17920
X2290 3 DigitalLDOLogic_VIA0 $T=91190 23600 0 0 $X=90940 $Y=23360
X2291 3 DigitalLDOLogic_VIA0 $T=91190 29040 0 0 $X=90940 $Y=28800
X2292 3 DigitalLDOLogic_VIA0 $T=91190 34480 0 0 $X=90940 $Y=34240
X2293 3 DigitalLDOLogic_VIA0 $T=91190 39920 0 0 $X=90940 $Y=39680
X2294 3 DigitalLDOLogic_VIA0 $T=91190 45360 0 0 $X=90940 $Y=45120
X2295 3 DigitalLDOLogic_VIA0 $T=91190 50800 0 0 $X=90940 $Y=50560
X2296 3 DigitalLDOLogic_VIA0 $T=91190 56240 0 0 $X=90940 $Y=56000
X2297 1 DigitalLDOLogic_VIA0 $T=92110 15440 0 0 $X=91860 $Y=15200
X2298 1 DigitalLDOLogic_VIA0 $T=92110 20880 0 0 $X=91860 $Y=20640
X2299 1 DigitalLDOLogic_VIA0 $T=92110 26320 0 0 $X=91860 $Y=26080
X2300 1 DigitalLDOLogic_VIA0 $T=92110 31760 0 0 $X=91860 $Y=31520
X2301 1 DigitalLDOLogic_VIA0 $T=92110 37200 0 0 $X=91860 $Y=36960
X2302 1 DigitalLDOLogic_VIA0 $T=92110 42640 0 0 $X=91860 $Y=42400
X2303 1 DigitalLDOLogic_VIA0 $T=92110 48080 0 0 $X=91860 $Y=47840
X2304 1 DigitalLDOLogic_VIA0 $T=92110 53520 0 0 $X=91860 $Y=53280
X2305 1 DigitalLDOLogic_VIA0 $T=92110 58960 0 0 $X=91860 $Y=58720
X2306 3 DigitalLDOLogic_VIA0 $T=93950 12720 0 0 $X=93700 $Y=12480
X2307 3 DigitalLDOLogic_VIA0 $T=93950 18160 0 0 $X=93700 $Y=17920
X2308 3 DigitalLDOLogic_VIA0 $T=93950 23600 0 0 $X=93700 $Y=23360
X2309 3 DigitalLDOLogic_VIA0 $T=93950 29040 0 0 $X=93700 $Y=28800
X2310 3 DigitalLDOLogic_VIA0 $T=93950 34480 0 0 $X=93700 $Y=34240
X2311 3 DigitalLDOLogic_VIA0 $T=93950 39920 0 0 $X=93700 $Y=39680
X2312 3 DigitalLDOLogic_VIA0 $T=93950 45360 0 0 $X=93700 $Y=45120
X2313 3 DigitalLDOLogic_VIA0 $T=93950 50800 0 0 $X=93700 $Y=50560
X2314 3 DigitalLDOLogic_VIA0 $T=93950 56240 0 0 $X=93700 $Y=56000
X2315 1 DigitalLDOLogic_VIA0 $T=94870 15440 0 0 $X=94620 $Y=15200
X2316 1 DigitalLDOLogic_VIA0 $T=94870 20880 0 0 $X=94620 $Y=20640
X2317 1 DigitalLDOLogic_VIA0 $T=94870 26320 0 0 $X=94620 $Y=26080
X2318 1 DigitalLDOLogic_VIA0 $T=94870 31760 0 0 $X=94620 $Y=31520
X2319 1 DigitalLDOLogic_VIA0 $T=94870 37200 0 0 $X=94620 $Y=36960
X2320 1 DigitalLDOLogic_VIA0 $T=94870 42640 0 0 $X=94620 $Y=42400
X2321 1 DigitalLDOLogic_VIA0 $T=94870 48080 0 0 $X=94620 $Y=47840
X2322 1 DigitalLDOLogic_VIA0 $T=94870 53520 0 0 $X=94620 $Y=53280
X2323 1 DigitalLDOLogic_VIA0 $T=94870 58960 0 0 $X=94620 $Y=58720
X2324 3 DigitalLDOLogic_VIA0 $T=96710 12720 0 0 $X=96460 $Y=12480
X2325 3 DigitalLDOLogic_VIA0 $T=96710 18160 0 0 $X=96460 $Y=17920
X2326 3 DigitalLDOLogic_VIA0 $T=96710 23600 0 0 $X=96460 $Y=23360
X2327 3 DigitalLDOLogic_VIA0 $T=96710 29040 0 0 $X=96460 $Y=28800
X2328 3 DigitalLDOLogic_VIA0 $T=96710 34480 0 0 $X=96460 $Y=34240
X2329 3 DigitalLDOLogic_VIA0 $T=96710 39920 0 0 $X=96460 $Y=39680
X2330 3 DigitalLDOLogic_VIA0 $T=96710 45360 0 0 $X=96460 $Y=45120
X2331 3 DigitalLDOLogic_VIA0 $T=96710 50800 0 0 $X=96460 $Y=50560
X2332 3 DigitalLDOLogic_VIA0 $T=96710 56240 0 0 $X=96460 $Y=56000
X2333 1 DigitalLDOLogic_VIA0 $T=97630 15440 0 0 $X=97380 $Y=15200
X2334 1 DigitalLDOLogic_VIA0 $T=97630 20880 0 0 $X=97380 $Y=20640
X2335 1 DigitalLDOLogic_VIA0 $T=97630 26320 0 0 $X=97380 $Y=26080
X2336 1 DigitalLDOLogic_VIA0 $T=97630 31760 0 0 $X=97380 $Y=31520
X2337 1 DigitalLDOLogic_VIA0 $T=97630 37200 0 0 $X=97380 $Y=36960
X2338 1 DigitalLDOLogic_VIA0 $T=97630 42640 0 0 $X=97380 $Y=42400
X2339 1 DigitalLDOLogic_VIA0 $T=97630 48080 0 0 $X=97380 $Y=47840
X2340 1 DigitalLDOLogic_VIA0 $T=97630 53520 0 0 $X=97380 $Y=53280
X2341 1 DigitalLDOLogic_VIA0 $T=97630 58960 0 0 $X=97380 $Y=58720
X2342 3 DigitalLDOLogic_VIA0 $T=99470 12720 0 0 $X=99220 $Y=12480
X2343 3 DigitalLDOLogic_VIA0 $T=99470 18160 0 0 $X=99220 $Y=17920
X2344 3 DigitalLDOLogic_VIA0 $T=99470 23600 0 0 $X=99220 $Y=23360
X2345 3 DigitalLDOLogic_VIA0 $T=99470 29040 0 0 $X=99220 $Y=28800
X2346 3 DigitalLDOLogic_VIA0 $T=99470 34480 0 0 $X=99220 $Y=34240
X2347 3 DigitalLDOLogic_VIA0 $T=99470 39920 0 0 $X=99220 $Y=39680
X2348 3 DigitalLDOLogic_VIA0 $T=99470 45360 0 0 $X=99220 $Y=45120
X2349 3 DigitalLDOLogic_VIA0 $T=99470 50800 0 0 $X=99220 $Y=50560
X2350 3 DigitalLDOLogic_VIA0 $T=99470 56240 0 0 $X=99220 $Y=56000
X2351 1 DigitalLDOLogic_VIA0 $T=100390 15440 0 0 $X=100140 $Y=15200
X2352 1 DigitalLDOLogic_VIA0 $T=100390 20880 0 0 $X=100140 $Y=20640
X2353 1 DigitalLDOLogic_VIA0 $T=100390 26320 0 0 $X=100140 $Y=26080
X2354 1 DigitalLDOLogic_VIA0 $T=100390 31760 0 0 $X=100140 $Y=31520
X2355 1 DigitalLDOLogic_VIA0 $T=100390 37200 0 0 $X=100140 $Y=36960
X2356 1 DigitalLDOLogic_VIA0 $T=100390 42640 0 0 $X=100140 $Y=42400
X2357 1 DigitalLDOLogic_VIA0 $T=100390 48080 0 0 $X=100140 $Y=47840
X2358 1 DigitalLDOLogic_VIA0 $T=100390 53520 0 0 $X=100140 $Y=53280
X2359 1 DigitalLDOLogic_VIA0 $T=100390 58960 0 0 $X=100140 $Y=58720
X2360 3 DigitalLDOLogic_VIA0 $T=102230 12720 0 0 $X=101980 $Y=12480
X2361 3 DigitalLDOLogic_VIA0 $T=102230 18160 0 0 $X=101980 $Y=17920
X2362 3 DigitalLDOLogic_VIA0 $T=102230 23600 0 0 $X=101980 $Y=23360
X2363 3 DigitalLDOLogic_VIA0 $T=102230 29040 0 0 $X=101980 $Y=28800
X2364 3 DigitalLDOLogic_VIA0 $T=102230 34480 0 0 $X=101980 $Y=34240
X2365 3 DigitalLDOLogic_VIA0 $T=102230 39920 0 0 $X=101980 $Y=39680
X2366 3 DigitalLDOLogic_VIA0 $T=102230 45360 0 0 $X=101980 $Y=45120
X2367 3 DigitalLDOLogic_VIA0 $T=102230 50800 0 0 $X=101980 $Y=50560
X2368 3 DigitalLDOLogic_VIA0 $T=102230 56240 0 0 $X=101980 $Y=56000
X2369 1 DigitalLDOLogic_VIA0 $T=103150 15440 0 0 $X=102900 $Y=15200
X2370 1 DigitalLDOLogic_VIA0 $T=103150 20880 0 0 $X=102900 $Y=20640
X2371 1 DigitalLDOLogic_VIA0 $T=103150 26320 0 0 $X=102900 $Y=26080
X2372 1 DigitalLDOLogic_VIA0 $T=103150 31760 0 0 $X=102900 $Y=31520
X2373 1 DigitalLDOLogic_VIA0 $T=103150 37200 0 0 $X=102900 $Y=36960
X2374 1 DigitalLDOLogic_VIA0 $T=103150 42640 0 0 $X=102900 $Y=42400
X2375 1 DigitalLDOLogic_VIA0 $T=103150 48080 0 0 $X=102900 $Y=47840
X2376 1 DigitalLDOLogic_VIA0 $T=103150 53520 0 0 $X=102900 $Y=53280
X2377 1 DigitalLDOLogic_VIA0 $T=103150 58960 0 0 $X=102900 $Y=58720
X2378 3 DigitalLDOLogic_VIA0 $T=104990 12720 0 0 $X=104740 $Y=12480
X2379 3 DigitalLDOLogic_VIA0 $T=104990 18160 0 0 $X=104740 $Y=17920
X2380 3 DigitalLDOLogic_VIA0 $T=104990 23600 0 0 $X=104740 $Y=23360
X2381 3 DigitalLDOLogic_VIA0 $T=104990 29040 0 0 $X=104740 $Y=28800
X2382 3 DigitalLDOLogic_VIA0 $T=104990 34480 0 0 $X=104740 $Y=34240
X2383 3 DigitalLDOLogic_VIA0 $T=104990 39920 0 0 $X=104740 $Y=39680
X2384 3 DigitalLDOLogic_VIA0 $T=104990 45360 0 0 $X=104740 $Y=45120
X2385 3 DigitalLDOLogic_VIA0 $T=104990 50800 0 0 $X=104740 $Y=50560
X2386 3 DigitalLDOLogic_VIA0 $T=104990 56240 0 0 $X=104740 $Y=56000
X2387 1 DigitalLDOLogic_VIA0 $T=105910 15440 0 0 $X=105660 $Y=15200
X2388 1 DigitalLDOLogic_VIA0 $T=105910 20880 0 0 $X=105660 $Y=20640
X2389 1 DigitalLDOLogic_VIA0 $T=105910 26320 0 0 $X=105660 $Y=26080
X2390 1 DigitalLDOLogic_VIA0 $T=105910 31760 0 0 $X=105660 $Y=31520
X2391 1 DigitalLDOLogic_VIA0 $T=105910 37200 0 0 $X=105660 $Y=36960
X2392 1 DigitalLDOLogic_VIA0 $T=105910 42640 0 0 $X=105660 $Y=42400
X2393 1 DigitalLDOLogic_VIA0 $T=105910 48080 0 0 $X=105660 $Y=47840
X2394 1 DigitalLDOLogic_VIA0 $T=105910 53520 0 0 $X=105660 $Y=53280
X2395 1 DigitalLDOLogic_VIA0 $T=105910 58960 0 0 $X=105660 $Y=58720
X2396 3 DigitalLDOLogic_VIA0 $T=107750 12720 0 0 $X=107500 $Y=12480
X2397 3 DigitalLDOLogic_VIA0 $T=107750 18160 0 0 $X=107500 $Y=17920
X2398 3 DigitalLDOLogic_VIA0 $T=107750 23600 0 0 $X=107500 $Y=23360
X2399 3 DigitalLDOLogic_VIA0 $T=107750 29040 0 0 $X=107500 $Y=28800
X2400 3 DigitalLDOLogic_VIA0 $T=107750 34480 0 0 $X=107500 $Y=34240
X2401 3 DigitalLDOLogic_VIA0 $T=107750 39920 0 0 $X=107500 $Y=39680
X2402 3 DigitalLDOLogic_VIA0 $T=107750 45360 0 0 $X=107500 $Y=45120
X2403 3 DigitalLDOLogic_VIA0 $T=107750 50800 0 0 $X=107500 $Y=50560
X2404 3 DigitalLDOLogic_VIA0 $T=107750 56240 0 0 $X=107500 $Y=56000
X2405 1 DigitalLDOLogic_VIA0 $T=108670 15440 0 0 $X=108420 $Y=15200
X2406 1 DigitalLDOLogic_VIA0 $T=108670 20880 0 0 $X=108420 $Y=20640
X2407 1 DigitalLDOLogic_VIA0 $T=108670 26320 0 0 $X=108420 $Y=26080
X2408 1 DigitalLDOLogic_VIA0 $T=108670 31760 0 0 $X=108420 $Y=31520
X2409 1 DigitalLDOLogic_VIA0 $T=108670 37200 0 0 $X=108420 $Y=36960
X2410 1 DigitalLDOLogic_VIA0 $T=108670 42640 0 0 $X=108420 $Y=42400
X2411 1 DigitalLDOLogic_VIA0 $T=108670 48080 0 0 $X=108420 $Y=47840
X2412 1 DigitalLDOLogic_VIA0 $T=108670 53520 0 0 $X=108420 $Y=53280
X2413 1 DigitalLDOLogic_VIA0 $T=108670 58960 0 0 $X=108420 $Y=58720
X2414 3 DigitalLDOLogic_VIA0 $T=110510 12720 0 0 $X=110260 $Y=12480
X2415 3 DigitalLDOLogic_VIA0 $T=110510 18160 0 0 $X=110260 $Y=17920
X2416 3 DigitalLDOLogic_VIA0 $T=110510 23600 0 0 $X=110260 $Y=23360
X2417 3 DigitalLDOLogic_VIA0 $T=110510 29040 0 0 $X=110260 $Y=28800
X2418 3 DigitalLDOLogic_VIA0 $T=110510 34480 0 0 $X=110260 $Y=34240
X2419 3 DigitalLDOLogic_VIA0 $T=110510 39920 0 0 $X=110260 $Y=39680
X2420 3 DigitalLDOLogic_VIA0 $T=110510 45360 0 0 $X=110260 $Y=45120
X2421 3 DigitalLDOLogic_VIA0 $T=110510 50800 0 0 $X=110260 $Y=50560
X2422 3 DigitalLDOLogic_VIA0 $T=110510 56240 0 0 $X=110260 $Y=56000
X2423 1 DigitalLDOLogic_VIA0 $T=111430 15440 0 0 $X=111180 $Y=15200
X2424 1 DigitalLDOLogic_VIA0 $T=111430 20880 0 0 $X=111180 $Y=20640
X2425 1 DigitalLDOLogic_VIA0 $T=111430 26320 0 0 $X=111180 $Y=26080
X2426 1 DigitalLDOLogic_VIA0 $T=111430 31760 0 0 $X=111180 $Y=31520
X2427 1 DigitalLDOLogic_VIA0 $T=111430 37200 0 0 $X=111180 $Y=36960
X2428 1 DigitalLDOLogic_VIA0 $T=111430 42640 0 0 $X=111180 $Y=42400
X2429 1 DigitalLDOLogic_VIA0 $T=111430 48080 0 0 $X=111180 $Y=47840
X2430 1 DigitalLDOLogic_VIA0 $T=111430 53520 0 0 $X=111180 $Y=53280
X2431 1 DigitalLDOLogic_VIA0 $T=111430 58960 0 0 $X=111180 $Y=58720
X2432 3 DigitalLDOLogic_VIA0 $T=113270 12720 0 0 $X=113020 $Y=12480
X2433 3 DigitalLDOLogic_VIA0 $T=113270 18160 0 0 $X=113020 $Y=17920
X2434 3 DigitalLDOLogic_VIA0 $T=113270 23600 0 0 $X=113020 $Y=23360
X2435 3 DigitalLDOLogic_VIA0 $T=113270 29040 0 0 $X=113020 $Y=28800
X2436 3 DigitalLDOLogic_VIA0 $T=113270 34480 0 0 $X=113020 $Y=34240
X2437 3 DigitalLDOLogic_VIA0 $T=113270 39920 0 0 $X=113020 $Y=39680
X2438 3 DigitalLDOLogic_VIA0 $T=113270 45360 0 0 $X=113020 $Y=45120
X2439 3 DigitalLDOLogic_VIA0 $T=113270 50800 0 0 $X=113020 $Y=50560
X2440 3 DigitalLDOLogic_VIA0 $T=113270 56240 0 0 $X=113020 $Y=56000
X2441 1 DigitalLDOLogic_VIA0 $T=114190 15440 0 0 $X=113940 $Y=15200
X2442 1 DigitalLDOLogic_VIA0 $T=114190 20880 0 0 $X=113940 $Y=20640
X2443 1 DigitalLDOLogic_VIA0 $T=114190 26320 0 0 $X=113940 $Y=26080
X2444 1 DigitalLDOLogic_VIA0 $T=114190 31760 0 0 $X=113940 $Y=31520
X2445 1 DigitalLDOLogic_VIA0 $T=114190 37200 0 0 $X=113940 $Y=36960
X2446 1 DigitalLDOLogic_VIA0 $T=114190 42640 0 0 $X=113940 $Y=42400
X2447 1 DigitalLDOLogic_VIA0 $T=114190 48080 0 0 $X=113940 $Y=47840
X2448 1 DigitalLDOLogic_VIA0 $T=114190 53520 0 0 $X=113940 $Y=53280
X2449 1 DigitalLDOLogic_VIA0 $T=114190 58960 0 0 $X=113940 $Y=58720
X2450 3 DigitalLDOLogic_VIA0 $T=116030 12720 0 0 $X=115780 $Y=12480
X2451 3 DigitalLDOLogic_VIA0 $T=116030 18160 0 0 $X=115780 $Y=17920
X2452 3 DigitalLDOLogic_VIA0 $T=116030 23600 0 0 $X=115780 $Y=23360
X2453 3 DigitalLDOLogic_VIA0 $T=116030 29040 0 0 $X=115780 $Y=28800
X2454 3 DigitalLDOLogic_VIA0 $T=116030 34480 0 0 $X=115780 $Y=34240
X2455 3 DigitalLDOLogic_VIA0 $T=116030 39920 0 0 $X=115780 $Y=39680
X2456 3 DigitalLDOLogic_VIA0 $T=116030 45360 0 0 $X=115780 $Y=45120
X2457 3 DigitalLDOLogic_VIA0 $T=116030 50800 0 0 $X=115780 $Y=50560
X2458 3 DigitalLDOLogic_VIA0 $T=116030 56240 0 0 $X=115780 $Y=56000
X2459 1 DigitalLDOLogic_VIA0 $T=116950 15440 0 0 $X=116700 $Y=15200
X2460 1 DigitalLDOLogic_VIA0 $T=116950 20880 0 0 $X=116700 $Y=20640
X2461 1 DigitalLDOLogic_VIA0 $T=116950 26320 0 0 $X=116700 $Y=26080
X2462 1 DigitalLDOLogic_VIA0 $T=116950 31760 0 0 $X=116700 $Y=31520
X2463 1 DigitalLDOLogic_VIA0 $T=116950 37200 0 0 $X=116700 $Y=36960
X2464 1 DigitalLDOLogic_VIA0 $T=116950 42640 0 0 $X=116700 $Y=42400
X2465 1 DigitalLDOLogic_VIA0 $T=116950 48080 0 0 $X=116700 $Y=47840
X2466 1 DigitalLDOLogic_VIA0 $T=116950 53520 0 0 $X=116700 $Y=53280
X2467 1 DigitalLDOLogic_VIA0 $T=116950 58960 0 0 $X=116700 $Y=58720
X2468 3 DigitalLDOLogic_VIA0 $T=118790 12720 0 0 $X=118540 $Y=12480
X2469 3 DigitalLDOLogic_VIA0 $T=118790 18160 0 0 $X=118540 $Y=17920
X2470 3 DigitalLDOLogic_VIA0 $T=118790 23600 0 0 $X=118540 $Y=23360
X2471 3 DigitalLDOLogic_VIA0 $T=118790 29040 0 0 $X=118540 $Y=28800
X2472 3 DigitalLDOLogic_VIA0 $T=118790 34480 0 0 $X=118540 $Y=34240
X2473 3 DigitalLDOLogic_VIA0 $T=118790 39920 0 0 $X=118540 $Y=39680
X2474 3 DigitalLDOLogic_VIA0 $T=118790 45360 0 0 $X=118540 $Y=45120
X2475 3 DigitalLDOLogic_VIA0 $T=118790 50800 0 0 $X=118540 $Y=50560
X2476 3 DigitalLDOLogic_VIA0 $T=118790 56240 0 0 $X=118540 $Y=56000
X2477 1 DigitalLDOLogic_VIA0 $T=119710 15440 0 0 $X=119460 $Y=15200
X2478 1 DigitalLDOLogic_VIA0 $T=119710 20880 0 0 $X=119460 $Y=20640
X2479 1 DigitalLDOLogic_VIA0 $T=119710 26320 0 0 $X=119460 $Y=26080
X2480 1 DigitalLDOLogic_VIA0 $T=119710 31760 0 0 $X=119460 $Y=31520
X2481 1 DigitalLDOLogic_VIA0 $T=119710 37200 0 0 $X=119460 $Y=36960
X2482 1 DigitalLDOLogic_VIA0 $T=119710 42640 0 0 $X=119460 $Y=42400
X2483 1 DigitalLDOLogic_VIA0 $T=119710 48080 0 0 $X=119460 $Y=47840
X2484 1 DigitalLDOLogic_VIA0 $T=119710 53520 0 0 $X=119460 $Y=53280
X2485 1 DigitalLDOLogic_VIA0 $T=119710 58960 0 0 $X=119460 $Y=58720
X2486 3 DigitalLDOLogic_VIA0 $T=121550 12720 0 0 $X=121300 $Y=12480
X2487 3 DigitalLDOLogic_VIA0 $T=121550 18160 0 0 $X=121300 $Y=17920
X2488 3 DigitalLDOLogic_VIA0 $T=121550 23600 0 0 $X=121300 $Y=23360
X2489 3 DigitalLDOLogic_VIA0 $T=121550 29040 0 0 $X=121300 $Y=28800
X2490 3 DigitalLDOLogic_VIA0 $T=121550 34480 0 0 $X=121300 $Y=34240
X2491 3 DigitalLDOLogic_VIA0 $T=121550 39920 0 0 $X=121300 $Y=39680
X2492 3 DigitalLDOLogic_VIA0 $T=121550 45360 0 0 $X=121300 $Y=45120
X2493 3 DigitalLDOLogic_VIA0 $T=121550 50800 0 0 $X=121300 $Y=50560
X2494 3 DigitalLDOLogic_VIA0 $T=121550 56240 0 0 $X=121300 $Y=56000
X2495 1 DigitalLDOLogic_VIA0 $T=122470 15440 0 0 $X=122220 $Y=15200
X2496 1 DigitalLDOLogic_VIA0 $T=122470 20880 0 0 $X=122220 $Y=20640
X2497 1 DigitalLDOLogic_VIA0 $T=122470 26320 0 0 $X=122220 $Y=26080
X2498 1 DigitalLDOLogic_VIA0 $T=122470 31760 0 0 $X=122220 $Y=31520
X2499 1 DigitalLDOLogic_VIA0 $T=122470 37200 0 0 $X=122220 $Y=36960
X2500 1 DigitalLDOLogic_VIA0 $T=122470 42640 0 0 $X=122220 $Y=42400
X2501 1 DigitalLDOLogic_VIA0 $T=122470 48080 0 0 $X=122220 $Y=47840
X2502 1 DigitalLDOLogic_VIA0 $T=122470 53520 0 0 $X=122220 $Y=53280
X2503 1 DigitalLDOLogic_VIA0 $T=122470 58960 0 0 $X=122220 $Y=58720
X2504 3 DigitalLDOLogic_VIA0 $T=124310 12720 0 0 $X=124060 $Y=12480
X2505 3 DigitalLDOLogic_VIA0 $T=124310 18160 0 0 $X=124060 $Y=17920
X2506 3 DigitalLDOLogic_VIA0 $T=124310 23600 0 0 $X=124060 $Y=23360
X2507 3 DigitalLDOLogic_VIA0 $T=124310 29040 0 0 $X=124060 $Y=28800
X2508 3 DigitalLDOLogic_VIA0 $T=124310 34480 0 0 $X=124060 $Y=34240
X2509 3 DigitalLDOLogic_VIA0 $T=124310 39920 0 0 $X=124060 $Y=39680
X2510 3 DigitalLDOLogic_VIA0 $T=124310 45360 0 0 $X=124060 $Y=45120
X2511 3 DigitalLDOLogic_VIA0 $T=124310 50800 0 0 $X=124060 $Y=50560
X2512 3 DigitalLDOLogic_VIA0 $T=124310 56240 0 0 $X=124060 $Y=56000
X2513 1 DigitalLDOLogic_VIA0 $T=125230 15440 0 0 $X=124980 $Y=15200
X2514 1 DigitalLDOLogic_VIA0 $T=125230 20880 0 0 $X=124980 $Y=20640
X2515 1 DigitalLDOLogic_VIA0 $T=125230 26320 0 0 $X=124980 $Y=26080
X2516 1 DigitalLDOLogic_VIA0 $T=125230 31760 0 0 $X=124980 $Y=31520
X2517 1 DigitalLDOLogic_VIA0 $T=125230 37200 0 0 $X=124980 $Y=36960
X2518 1 DigitalLDOLogic_VIA0 $T=125230 42640 0 0 $X=124980 $Y=42400
X2519 1 DigitalLDOLogic_VIA0 $T=125230 48080 0 0 $X=124980 $Y=47840
X2520 1 DigitalLDOLogic_VIA0 $T=125230 53520 0 0 $X=124980 $Y=53280
X2521 1 DigitalLDOLogic_VIA0 $T=125230 58960 0 0 $X=124980 $Y=58720
X2522 3 DigitalLDOLogic_VIA0 $T=127070 12720 0 0 $X=126820 $Y=12480
X2523 3 DigitalLDOLogic_VIA0 $T=127070 18160 0 0 $X=126820 $Y=17920
X2524 3 DigitalLDOLogic_VIA0 $T=127070 23600 0 0 $X=126820 $Y=23360
X2525 3 DigitalLDOLogic_VIA0 $T=127070 29040 0 0 $X=126820 $Y=28800
X2526 3 DigitalLDOLogic_VIA0 $T=127070 34480 0 0 $X=126820 $Y=34240
X2527 3 DigitalLDOLogic_VIA0 $T=127070 39920 0 0 $X=126820 $Y=39680
X2528 3 DigitalLDOLogic_VIA0 $T=127070 45360 0 0 $X=126820 $Y=45120
X2529 3 DigitalLDOLogic_VIA0 $T=127070 50800 0 0 $X=126820 $Y=50560
X2530 3 DigitalLDOLogic_VIA0 $T=127070 56240 0 0 $X=126820 $Y=56000
X2531 1 DigitalLDOLogic_VIA0 $T=127990 15440 0 0 $X=127740 $Y=15200
X2532 1 DigitalLDOLogic_VIA0 $T=127990 20880 0 0 $X=127740 $Y=20640
X2533 1 DigitalLDOLogic_VIA0 $T=127990 26320 0 0 $X=127740 $Y=26080
X2534 1 DigitalLDOLogic_VIA0 $T=127990 31760 0 0 $X=127740 $Y=31520
X2535 1 DigitalLDOLogic_VIA0 $T=127990 37200 0 0 $X=127740 $Y=36960
X2536 1 DigitalLDOLogic_VIA0 $T=127990 42640 0 0 $X=127740 $Y=42400
X2537 1 DigitalLDOLogic_VIA0 $T=127990 48080 0 0 $X=127740 $Y=47840
X2538 1 DigitalLDOLogic_VIA0 $T=127990 53520 0 0 $X=127740 $Y=53280
X2539 1 DigitalLDOLogic_VIA0 $T=127990 58960 0 0 $X=127740 $Y=58720
X2540 3 DigitalLDOLogic_VIA0 $T=129830 12720 0 0 $X=129580 $Y=12480
X2541 3 DigitalLDOLogic_VIA0 $T=129830 18160 0 0 $X=129580 $Y=17920
X2542 3 DigitalLDOLogic_VIA0 $T=129830 23600 0 0 $X=129580 $Y=23360
X2543 3 DigitalLDOLogic_VIA0 $T=129830 29040 0 0 $X=129580 $Y=28800
X2544 3 DigitalLDOLogic_VIA0 $T=129830 34480 0 0 $X=129580 $Y=34240
X2545 3 DigitalLDOLogic_VIA0 $T=129830 39920 0 0 $X=129580 $Y=39680
X2546 3 DigitalLDOLogic_VIA0 $T=129830 45360 0 0 $X=129580 $Y=45120
X2547 3 DigitalLDOLogic_VIA0 $T=129830 50800 0 0 $X=129580 $Y=50560
X2548 3 DigitalLDOLogic_VIA0 $T=129830 56240 0 0 $X=129580 $Y=56000
X2549 1 DigitalLDOLogic_VIA0 $T=130750 15440 0 0 $X=130500 $Y=15200
X2550 1 DigitalLDOLogic_VIA0 $T=130750 20880 0 0 $X=130500 $Y=20640
X2551 1 DigitalLDOLogic_VIA0 $T=130750 26320 0 0 $X=130500 $Y=26080
X2552 1 DigitalLDOLogic_VIA0 $T=130750 31760 0 0 $X=130500 $Y=31520
X2553 1 DigitalLDOLogic_VIA0 $T=130750 37200 0 0 $X=130500 $Y=36960
X2554 1 DigitalLDOLogic_VIA0 $T=130750 42640 0 0 $X=130500 $Y=42400
X2555 1 DigitalLDOLogic_VIA0 $T=130750 48080 0 0 $X=130500 $Y=47840
X2556 1 DigitalLDOLogic_VIA0 $T=130750 53520 0 0 $X=130500 $Y=53280
X2557 1 DigitalLDOLogic_VIA0 $T=130750 58960 0 0 $X=130500 $Y=58720
X2558 3 DigitalLDOLogic_VIA0 $T=132590 12720 0 0 $X=132340 $Y=12480
X2559 3 DigitalLDOLogic_VIA0 $T=132590 18160 0 0 $X=132340 $Y=17920
X2560 3 DigitalLDOLogic_VIA0 $T=132590 23600 0 0 $X=132340 $Y=23360
X2561 3 DigitalLDOLogic_VIA0 $T=132590 29040 0 0 $X=132340 $Y=28800
X2562 3 DigitalLDOLogic_VIA0 $T=132590 34480 0 0 $X=132340 $Y=34240
X2563 3 DigitalLDOLogic_VIA0 $T=132590 39920 0 0 $X=132340 $Y=39680
X2564 3 DigitalLDOLogic_VIA0 $T=132590 45360 0 0 $X=132340 $Y=45120
X2565 3 DigitalLDOLogic_VIA0 $T=132590 50800 0 0 $X=132340 $Y=50560
X2566 3 DigitalLDOLogic_VIA0 $T=132590 56240 0 0 $X=132340 $Y=56000
X2567 1 DigitalLDOLogic_VIA0 $T=133510 15440 0 0 $X=133260 $Y=15200
X2568 1 DigitalLDOLogic_VIA0 $T=133510 20880 0 0 $X=133260 $Y=20640
X2569 1 DigitalLDOLogic_VIA0 $T=133510 26320 0 0 $X=133260 $Y=26080
X2570 1 DigitalLDOLogic_VIA0 $T=133510 31760 0 0 $X=133260 $Y=31520
X2571 1 DigitalLDOLogic_VIA0 $T=133510 37200 0 0 $X=133260 $Y=36960
X2572 1 DigitalLDOLogic_VIA0 $T=133510 42640 0 0 $X=133260 $Y=42400
X2573 1 DigitalLDOLogic_VIA0 $T=133510 48080 0 0 $X=133260 $Y=47840
X2574 1 DigitalLDOLogic_VIA0 $T=133510 53520 0 0 $X=133260 $Y=53280
X2575 1 DigitalLDOLogic_VIA0 $T=133510 58960 0 0 $X=133260 $Y=58720
X2576 3 DigitalLDOLogic_VIA0 $T=135350 12720 0 0 $X=135100 $Y=12480
X2577 3 DigitalLDOLogic_VIA0 $T=135350 18160 0 0 $X=135100 $Y=17920
X2578 3 DigitalLDOLogic_VIA0 $T=135350 23600 0 0 $X=135100 $Y=23360
X2579 3 DigitalLDOLogic_VIA0 $T=135350 29040 0 0 $X=135100 $Y=28800
X2580 3 DigitalLDOLogic_VIA0 $T=135350 34480 0 0 $X=135100 $Y=34240
X2581 3 DigitalLDOLogic_VIA0 $T=135350 39920 0 0 $X=135100 $Y=39680
X2582 3 DigitalLDOLogic_VIA0 $T=135350 45360 0 0 $X=135100 $Y=45120
X2583 3 DigitalLDOLogic_VIA0 $T=135350 50800 0 0 $X=135100 $Y=50560
X2584 3 DigitalLDOLogic_VIA0 $T=135350 56240 0 0 $X=135100 $Y=56000
X2585 1 DigitalLDOLogic_VIA0 $T=136270 15440 0 0 $X=136020 $Y=15200
X2586 1 DigitalLDOLogic_VIA0 $T=136270 20880 0 0 $X=136020 $Y=20640
X2587 1 DigitalLDOLogic_VIA0 $T=136270 26320 0 0 $X=136020 $Y=26080
X2588 1 DigitalLDOLogic_VIA0 $T=136270 31760 0 0 $X=136020 $Y=31520
X2589 1 DigitalLDOLogic_VIA0 $T=136270 37200 0 0 $X=136020 $Y=36960
X2590 1 DigitalLDOLogic_VIA0 $T=136270 42640 0 0 $X=136020 $Y=42400
X2591 1 DigitalLDOLogic_VIA0 $T=136270 48080 0 0 $X=136020 $Y=47840
X2592 1 DigitalLDOLogic_VIA0 $T=136270 53520 0 0 $X=136020 $Y=53280
X2593 1 DigitalLDOLogic_VIA0 $T=136270 58960 0 0 $X=136020 $Y=58720
X2594 3 DigitalLDOLogic_VIA0 $T=138110 12720 0 0 $X=137860 $Y=12480
X2595 3 DigitalLDOLogic_VIA0 $T=138110 18160 0 0 $X=137860 $Y=17920
X2596 3 DigitalLDOLogic_VIA0 $T=138110 23600 0 0 $X=137860 $Y=23360
X2597 3 DigitalLDOLogic_VIA0 $T=138110 29040 0 0 $X=137860 $Y=28800
X2598 3 DigitalLDOLogic_VIA0 $T=138110 34480 0 0 $X=137860 $Y=34240
X2599 3 DigitalLDOLogic_VIA0 $T=138110 39920 0 0 $X=137860 $Y=39680
X2600 3 DigitalLDOLogic_VIA0 $T=138110 45360 0 0 $X=137860 $Y=45120
X2601 3 DigitalLDOLogic_VIA0 $T=138110 50800 0 0 $X=137860 $Y=50560
X2602 3 DigitalLDOLogic_VIA0 $T=138110 56240 0 0 $X=137860 $Y=56000
X2603 1 DigitalLDOLogic_VIA0 $T=139030 15440 0 0 $X=138780 $Y=15200
X2604 1 DigitalLDOLogic_VIA0 $T=139030 20880 0 0 $X=138780 $Y=20640
X2605 1 DigitalLDOLogic_VIA0 $T=139030 26320 0 0 $X=138780 $Y=26080
X2606 1 DigitalLDOLogic_VIA0 $T=139030 31760 0 0 $X=138780 $Y=31520
X2607 1 DigitalLDOLogic_VIA0 $T=139030 37200 0 0 $X=138780 $Y=36960
X2608 1 DigitalLDOLogic_VIA0 $T=139030 42640 0 0 $X=138780 $Y=42400
X2609 1 DigitalLDOLogic_VIA0 $T=139030 48080 0 0 $X=138780 $Y=47840
X2610 1 DigitalLDOLogic_VIA0 $T=139030 53520 0 0 $X=138780 $Y=53280
X2611 1 DigitalLDOLogic_VIA0 $T=139030 58960 0 0 $X=138780 $Y=58720
X2612 3 DigitalLDOLogic_VIA0 $T=140870 12720 0 0 $X=140620 $Y=12480
X2613 3 DigitalLDOLogic_VIA0 $T=140870 18160 0 0 $X=140620 $Y=17920
X2614 3 DigitalLDOLogic_VIA0 $T=140870 23600 0 0 $X=140620 $Y=23360
X2615 3 DigitalLDOLogic_VIA0 $T=140870 29040 0 0 $X=140620 $Y=28800
X2616 3 DigitalLDOLogic_VIA0 $T=140870 34480 0 0 $X=140620 $Y=34240
X2617 3 DigitalLDOLogic_VIA0 $T=140870 39920 0 0 $X=140620 $Y=39680
X2618 3 DigitalLDOLogic_VIA0 $T=140870 45360 0 0 $X=140620 $Y=45120
X2619 3 DigitalLDOLogic_VIA0 $T=140870 50800 0 0 $X=140620 $Y=50560
X2620 3 DigitalLDOLogic_VIA0 $T=140870 56240 0 0 $X=140620 $Y=56000
X2621 1 DigitalLDOLogic_VIA0 $T=141790 15440 0 0 $X=141540 $Y=15200
X2622 1 DigitalLDOLogic_VIA0 $T=141790 20880 0 0 $X=141540 $Y=20640
X2623 1 DigitalLDOLogic_VIA0 $T=141790 26320 0 0 $X=141540 $Y=26080
X2624 1 DigitalLDOLogic_VIA0 $T=141790 31760 0 0 $X=141540 $Y=31520
X2625 1 DigitalLDOLogic_VIA0 $T=141790 37200 0 0 $X=141540 $Y=36960
X2626 1 DigitalLDOLogic_VIA0 $T=141790 42640 0 0 $X=141540 $Y=42400
X2627 1 DigitalLDOLogic_VIA0 $T=141790 48080 0 0 $X=141540 $Y=47840
X2628 1 DigitalLDOLogic_VIA0 $T=141790 53520 0 0 $X=141540 $Y=53280
X2629 1 DigitalLDOLogic_VIA0 $T=141790 58960 0 0 $X=141540 $Y=58720
X2630 3 DigitalLDOLogic_VIA0 $T=143630 12720 0 0 $X=143380 $Y=12480
X2631 3 DigitalLDOLogic_VIA0 $T=143630 18160 0 0 $X=143380 $Y=17920
X2632 3 DigitalLDOLogic_VIA0 $T=143630 23600 0 0 $X=143380 $Y=23360
X2633 3 DigitalLDOLogic_VIA0 $T=143630 29040 0 0 $X=143380 $Y=28800
X2634 3 DigitalLDOLogic_VIA0 $T=143630 34480 0 0 $X=143380 $Y=34240
X2635 3 DigitalLDOLogic_VIA0 $T=143630 39920 0 0 $X=143380 $Y=39680
X2636 3 DigitalLDOLogic_VIA0 $T=143630 45360 0 0 $X=143380 $Y=45120
X2637 3 DigitalLDOLogic_VIA0 $T=143630 50800 0 0 $X=143380 $Y=50560
X2638 3 DigitalLDOLogic_VIA0 $T=143630 56240 0 0 $X=143380 $Y=56000
X2639 1 DigitalLDOLogic_VIA0 $T=144550 15440 0 0 $X=144300 $Y=15200
X2640 1 DigitalLDOLogic_VIA0 $T=144550 20880 0 0 $X=144300 $Y=20640
X2641 1 DigitalLDOLogic_VIA0 $T=144550 26320 0 0 $X=144300 $Y=26080
X2642 1 DigitalLDOLogic_VIA0 $T=144550 31760 0 0 $X=144300 $Y=31520
X2643 1 DigitalLDOLogic_VIA0 $T=144550 37200 0 0 $X=144300 $Y=36960
X2644 1 DigitalLDOLogic_VIA0 $T=144550 42640 0 0 $X=144300 $Y=42400
X2645 1 DigitalLDOLogic_VIA0 $T=144550 48080 0 0 $X=144300 $Y=47840
X2646 1 DigitalLDOLogic_VIA0 $T=144550 53520 0 0 $X=144300 $Y=53280
X2647 1 DigitalLDOLogic_VIA0 $T=144550 58960 0 0 $X=144300 $Y=58720
X2648 3 DigitalLDOLogic_VIA0 $T=146390 12720 0 0 $X=146140 $Y=12480
X2649 3 DigitalLDOLogic_VIA0 $T=146390 18160 0 0 $X=146140 $Y=17920
X2650 3 DigitalLDOLogic_VIA0 $T=146390 23600 0 0 $X=146140 $Y=23360
X2651 3 DigitalLDOLogic_VIA0 $T=146390 29040 0 0 $X=146140 $Y=28800
X2652 3 DigitalLDOLogic_VIA0 $T=146390 34480 0 0 $X=146140 $Y=34240
X2653 3 DigitalLDOLogic_VIA0 $T=146390 39920 0 0 $X=146140 $Y=39680
X2654 3 DigitalLDOLogic_VIA0 $T=146390 45360 0 0 $X=146140 $Y=45120
X2655 3 DigitalLDOLogic_VIA0 $T=146390 50800 0 0 $X=146140 $Y=50560
X2656 3 DigitalLDOLogic_VIA0 $T=146390 56240 0 0 $X=146140 $Y=56000
X2657 1 DigitalLDOLogic_VIA0 $T=147310 15440 0 0 $X=147060 $Y=15200
X2658 1 DigitalLDOLogic_VIA0 $T=147310 20880 0 0 $X=147060 $Y=20640
X2659 1 DigitalLDOLogic_VIA0 $T=147310 26320 0 0 $X=147060 $Y=26080
X2660 1 DigitalLDOLogic_VIA0 $T=147310 31760 0 0 $X=147060 $Y=31520
X2661 1 DigitalLDOLogic_VIA0 $T=147310 37200 0 0 $X=147060 $Y=36960
X2662 1 DigitalLDOLogic_VIA0 $T=147310 42640 0 0 $X=147060 $Y=42400
X2663 1 DigitalLDOLogic_VIA0 $T=147310 48080 0 0 $X=147060 $Y=47840
X2664 1 DigitalLDOLogic_VIA0 $T=147310 53520 0 0 $X=147060 $Y=53280
X2665 1 DigitalLDOLogic_VIA0 $T=147310 58960 0 0 $X=147060 $Y=58720
X2666 3 DigitalLDOLogic_VIA0 $T=149150 12720 0 0 $X=148900 $Y=12480
X2667 3 DigitalLDOLogic_VIA0 $T=149150 18160 0 0 $X=148900 $Y=17920
X2668 3 DigitalLDOLogic_VIA0 $T=149150 23600 0 0 $X=148900 $Y=23360
X2669 3 DigitalLDOLogic_VIA0 $T=149150 29040 0 0 $X=148900 $Y=28800
X2670 3 DigitalLDOLogic_VIA0 $T=149150 34480 0 0 $X=148900 $Y=34240
X2671 3 DigitalLDOLogic_VIA0 $T=149150 39920 0 0 $X=148900 $Y=39680
X2672 3 DigitalLDOLogic_VIA0 $T=149150 45360 0 0 $X=148900 $Y=45120
X2673 3 DigitalLDOLogic_VIA0 $T=149150 50800 0 0 $X=148900 $Y=50560
X2674 3 DigitalLDOLogic_VIA0 $T=149150 56240 0 0 $X=148900 $Y=56000
X2675 1 DigitalLDOLogic_VIA0 $T=150070 15440 0 0 $X=149820 $Y=15200
X2676 1 DigitalLDOLogic_VIA0 $T=150070 20880 0 0 $X=149820 $Y=20640
X2677 1 DigitalLDOLogic_VIA0 $T=150070 26320 0 0 $X=149820 $Y=26080
X2678 1 DigitalLDOLogic_VIA0 $T=150070 31760 0 0 $X=149820 $Y=31520
X2679 1 DigitalLDOLogic_VIA0 $T=150070 37200 0 0 $X=149820 $Y=36960
X2680 1 DigitalLDOLogic_VIA0 $T=150070 42640 0 0 $X=149820 $Y=42400
X2681 1 DigitalLDOLogic_VIA0 $T=150070 48080 0 0 $X=149820 $Y=47840
X2682 1 DigitalLDOLogic_VIA0 $T=150070 53520 0 0 $X=149820 $Y=53280
X2683 1 DigitalLDOLogic_VIA0 $T=150070 58960 0 0 $X=149820 $Y=58720
X2684 3 DigitalLDOLogic_VIA0 $T=151910 12720 0 0 $X=151660 $Y=12480
X2685 3 DigitalLDOLogic_VIA0 $T=151910 18160 0 0 $X=151660 $Y=17920
X2686 3 DigitalLDOLogic_VIA0 $T=151910 23600 0 0 $X=151660 $Y=23360
X2687 3 DigitalLDOLogic_VIA0 $T=151910 29040 0 0 $X=151660 $Y=28800
X2688 3 DigitalLDOLogic_VIA0 $T=151910 34480 0 0 $X=151660 $Y=34240
X2689 3 DigitalLDOLogic_VIA0 $T=151910 39920 0 0 $X=151660 $Y=39680
X2690 3 DigitalLDOLogic_VIA0 $T=151910 45360 0 0 $X=151660 $Y=45120
X2691 3 DigitalLDOLogic_VIA0 $T=151910 50800 0 0 $X=151660 $Y=50560
X2692 3 DigitalLDOLogic_VIA0 $T=151910 56240 0 0 $X=151660 $Y=56000
X2693 1 DigitalLDOLogic_VIA0 $T=152830 15440 0 0 $X=152580 $Y=15200
X2694 1 DigitalLDOLogic_VIA0 $T=152830 20880 0 0 $X=152580 $Y=20640
X2695 1 DigitalLDOLogic_VIA0 $T=152830 26320 0 0 $X=152580 $Y=26080
X2696 1 DigitalLDOLogic_VIA0 $T=152830 31760 0 0 $X=152580 $Y=31520
X2697 1 DigitalLDOLogic_VIA0 $T=152830 37200 0 0 $X=152580 $Y=36960
X2698 1 DigitalLDOLogic_VIA0 $T=152830 42640 0 0 $X=152580 $Y=42400
X2699 1 DigitalLDOLogic_VIA0 $T=152830 48080 0 0 $X=152580 $Y=47840
X2700 1 DigitalLDOLogic_VIA0 $T=152830 53520 0 0 $X=152580 $Y=53280
X2701 1 DigitalLDOLogic_VIA0 $T=152830 58960 0 0 $X=152580 $Y=58720
X2702 3 DigitalLDOLogic_VIA0 $T=154670 12720 0 0 $X=154420 $Y=12480
X2703 3 DigitalLDOLogic_VIA0 $T=154670 18160 0 0 $X=154420 $Y=17920
X2704 3 DigitalLDOLogic_VIA0 $T=154670 23600 0 0 $X=154420 $Y=23360
X2705 3 DigitalLDOLogic_VIA0 $T=154670 29040 0 0 $X=154420 $Y=28800
X2706 3 DigitalLDOLogic_VIA0 $T=154670 34480 0 0 $X=154420 $Y=34240
X2707 3 DigitalLDOLogic_VIA0 $T=154670 39920 0 0 $X=154420 $Y=39680
X2708 3 DigitalLDOLogic_VIA0 $T=154670 45360 0 0 $X=154420 $Y=45120
X2709 3 DigitalLDOLogic_VIA0 $T=154670 50800 0 0 $X=154420 $Y=50560
X2710 3 DigitalLDOLogic_VIA0 $T=154670 56240 0 0 $X=154420 $Y=56000
X2711 1 DigitalLDOLogic_VIA0 $T=155590 15440 0 0 $X=155340 $Y=15200
X2712 1 DigitalLDOLogic_VIA0 $T=155590 20880 0 0 $X=155340 $Y=20640
X2713 1 DigitalLDOLogic_VIA0 $T=155590 26320 0 0 $X=155340 $Y=26080
X2714 1 DigitalLDOLogic_VIA0 $T=155590 31760 0 0 $X=155340 $Y=31520
X2715 1 DigitalLDOLogic_VIA0 $T=155590 37200 0 0 $X=155340 $Y=36960
X2716 1 DigitalLDOLogic_VIA0 $T=155590 42640 0 0 $X=155340 $Y=42400
X2717 1 DigitalLDOLogic_VIA0 $T=155590 48080 0 0 $X=155340 $Y=47840
X2718 1 DigitalLDOLogic_VIA0 $T=155590 53520 0 0 $X=155340 $Y=53280
X2719 1 DigitalLDOLogic_VIA0 $T=155590 58960 0 0 $X=155340 $Y=58720
X2720 3 DigitalLDOLogic_VIA0 $T=157430 12720 0 0 $X=157180 $Y=12480
X2721 3 DigitalLDOLogic_VIA0 $T=157430 18160 0 0 $X=157180 $Y=17920
X2722 3 DigitalLDOLogic_VIA0 $T=157430 23600 0 0 $X=157180 $Y=23360
X2723 3 DigitalLDOLogic_VIA0 $T=157430 29040 0 0 $X=157180 $Y=28800
X2724 3 DigitalLDOLogic_VIA0 $T=157430 34480 0 0 $X=157180 $Y=34240
X2725 3 DigitalLDOLogic_VIA0 $T=157430 39920 0 0 $X=157180 $Y=39680
X2726 3 DigitalLDOLogic_VIA0 $T=157430 45360 0 0 $X=157180 $Y=45120
X2727 3 DigitalLDOLogic_VIA0 $T=157430 50800 0 0 $X=157180 $Y=50560
X2728 3 DigitalLDOLogic_VIA0 $T=157430 56240 0 0 $X=157180 $Y=56000
X2729 1 DigitalLDOLogic_VIA0 $T=158350 15440 0 0 $X=158100 $Y=15200
X2730 1 DigitalLDOLogic_VIA0 $T=158350 20880 0 0 $X=158100 $Y=20640
X2731 1 DigitalLDOLogic_VIA0 $T=158350 26320 0 0 $X=158100 $Y=26080
X2732 1 DigitalLDOLogic_VIA0 $T=158350 31760 0 0 $X=158100 $Y=31520
X2733 1 DigitalLDOLogic_VIA0 $T=158350 37200 0 0 $X=158100 $Y=36960
X2734 1 DigitalLDOLogic_VIA0 $T=158350 42640 0 0 $X=158100 $Y=42400
X2735 1 DigitalLDOLogic_VIA0 $T=158350 48080 0 0 $X=158100 $Y=47840
X2736 1 DigitalLDOLogic_VIA0 $T=158350 53520 0 0 $X=158100 $Y=53280
X2737 1 DigitalLDOLogic_VIA0 $T=158350 58960 0 0 $X=158100 $Y=58720
X2738 3 DigitalLDOLogic_VIA0 $T=160190 12720 0 0 $X=159940 $Y=12480
X2739 3 DigitalLDOLogic_VIA0 $T=160190 18160 0 0 $X=159940 $Y=17920
X2740 3 DigitalLDOLogic_VIA0 $T=160190 23600 0 0 $X=159940 $Y=23360
X2741 3 DigitalLDOLogic_VIA0 $T=160190 29040 0 0 $X=159940 $Y=28800
X2742 3 DigitalLDOLogic_VIA0 $T=160190 34480 0 0 $X=159940 $Y=34240
X2743 3 DigitalLDOLogic_VIA0 $T=160190 39920 0 0 $X=159940 $Y=39680
X2744 3 DigitalLDOLogic_VIA0 $T=160190 45360 0 0 $X=159940 $Y=45120
X2745 3 DigitalLDOLogic_VIA0 $T=160190 50800 0 0 $X=159940 $Y=50560
X2746 3 DigitalLDOLogic_VIA0 $T=160190 56240 0 0 $X=159940 $Y=56000
X2747 1 DigitalLDOLogic_VIA0 $T=161110 15440 0 0 $X=160860 $Y=15200
X2748 1 DigitalLDOLogic_VIA0 $T=161110 20880 0 0 $X=160860 $Y=20640
X2749 1 DigitalLDOLogic_VIA0 $T=161110 26320 0 0 $X=160860 $Y=26080
X2750 1 DigitalLDOLogic_VIA0 $T=161110 31760 0 0 $X=160860 $Y=31520
X2751 1 DigitalLDOLogic_VIA0 $T=161110 37200 0 0 $X=160860 $Y=36960
X2752 1 DigitalLDOLogic_VIA0 $T=161110 42640 0 0 $X=160860 $Y=42400
X2753 1 DigitalLDOLogic_VIA0 $T=161110 48080 0 0 $X=160860 $Y=47840
X2754 1 DigitalLDOLogic_VIA0 $T=161110 53520 0 0 $X=160860 $Y=53280
X2755 1 DigitalLDOLogic_VIA0 $T=161110 58960 0 0 $X=160860 $Y=58720
X2756 3 DigitalLDOLogic_VIA0 $T=162950 12720 0 0 $X=162700 $Y=12480
X2757 3 DigitalLDOLogic_VIA0 $T=162950 18160 0 0 $X=162700 $Y=17920
X2758 3 DigitalLDOLogic_VIA0 $T=162950 23600 0 0 $X=162700 $Y=23360
X2759 3 DigitalLDOLogic_VIA0 $T=162950 29040 0 0 $X=162700 $Y=28800
X2760 3 DigitalLDOLogic_VIA0 $T=162950 34480 0 0 $X=162700 $Y=34240
X2761 3 DigitalLDOLogic_VIA0 $T=162950 39920 0 0 $X=162700 $Y=39680
X2762 3 DigitalLDOLogic_VIA0 $T=162950 45360 0 0 $X=162700 $Y=45120
X2763 3 DigitalLDOLogic_VIA0 $T=162950 50800 0 0 $X=162700 $Y=50560
X2764 3 DigitalLDOLogic_VIA0 $T=162950 56240 0 0 $X=162700 $Y=56000
X2765 1 DigitalLDOLogic_VIA0 $T=163870 15440 0 0 $X=163620 $Y=15200
X2766 1 DigitalLDOLogic_VIA0 $T=163870 20880 0 0 $X=163620 $Y=20640
X2767 1 DigitalLDOLogic_VIA0 $T=163870 26320 0 0 $X=163620 $Y=26080
X2768 1 DigitalLDOLogic_VIA0 $T=163870 31760 0 0 $X=163620 $Y=31520
X2769 1 DigitalLDOLogic_VIA0 $T=163870 37200 0 0 $X=163620 $Y=36960
X2770 1 DigitalLDOLogic_VIA0 $T=163870 42640 0 0 $X=163620 $Y=42400
X2771 1 DigitalLDOLogic_VIA0 $T=163870 48080 0 0 $X=163620 $Y=47840
X2772 1 DigitalLDOLogic_VIA0 $T=163870 53520 0 0 $X=163620 $Y=53280
X2773 1 DigitalLDOLogic_VIA0 $T=163870 58960 0 0 $X=163620 $Y=58720
X2774 3 DigitalLDOLogic_VIA0 $T=165710 12720 0 0 $X=165460 $Y=12480
X2775 3 DigitalLDOLogic_VIA0 $T=165710 18160 0 0 $X=165460 $Y=17920
X2776 3 DigitalLDOLogic_VIA0 $T=165710 23600 0 0 $X=165460 $Y=23360
X2777 3 DigitalLDOLogic_VIA0 $T=165710 29040 0 0 $X=165460 $Y=28800
X2778 3 DigitalLDOLogic_VIA0 $T=165710 34480 0 0 $X=165460 $Y=34240
X2779 3 DigitalLDOLogic_VIA0 $T=165710 39920 0 0 $X=165460 $Y=39680
X2780 3 DigitalLDOLogic_VIA0 $T=165710 45360 0 0 $X=165460 $Y=45120
X2781 3 DigitalLDOLogic_VIA0 $T=165710 50800 0 0 $X=165460 $Y=50560
X2782 3 DigitalLDOLogic_VIA0 $T=165710 56240 0 0 $X=165460 $Y=56000
X2783 1 DigitalLDOLogic_VIA0 $T=166630 15440 0 0 $X=166380 $Y=15200
X2784 1 DigitalLDOLogic_VIA0 $T=166630 20880 0 0 $X=166380 $Y=20640
X2785 1 DigitalLDOLogic_VIA0 $T=166630 26320 0 0 $X=166380 $Y=26080
X2786 1 DigitalLDOLogic_VIA0 $T=166630 31760 0 0 $X=166380 $Y=31520
X2787 1 DigitalLDOLogic_VIA0 $T=166630 37200 0 0 $X=166380 $Y=36960
X2788 1 DigitalLDOLogic_VIA0 $T=166630 42640 0 0 $X=166380 $Y=42400
X2789 1 DigitalLDOLogic_VIA0 $T=166630 48080 0 0 $X=166380 $Y=47840
X2790 1 DigitalLDOLogic_VIA0 $T=166630 53520 0 0 $X=166380 $Y=53280
X2791 1 DigitalLDOLogic_VIA0 $T=166630 58960 0 0 $X=166380 $Y=58720
X2792 3 DigitalLDOLogic_VIA0 $T=168470 12720 0 0 $X=168220 $Y=12480
X2793 3 DigitalLDOLogic_VIA0 $T=168470 18160 0 0 $X=168220 $Y=17920
X2794 3 DigitalLDOLogic_VIA0 $T=168470 23600 0 0 $X=168220 $Y=23360
X2795 3 DigitalLDOLogic_VIA0 $T=168470 29040 0 0 $X=168220 $Y=28800
X2796 3 DigitalLDOLogic_VIA0 $T=168470 34480 0 0 $X=168220 $Y=34240
X2797 3 DigitalLDOLogic_VIA0 $T=168470 39920 0 0 $X=168220 $Y=39680
X2798 3 DigitalLDOLogic_VIA0 $T=168470 45360 0 0 $X=168220 $Y=45120
X2799 3 DigitalLDOLogic_VIA0 $T=168470 50800 0 0 $X=168220 $Y=50560
X2800 3 DigitalLDOLogic_VIA0 $T=168470 56240 0 0 $X=168220 $Y=56000
X2801 1 DigitalLDOLogic_VIA0 $T=169390 15440 0 0 $X=169140 $Y=15200
X2802 1 DigitalLDOLogic_VIA0 $T=169390 20880 0 0 $X=169140 $Y=20640
X2803 1 DigitalLDOLogic_VIA0 $T=169390 26320 0 0 $X=169140 $Y=26080
X2804 1 DigitalLDOLogic_VIA0 $T=169390 31760 0 0 $X=169140 $Y=31520
X2805 1 DigitalLDOLogic_VIA0 $T=169390 37200 0 0 $X=169140 $Y=36960
X2806 1 DigitalLDOLogic_VIA0 $T=169390 42640 0 0 $X=169140 $Y=42400
X2807 1 DigitalLDOLogic_VIA0 $T=169390 48080 0 0 $X=169140 $Y=47840
X2808 1 DigitalLDOLogic_VIA0 $T=169390 53520 0 0 $X=169140 $Y=53280
X2809 1 DigitalLDOLogic_VIA0 $T=169390 58960 0 0 $X=169140 $Y=58720
X2810 3 DigitalLDOLogic_VIA0 $T=171230 12720 0 0 $X=170980 $Y=12480
X2811 3 DigitalLDOLogic_VIA0 $T=171230 18160 0 0 $X=170980 $Y=17920
X2812 3 DigitalLDOLogic_VIA0 $T=171230 23600 0 0 $X=170980 $Y=23360
X2813 3 DigitalLDOLogic_VIA0 $T=171230 29040 0 0 $X=170980 $Y=28800
X2814 3 DigitalLDOLogic_VIA0 $T=171230 34480 0 0 $X=170980 $Y=34240
X2815 3 DigitalLDOLogic_VIA0 $T=171230 39920 0 0 $X=170980 $Y=39680
X2816 3 DigitalLDOLogic_VIA0 $T=171230 45360 0 0 $X=170980 $Y=45120
X2817 3 DigitalLDOLogic_VIA0 $T=171230 50800 0 0 $X=170980 $Y=50560
X2818 3 DigitalLDOLogic_VIA0 $T=171230 56240 0 0 $X=170980 $Y=56000
X2819 1 DigitalLDOLogic_VIA0 $T=172150 15440 0 0 $X=171900 $Y=15200
X2820 1 DigitalLDOLogic_VIA0 $T=172150 20880 0 0 $X=171900 $Y=20640
X2821 1 DigitalLDOLogic_VIA0 $T=172150 26320 0 0 $X=171900 $Y=26080
X2822 1 DigitalLDOLogic_VIA0 $T=172150 31760 0 0 $X=171900 $Y=31520
X2823 1 DigitalLDOLogic_VIA0 $T=172150 37200 0 0 $X=171900 $Y=36960
X2824 1 DigitalLDOLogic_VIA0 $T=172150 42640 0 0 $X=171900 $Y=42400
X2825 1 DigitalLDOLogic_VIA0 $T=172150 48080 0 0 $X=171900 $Y=47840
X2826 1 DigitalLDOLogic_VIA0 $T=172150 53520 0 0 $X=171900 $Y=53280
X2827 1 DigitalLDOLogic_VIA0 $T=172150 58960 0 0 $X=171900 $Y=58720
X2828 3 DigitalLDOLogic_VIA0 $T=173990 12720 0 0 $X=173740 $Y=12480
X2829 3 DigitalLDOLogic_VIA0 $T=173990 18160 0 0 $X=173740 $Y=17920
X2830 3 DigitalLDOLogic_VIA0 $T=173990 23600 0 0 $X=173740 $Y=23360
X2831 3 DigitalLDOLogic_VIA0 $T=173990 29040 0 0 $X=173740 $Y=28800
X2832 3 DigitalLDOLogic_VIA0 $T=173990 34480 0 0 $X=173740 $Y=34240
X2833 3 DigitalLDOLogic_VIA0 $T=173990 39920 0 0 $X=173740 $Y=39680
X2834 3 DigitalLDOLogic_VIA0 $T=173990 45360 0 0 $X=173740 $Y=45120
X2835 3 DigitalLDOLogic_VIA0 $T=173990 50800 0 0 $X=173740 $Y=50560
X2836 3 DigitalLDOLogic_VIA0 $T=173990 56240 0 0 $X=173740 $Y=56000
X2837 1 DigitalLDOLogic_VIA0 $T=174910 15440 0 0 $X=174660 $Y=15200
X2838 1 DigitalLDOLogic_VIA0 $T=174910 20880 0 0 $X=174660 $Y=20640
X2839 1 DigitalLDOLogic_VIA0 $T=174910 26320 0 0 $X=174660 $Y=26080
X2840 1 DigitalLDOLogic_VIA0 $T=174910 31760 0 0 $X=174660 $Y=31520
X2841 1 DigitalLDOLogic_VIA0 $T=174910 37200 0 0 $X=174660 $Y=36960
X2842 1 DigitalLDOLogic_VIA0 $T=174910 42640 0 0 $X=174660 $Y=42400
X2843 1 DigitalLDOLogic_VIA0 $T=174910 48080 0 0 $X=174660 $Y=47840
X2844 1 DigitalLDOLogic_VIA0 $T=174910 53520 0 0 $X=174660 $Y=53280
X2845 1 DigitalLDOLogic_VIA0 $T=174910 58960 0 0 $X=174660 $Y=58720
X2846 3 DigitalLDOLogic_VIA0 $T=176750 12720 0 0 $X=176500 $Y=12480
X2847 3 DigitalLDOLogic_VIA0 $T=176750 18160 0 0 $X=176500 $Y=17920
X2848 3 DigitalLDOLogic_VIA0 $T=176750 23600 0 0 $X=176500 $Y=23360
X2849 3 DigitalLDOLogic_VIA0 $T=176750 29040 0 0 $X=176500 $Y=28800
X2850 3 DigitalLDOLogic_VIA0 $T=176750 34480 0 0 $X=176500 $Y=34240
X2851 3 DigitalLDOLogic_VIA0 $T=176750 39920 0 0 $X=176500 $Y=39680
X2852 3 DigitalLDOLogic_VIA0 $T=176750 45360 0 0 $X=176500 $Y=45120
X2853 3 DigitalLDOLogic_VIA0 $T=176750 50800 0 0 $X=176500 $Y=50560
X2854 3 DigitalLDOLogic_VIA0 $T=176750 56240 0 0 $X=176500 $Y=56000
X2855 1 DigitalLDOLogic_VIA0 $T=177670 15440 0 0 $X=177420 $Y=15200
X2856 1 DigitalLDOLogic_VIA0 $T=177670 20880 0 0 $X=177420 $Y=20640
X2857 1 DigitalLDOLogic_VIA0 $T=177670 26320 0 0 $X=177420 $Y=26080
X2858 1 DigitalLDOLogic_VIA0 $T=177670 31760 0 0 $X=177420 $Y=31520
X2859 1 DigitalLDOLogic_VIA0 $T=177670 37200 0 0 $X=177420 $Y=36960
X2860 1 DigitalLDOLogic_VIA0 $T=177670 42640 0 0 $X=177420 $Y=42400
X2861 1 DigitalLDOLogic_VIA0 $T=177670 48080 0 0 $X=177420 $Y=47840
X2862 1 DigitalLDOLogic_VIA0 $T=177670 53520 0 0 $X=177420 $Y=53280
X2863 1 DigitalLDOLogic_VIA0 $T=177670 58960 0 0 $X=177420 $Y=58720
X2864 3 DigitalLDOLogic_VIA0 $T=179510 12720 0 0 $X=179260 $Y=12480
X2865 3 DigitalLDOLogic_VIA0 $T=179510 18160 0 0 $X=179260 $Y=17920
X2866 3 DigitalLDOLogic_VIA0 $T=179510 23600 0 0 $X=179260 $Y=23360
X2867 3 DigitalLDOLogic_VIA0 $T=179510 29040 0 0 $X=179260 $Y=28800
X2868 3 DigitalLDOLogic_VIA0 $T=179510 34480 0 0 $X=179260 $Y=34240
X2869 3 DigitalLDOLogic_VIA0 $T=179510 39920 0 0 $X=179260 $Y=39680
X2870 3 DigitalLDOLogic_VIA0 $T=179510 45360 0 0 $X=179260 $Y=45120
X2871 3 DigitalLDOLogic_VIA0 $T=179510 50800 0 0 $X=179260 $Y=50560
X2872 3 DigitalLDOLogic_VIA0 $T=179510 56240 0 0 $X=179260 $Y=56000
X2873 1 DigitalLDOLogic_VIA0 $T=180430 15440 0 0 $X=180180 $Y=15200
X2874 1 DigitalLDOLogic_VIA0 $T=180430 20880 0 0 $X=180180 $Y=20640
X2875 1 DigitalLDOLogic_VIA0 $T=180430 26320 0 0 $X=180180 $Y=26080
X2876 1 DigitalLDOLogic_VIA0 $T=180430 31760 0 0 $X=180180 $Y=31520
X2877 1 DigitalLDOLogic_VIA0 $T=180430 37200 0 0 $X=180180 $Y=36960
X2878 1 DigitalLDOLogic_VIA0 $T=180430 42640 0 0 $X=180180 $Y=42400
X2879 1 DigitalLDOLogic_VIA0 $T=180430 48080 0 0 $X=180180 $Y=47840
X2880 1 DigitalLDOLogic_VIA0 $T=180430 53520 0 0 $X=180180 $Y=53280
X2881 1 DigitalLDOLogic_VIA0 $T=180430 58960 0 0 $X=180180 $Y=58720
X2882 3 DigitalLDOLogic_VIA0 $T=182270 12720 0 0 $X=182020 $Y=12480
X2883 3 DigitalLDOLogic_VIA0 $T=182270 18160 0 0 $X=182020 $Y=17920
X2884 3 DigitalLDOLogic_VIA0 $T=182270 23600 0 0 $X=182020 $Y=23360
X2885 3 DigitalLDOLogic_VIA0 $T=182270 29040 0 0 $X=182020 $Y=28800
X2886 3 DigitalLDOLogic_VIA0 $T=182270 34480 0 0 $X=182020 $Y=34240
X2887 3 DigitalLDOLogic_VIA0 $T=182270 39920 0 0 $X=182020 $Y=39680
X2888 3 DigitalLDOLogic_VIA0 $T=182270 45360 0 0 $X=182020 $Y=45120
X2889 3 DigitalLDOLogic_VIA0 $T=182270 50800 0 0 $X=182020 $Y=50560
X2890 3 DigitalLDOLogic_VIA0 $T=182270 56240 0 0 $X=182020 $Y=56000
X2891 1 DigitalLDOLogic_VIA0 $T=183190 15440 0 0 $X=182940 $Y=15200
X2892 1 DigitalLDOLogic_VIA0 $T=183190 20880 0 0 $X=182940 $Y=20640
X2893 1 DigitalLDOLogic_VIA0 $T=183190 26320 0 0 $X=182940 $Y=26080
X2894 1 DigitalLDOLogic_VIA0 $T=183190 31760 0 0 $X=182940 $Y=31520
X2895 1 DigitalLDOLogic_VIA0 $T=183190 37200 0 0 $X=182940 $Y=36960
X2896 1 DigitalLDOLogic_VIA0 $T=183190 42640 0 0 $X=182940 $Y=42400
X2897 1 DigitalLDOLogic_VIA0 $T=183190 48080 0 0 $X=182940 $Y=47840
X2898 1 DigitalLDOLogic_VIA0 $T=183190 53520 0 0 $X=182940 $Y=53280
X2899 1 DigitalLDOLogic_VIA0 $T=183190 58960 0 0 $X=182940 $Y=58720
X2900 3 DigitalLDOLogic_VIA0 $T=185030 12720 0 0 $X=184780 $Y=12480
X2901 3 DigitalLDOLogic_VIA0 $T=185030 18160 0 0 $X=184780 $Y=17920
X2902 3 DigitalLDOLogic_VIA0 $T=185030 23600 0 0 $X=184780 $Y=23360
X2903 3 DigitalLDOLogic_VIA0 $T=185030 29040 0 0 $X=184780 $Y=28800
X2904 3 DigitalLDOLogic_VIA0 $T=185030 34480 0 0 $X=184780 $Y=34240
X2905 3 DigitalLDOLogic_VIA0 $T=185030 39920 0 0 $X=184780 $Y=39680
X2906 3 DigitalLDOLogic_VIA0 $T=185030 45360 0 0 $X=184780 $Y=45120
X2907 3 DigitalLDOLogic_VIA0 $T=185030 50800 0 0 $X=184780 $Y=50560
X2908 3 DigitalLDOLogic_VIA0 $T=185030 56240 0 0 $X=184780 $Y=56000
X2909 1 DigitalLDOLogic_VIA0 $T=185950 15440 0 0 $X=185700 $Y=15200
X2910 1 DigitalLDOLogic_VIA0 $T=185950 20880 0 0 $X=185700 $Y=20640
X2911 1 DigitalLDOLogic_VIA0 $T=185950 26320 0 0 $X=185700 $Y=26080
X2912 1 DigitalLDOLogic_VIA0 $T=185950 31760 0 0 $X=185700 $Y=31520
X2913 1 DigitalLDOLogic_VIA0 $T=185950 37200 0 0 $X=185700 $Y=36960
X2914 1 DigitalLDOLogic_VIA0 $T=185950 42640 0 0 $X=185700 $Y=42400
X2915 1 DigitalLDOLogic_VIA0 $T=185950 48080 0 0 $X=185700 $Y=47840
X2916 1 DigitalLDOLogic_VIA0 $T=185950 53520 0 0 $X=185700 $Y=53280
X2917 1 DigitalLDOLogic_VIA0 $T=185950 58960 0 0 $X=185700 $Y=58720
X2918 3 DigitalLDOLogic_VIA0 $T=187790 12720 0 0 $X=187540 $Y=12480
X2919 3 DigitalLDOLogic_VIA0 $T=187790 18160 0 0 $X=187540 $Y=17920
X2920 3 DigitalLDOLogic_VIA0 $T=187790 23600 0 0 $X=187540 $Y=23360
X2921 3 DigitalLDOLogic_VIA0 $T=187790 29040 0 0 $X=187540 $Y=28800
X2922 3 DigitalLDOLogic_VIA0 $T=187790 34480 0 0 $X=187540 $Y=34240
X2923 3 DigitalLDOLogic_VIA0 $T=187790 39920 0 0 $X=187540 $Y=39680
X2924 3 DigitalLDOLogic_VIA0 $T=187790 45360 0 0 $X=187540 $Y=45120
X2925 3 DigitalLDOLogic_VIA0 $T=187790 50800 0 0 $X=187540 $Y=50560
X2926 3 DigitalLDOLogic_VIA0 $T=187790 56240 0 0 $X=187540 $Y=56000
X2927 1 DigitalLDOLogic_VIA0 $T=188710 15440 0 0 $X=188460 $Y=15200
X2928 1 DigitalLDOLogic_VIA0 $T=188710 20880 0 0 $X=188460 $Y=20640
X2929 1 DigitalLDOLogic_VIA0 $T=188710 26320 0 0 $X=188460 $Y=26080
X2930 1 DigitalLDOLogic_VIA0 $T=188710 31760 0 0 $X=188460 $Y=31520
X2931 1 DigitalLDOLogic_VIA0 $T=188710 37200 0 0 $X=188460 $Y=36960
X2932 1 DigitalLDOLogic_VIA0 $T=188710 42640 0 0 $X=188460 $Y=42400
X2933 1 DigitalLDOLogic_VIA0 $T=188710 48080 0 0 $X=188460 $Y=47840
X2934 1 DigitalLDOLogic_VIA0 $T=188710 53520 0 0 $X=188460 $Y=53280
X2935 1 DigitalLDOLogic_VIA0 $T=188710 58960 0 0 $X=188460 $Y=58720
X2936 3 DigitalLDOLogic_VIA1 $T=11150 11700 0 0 $X=10900 $Y=11470
X2937 3 DigitalLDOLogic_VIA1 $T=11150 15780 0 0 $X=10900 $Y=15550
X2938 3 DigitalLDOLogic_VIA1 $T=11150 19860 0 0 $X=10900 $Y=19630
X2939 3 DigitalLDOLogic_VIA1 $T=11150 23940 0 0 $X=10900 $Y=23710
X2940 3 DigitalLDOLogic_VIA1 $T=11150 28020 0 0 $X=10900 $Y=27790
X2941 3 DigitalLDOLogic_VIA1 $T=11150 32100 0 0 $X=10900 $Y=31870
X2942 3 DigitalLDOLogic_VIA1 $T=11150 36180 0 0 $X=10900 $Y=35950
X2943 3 DigitalLDOLogic_VIA1 $T=11150 40260 0 0 $X=10900 $Y=40030
X2944 3 DigitalLDOLogic_VIA1 $T=11150 44340 0 0 $X=10900 $Y=44110
X2945 3 DigitalLDOLogic_VIA1 $T=11150 48420 0 0 $X=10900 $Y=48190
X2946 3 DigitalLDOLogic_VIA1 $T=11150 52500 0 0 $X=10900 $Y=52270
X2947 3 DigitalLDOLogic_VIA1 $T=11150 56580 0 0 $X=10900 $Y=56350
X2948 1 DigitalLDOLogic_VIA1 $T=12070 13060 0 0 $X=11820 $Y=12830
X2949 1 DigitalLDOLogic_VIA1 $T=12070 17140 0 0 $X=11820 $Y=16910
X2950 1 DigitalLDOLogic_VIA1 $T=12070 21220 0 0 $X=11820 $Y=20990
X2951 1 DigitalLDOLogic_VIA1 $T=12070 25300 0 0 $X=11820 $Y=25070
X2952 1 DigitalLDOLogic_VIA1 $T=12070 29380 0 0 $X=11820 $Y=29150
X2953 1 DigitalLDOLogic_VIA1 $T=12070 33460 0 0 $X=11820 $Y=33230
X2954 1 DigitalLDOLogic_VIA1 $T=12070 37540 0 0 $X=11820 $Y=37310
X2955 1 DigitalLDOLogic_VIA1 $T=12070 41620 0 0 $X=11820 $Y=41390
X2956 1 DigitalLDOLogic_VIA1 $T=12070 45700 0 0 $X=11820 $Y=45470
X2957 1 DigitalLDOLogic_VIA1 $T=12070 49780 0 0 $X=11820 $Y=49550
X2958 1 DigitalLDOLogic_VIA1 $T=12070 53860 0 0 $X=11820 $Y=53630
X2959 1 DigitalLDOLogic_VIA1 $T=12070 57940 0 0 $X=11820 $Y=57710
X2960 3 DigitalLDOLogic_VIA1 $T=13910 11700 0 0 $X=13660 $Y=11470
X2961 3 DigitalLDOLogic_VIA1 $T=13910 15780 0 0 $X=13660 $Y=15550
X2962 3 DigitalLDOLogic_VIA1 $T=13910 19860 0 0 $X=13660 $Y=19630
X2963 3 DigitalLDOLogic_VIA1 $T=13910 23940 0 0 $X=13660 $Y=23710
X2964 3 DigitalLDOLogic_VIA1 $T=13910 28020 0 0 $X=13660 $Y=27790
X2965 3 DigitalLDOLogic_VIA1 $T=13910 32100 0 0 $X=13660 $Y=31870
X2966 3 DigitalLDOLogic_VIA1 $T=13910 36180 0 0 $X=13660 $Y=35950
X2967 3 DigitalLDOLogic_VIA1 $T=13910 40260 0 0 $X=13660 $Y=40030
X2968 3 DigitalLDOLogic_VIA1 $T=13910 44340 0 0 $X=13660 $Y=44110
X2969 3 DigitalLDOLogic_VIA1 $T=13910 48420 0 0 $X=13660 $Y=48190
X2970 3 DigitalLDOLogic_VIA1 $T=13910 52500 0 0 $X=13660 $Y=52270
X2971 3 DigitalLDOLogic_VIA1 $T=13910 56580 0 0 $X=13660 $Y=56350
X2972 1 DigitalLDOLogic_VIA1 $T=14830 13060 0 0 $X=14580 $Y=12830
X2973 1 DigitalLDOLogic_VIA1 $T=14830 17140 0 0 $X=14580 $Y=16910
X2974 1 DigitalLDOLogic_VIA1 $T=14830 21220 0 0 $X=14580 $Y=20990
X2975 1 DigitalLDOLogic_VIA1 $T=14830 25300 0 0 $X=14580 $Y=25070
X2976 1 DigitalLDOLogic_VIA1 $T=14830 29380 0 0 $X=14580 $Y=29150
X2977 1 DigitalLDOLogic_VIA1 $T=14830 33460 0 0 $X=14580 $Y=33230
X2978 1 DigitalLDOLogic_VIA1 $T=14830 37540 0 0 $X=14580 $Y=37310
X2979 1 DigitalLDOLogic_VIA1 $T=14830 41620 0 0 $X=14580 $Y=41390
X2980 1 DigitalLDOLogic_VIA1 $T=14830 45700 0 0 $X=14580 $Y=45470
X2981 1 DigitalLDOLogic_VIA1 $T=14830 49780 0 0 $X=14580 $Y=49550
X2982 1 DigitalLDOLogic_VIA1 $T=14830 53860 0 0 $X=14580 $Y=53630
X2983 1 DigitalLDOLogic_VIA1 $T=14830 57940 0 0 $X=14580 $Y=57710
X2984 3 DigitalLDOLogic_VIA1 $T=16670 11700 0 0 $X=16420 $Y=11470
X2985 3 DigitalLDOLogic_VIA1 $T=16670 15780 0 0 $X=16420 $Y=15550
X2986 3 DigitalLDOLogic_VIA1 $T=16670 19860 0 0 $X=16420 $Y=19630
X2987 3 DigitalLDOLogic_VIA1 $T=16670 23940 0 0 $X=16420 $Y=23710
X2988 3 DigitalLDOLogic_VIA1 $T=16670 28020 0 0 $X=16420 $Y=27790
X2989 3 DigitalLDOLogic_VIA1 $T=16670 32100 0 0 $X=16420 $Y=31870
X2990 3 DigitalLDOLogic_VIA1 $T=16670 36180 0 0 $X=16420 $Y=35950
X2991 3 DigitalLDOLogic_VIA1 $T=16670 40260 0 0 $X=16420 $Y=40030
X2992 3 DigitalLDOLogic_VIA1 $T=16670 44340 0 0 $X=16420 $Y=44110
X2993 3 DigitalLDOLogic_VIA1 $T=16670 48420 0 0 $X=16420 $Y=48190
X2994 3 DigitalLDOLogic_VIA1 $T=16670 52500 0 0 $X=16420 $Y=52270
X2995 3 DigitalLDOLogic_VIA1 $T=16670 56580 0 0 $X=16420 $Y=56350
X2996 1 DigitalLDOLogic_VIA1 $T=17590 13060 0 0 $X=17340 $Y=12830
X2997 1 DigitalLDOLogic_VIA1 $T=17590 17140 0 0 $X=17340 $Y=16910
X2998 1 DigitalLDOLogic_VIA1 $T=17590 21220 0 0 $X=17340 $Y=20990
X2999 1 DigitalLDOLogic_VIA1 $T=17590 25300 0 0 $X=17340 $Y=25070
X3000 1 DigitalLDOLogic_VIA1 $T=17590 29380 0 0 $X=17340 $Y=29150
X3001 1 DigitalLDOLogic_VIA1 $T=17590 33460 0 0 $X=17340 $Y=33230
X3002 1 DigitalLDOLogic_VIA1 $T=17590 37540 0 0 $X=17340 $Y=37310
X3003 1 DigitalLDOLogic_VIA1 $T=17590 41620 0 0 $X=17340 $Y=41390
X3004 1 DigitalLDOLogic_VIA1 $T=17590 45700 0 0 $X=17340 $Y=45470
X3005 1 DigitalLDOLogic_VIA1 $T=17590 49780 0 0 $X=17340 $Y=49550
X3006 1 DigitalLDOLogic_VIA1 $T=17590 53860 0 0 $X=17340 $Y=53630
X3007 1 DigitalLDOLogic_VIA1 $T=17590 57940 0 0 $X=17340 $Y=57710
X3008 3 DigitalLDOLogic_VIA1 $T=19430 11700 0 0 $X=19180 $Y=11470
X3009 3 DigitalLDOLogic_VIA1 $T=19430 15780 0 0 $X=19180 $Y=15550
X3010 3 DigitalLDOLogic_VIA1 $T=19430 19860 0 0 $X=19180 $Y=19630
X3011 3 DigitalLDOLogic_VIA1 $T=19430 23940 0 0 $X=19180 $Y=23710
X3012 3 DigitalLDOLogic_VIA1 $T=19430 28020 0 0 $X=19180 $Y=27790
X3013 3 DigitalLDOLogic_VIA1 $T=19430 32100 0 0 $X=19180 $Y=31870
X3014 3 DigitalLDOLogic_VIA1 $T=19430 36180 0 0 $X=19180 $Y=35950
X3015 3 DigitalLDOLogic_VIA1 $T=19430 40260 0 0 $X=19180 $Y=40030
X3016 3 DigitalLDOLogic_VIA1 $T=19430 44340 0 0 $X=19180 $Y=44110
X3017 3 DigitalLDOLogic_VIA1 $T=19430 48420 0 0 $X=19180 $Y=48190
X3018 3 DigitalLDOLogic_VIA1 $T=19430 52500 0 0 $X=19180 $Y=52270
X3019 3 DigitalLDOLogic_VIA1 $T=19430 56580 0 0 $X=19180 $Y=56350
X3020 1 DigitalLDOLogic_VIA1 $T=20350 13060 0 0 $X=20100 $Y=12830
X3021 1 DigitalLDOLogic_VIA1 $T=20350 17140 0 0 $X=20100 $Y=16910
X3022 1 DigitalLDOLogic_VIA1 $T=20350 21220 0 0 $X=20100 $Y=20990
X3023 1 DigitalLDOLogic_VIA1 $T=20350 25300 0 0 $X=20100 $Y=25070
X3024 1 DigitalLDOLogic_VIA1 $T=20350 29380 0 0 $X=20100 $Y=29150
X3025 1 DigitalLDOLogic_VIA1 $T=20350 33460 0 0 $X=20100 $Y=33230
X3026 1 DigitalLDOLogic_VIA1 $T=20350 37540 0 0 $X=20100 $Y=37310
X3027 1 DigitalLDOLogic_VIA1 $T=20350 41620 0 0 $X=20100 $Y=41390
X3028 1 DigitalLDOLogic_VIA1 $T=20350 45700 0 0 $X=20100 $Y=45470
X3029 1 DigitalLDOLogic_VIA1 $T=20350 49780 0 0 $X=20100 $Y=49550
X3030 1 DigitalLDOLogic_VIA1 $T=20350 53860 0 0 $X=20100 $Y=53630
X3031 1 DigitalLDOLogic_VIA1 $T=20350 57940 0 0 $X=20100 $Y=57710
X3032 3 DigitalLDOLogic_VIA1 $T=22190 11700 0 0 $X=21940 $Y=11470
X3033 3 DigitalLDOLogic_VIA1 $T=22190 15780 0 0 $X=21940 $Y=15550
X3034 3 DigitalLDOLogic_VIA1 $T=22190 19860 0 0 $X=21940 $Y=19630
X3035 3 DigitalLDOLogic_VIA1 $T=22190 23940 0 0 $X=21940 $Y=23710
X3036 3 DigitalLDOLogic_VIA1 $T=22190 28020 0 0 $X=21940 $Y=27790
X3037 3 DigitalLDOLogic_VIA1 $T=22190 32100 0 0 $X=21940 $Y=31870
X3038 3 DigitalLDOLogic_VIA1 $T=22190 36180 0 0 $X=21940 $Y=35950
X3039 3 DigitalLDOLogic_VIA1 $T=22190 40260 0 0 $X=21940 $Y=40030
X3040 3 DigitalLDOLogic_VIA1 $T=22190 44340 0 0 $X=21940 $Y=44110
X3041 3 DigitalLDOLogic_VIA1 $T=22190 48420 0 0 $X=21940 $Y=48190
X3042 3 DigitalLDOLogic_VIA1 $T=22190 52500 0 0 $X=21940 $Y=52270
X3043 3 DigitalLDOLogic_VIA1 $T=22190 56580 0 0 $X=21940 $Y=56350
X3044 1 DigitalLDOLogic_VIA1 $T=23110 13060 0 0 $X=22860 $Y=12830
X3045 1 DigitalLDOLogic_VIA1 $T=23110 17140 0 0 $X=22860 $Y=16910
X3046 1 DigitalLDOLogic_VIA1 $T=23110 21220 0 0 $X=22860 $Y=20990
X3047 1 DigitalLDOLogic_VIA1 $T=23110 25300 0 0 $X=22860 $Y=25070
X3048 1 DigitalLDOLogic_VIA1 $T=23110 29380 0 0 $X=22860 $Y=29150
X3049 1 DigitalLDOLogic_VIA1 $T=23110 33460 0 0 $X=22860 $Y=33230
X3050 1 DigitalLDOLogic_VIA1 $T=23110 37540 0 0 $X=22860 $Y=37310
X3051 1 DigitalLDOLogic_VIA1 $T=23110 41620 0 0 $X=22860 $Y=41390
X3052 1 DigitalLDOLogic_VIA1 $T=23110 45700 0 0 $X=22860 $Y=45470
X3053 1 DigitalLDOLogic_VIA1 $T=23110 49780 0 0 $X=22860 $Y=49550
X3054 1 DigitalLDOLogic_VIA1 $T=23110 53860 0 0 $X=22860 $Y=53630
X3055 1 DigitalLDOLogic_VIA1 $T=23110 57940 0 0 $X=22860 $Y=57710
X3056 3 DigitalLDOLogic_VIA1 $T=24950 11700 0 0 $X=24700 $Y=11470
X3057 3 DigitalLDOLogic_VIA1 $T=24950 15780 0 0 $X=24700 $Y=15550
X3058 3 DigitalLDOLogic_VIA1 $T=24950 19860 0 0 $X=24700 $Y=19630
X3059 3 DigitalLDOLogic_VIA1 $T=24950 23940 0 0 $X=24700 $Y=23710
X3060 3 DigitalLDOLogic_VIA1 $T=24950 28020 0 0 $X=24700 $Y=27790
X3061 3 DigitalLDOLogic_VIA1 $T=24950 32100 0 0 $X=24700 $Y=31870
X3062 3 DigitalLDOLogic_VIA1 $T=24950 36180 0 0 $X=24700 $Y=35950
X3063 3 DigitalLDOLogic_VIA1 $T=24950 40260 0 0 $X=24700 $Y=40030
X3064 3 DigitalLDOLogic_VIA1 $T=24950 44340 0 0 $X=24700 $Y=44110
X3065 3 DigitalLDOLogic_VIA1 $T=24950 48420 0 0 $X=24700 $Y=48190
X3066 3 DigitalLDOLogic_VIA1 $T=24950 52500 0 0 $X=24700 $Y=52270
X3067 3 DigitalLDOLogic_VIA1 $T=24950 56580 0 0 $X=24700 $Y=56350
X3068 1 DigitalLDOLogic_VIA1 $T=25870 13060 0 0 $X=25620 $Y=12830
X3069 1 DigitalLDOLogic_VIA1 $T=25870 17140 0 0 $X=25620 $Y=16910
X3070 1 DigitalLDOLogic_VIA1 $T=25870 21220 0 0 $X=25620 $Y=20990
X3071 1 DigitalLDOLogic_VIA1 $T=25870 25300 0 0 $X=25620 $Y=25070
X3072 1 DigitalLDOLogic_VIA1 $T=25870 29380 0 0 $X=25620 $Y=29150
X3073 1 DigitalLDOLogic_VIA1 $T=25870 33460 0 0 $X=25620 $Y=33230
X3074 1 DigitalLDOLogic_VIA1 $T=25870 37540 0 0 $X=25620 $Y=37310
X3075 1 DigitalLDOLogic_VIA1 $T=25870 41620 0 0 $X=25620 $Y=41390
X3076 1 DigitalLDOLogic_VIA1 $T=25870 45700 0 0 $X=25620 $Y=45470
X3077 1 DigitalLDOLogic_VIA1 $T=25870 49780 0 0 $X=25620 $Y=49550
X3078 1 DigitalLDOLogic_VIA1 $T=25870 53860 0 0 $X=25620 $Y=53630
X3079 1 DigitalLDOLogic_VIA1 $T=25870 57940 0 0 $X=25620 $Y=57710
X3080 3 DigitalLDOLogic_VIA1 $T=27710 11700 0 0 $X=27460 $Y=11470
X3081 3 DigitalLDOLogic_VIA1 $T=27710 15780 0 0 $X=27460 $Y=15550
X3082 3 DigitalLDOLogic_VIA1 $T=27710 19860 0 0 $X=27460 $Y=19630
X3083 3 DigitalLDOLogic_VIA1 $T=27710 23940 0 0 $X=27460 $Y=23710
X3084 3 DigitalLDOLogic_VIA1 $T=27710 28020 0 0 $X=27460 $Y=27790
X3085 3 DigitalLDOLogic_VIA1 $T=27710 32100 0 0 $X=27460 $Y=31870
X3086 3 DigitalLDOLogic_VIA1 $T=27710 36180 0 0 $X=27460 $Y=35950
X3087 3 DigitalLDOLogic_VIA1 $T=27710 40260 0 0 $X=27460 $Y=40030
X3088 3 DigitalLDOLogic_VIA1 $T=27710 44340 0 0 $X=27460 $Y=44110
X3089 3 DigitalLDOLogic_VIA1 $T=27710 48420 0 0 $X=27460 $Y=48190
X3090 3 DigitalLDOLogic_VIA1 $T=27710 52500 0 0 $X=27460 $Y=52270
X3091 3 DigitalLDOLogic_VIA1 $T=27710 56580 0 0 $X=27460 $Y=56350
X3092 1 DigitalLDOLogic_VIA1 $T=28630 13060 0 0 $X=28380 $Y=12830
X3093 1 DigitalLDOLogic_VIA1 $T=28630 17140 0 0 $X=28380 $Y=16910
X3094 1 DigitalLDOLogic_VIA1 $T=28630 21220 0 0 $X=28380 $Y=20990
X3095 1 DigitalLDOLogic_VIA1 $T=28630 25300 0 0 $X=28380 $Y=25070
X3096 1 DigitalLDOLogic_VIA1 $T=28630 29380 0 0 $X=28380 $Y=29150
X3097 1 DigitalLDOLogic_VIA1 $T=28630 33460 0 0 $X=28380 $Y=33230
X3098 1 DigitalLDOLogic_VIA1 $T=28630 37540 0 0 $X=28380 $Y=37310
X3099 1 DigitalLDOLogic_VIA1 $T=28630 41620 0 0 $X=28380 $Y=41390
X3100 1 DigitalLDOLogic_VIA1 $T=28630 45700 0 0 $X=28380 $Y=45470
X3101 1 DigitalLDOLogic_VIA1 $T=28630 49780 0 0 $X=28380 $Y=49550
X3102 1 DigitalLDOLogic_VIA1 $T=28630 53860 0 0 $X=28380 $Y=53630
X3103 1 DigitalLDOLogic_VIA1 $T=28630 57940 0 0 $X=28380 $Y=57710
X3104 3 DigitalLDOLogic_VIA1 $T=30470 11700 0 0 $X=30220 $Y=11470
X3105 3 DigitalLDOLogic_VIA1 $T=30470 15780 0 0 $X=30220 $Y=15550
X3106 3 DigitalLDOLogic_VIA1 $T=30470 19860 0 0 $X=30220 $Y=19630
X3107 3 DigitalLDOLogic_VIA1 $T=30470 23940 0 0 $X=30220 $Y=23710
X3108 3 DigitalLDOLogic_VIA1 $T=30470 28020 0 0 $X=30220 $Y=27790
X3109 3 DigitalLDOLogic_VIA1 $T=30470 32100 0 0 $X=30220 $Y=31870
X3110 3 DigitalLDOLogic_VIA1 $T=30470 36180 0 0 $X=30220 $Y=35950
X3111 3 DigitalLDOLogic_VIA1 $T=30470 40260 0 0 $X=30220 $Y=40030
X3112 3 DigitalLDOLogic_VIA1 $T=30470 44340 0 0 $X=30220 $Y=44110
X3113 3 DigitalLDOLogic_VIA1 $T=30470 48420 0 0 $X=30220 $Y=48190
X3114 3 DigitalLDOLogic_VIA1 $T=30470 52500 0 0 $X=30220 $Y=52270
X3115 3 DigitalLDOLogic_VIA1 $T=30470 56580 0 0 $X=30220 $Y=56350
X3116 1 DigitalLDOLogic_VIA1 $T=31390 13060 0 0 $X=31140 $Y=12830
X3117 1 DigitalLDOLogic_VIA1 $T=31390 17140 0 0 $X=31140 $Y=16910
X3118 1 DigitalLDOLogic_VIA1 $T=31390 21220 0 0 $X=31140 $Y=20990
X3119 1 DigitalLDOLogic_VIA1 $T=31390 25300 0 0 $X=31140 $Y=25070
X3120 1 DigitalLDOLogic_VIA1 $T=31390 29380 0 0 $X=31140 $Y=29150
X3121 1 DigitalLDOLogic_VIA1 $T=31390 33460 0 0 $X=31140 $Y=33230
X3122 1 DigitalLDOLogic_VIA1 $T=31390 37540 0 0 $X=31140 $Y=37310
X3123 1 DigitalLDOLogic_VIA1 $T=31390 41620 0 0 $X=31140 $Y=41390
X3124 1 DigitalLDOLogic_VIA1 $T=31390 45700 0 0 $X=31140 $Y=45470
X3125 1 DigitalLDOLogic_VIA1 $T=31390 49780 0 0 $X=31140 $Y=49550
X3126 1 DigitalLDOLogic_VIA1 $T=31390 53860 0 0 $X=31140 $Y=53630
X3127 1 DigitalLDOLogic_VIA1 $T=31390 57940 0 0 $X=31140 $Y=57710
X3128 3 DigitalLDOLogic_VIA1 $T=33230 11700 0 0 $X=32980 $Y=11470
X3129 3 DigitalLDOLogic_VIA1 $T=33230 15780 0 0 $X=32980 $Y=15550
X3130 3 DigitalLDOLogic_VIA1 $T=33230 19860 0 0 $X=32980 $Y=19630
X3131 3 DigitalLDOLogic_VIA1 $T=33230 23940 0 0 $X=32980 $Y=23710
X3132 3 DigitalLDOLogic_VIA1 $T=33230 28020 0 0 $X=32980 $Y=27790
X3133 3 DigitalLDOLogic_VIA1 $T=33230 32100 0 0 $X=32980 $Y=31870
X3134 3 DigitalLDOLogic_VIA1 $T=33230 36180 0 0 $X=32980 $Y=35950
X3135 3 DigitalLDOLogic_VIA1 $T=33230 40260 0 0 $X=32980 $Y=40030
X3136 3 DigitalLDOLogic_VIA1 $T=33230 44340 0 0 $X=32980 $Y=44110
X3137 3 DigitalLDOLogic_VIA1 $T=33230 48420 0 0 $X=32980 $Y=48190
X3138 3 DigitalLDOLogic_VIA1 $T=33230 52500 0 0 $X=32980 $Y=52270
X3139 3 DigitalLDOLogic_VIA1 $T=33230 56580 0 0 $X=32980 $Y=56350
X3140 1 DigitalLDOLogic_VIA1 $T=34150 13060 0 0 $X=33900 $Y=12830
X3141 1 DigitalLDOLogic_VIA1 $T=34150 17140 0 0 $X=33900 $Y=16910
X3142 1 DigitalLDOLogic_VIA1 $T=34150 21220 0 0 $X=33900 $Y=20990
X3143 1 DigitalLDOLogic_VIA1 $T=34150 25300 0 0 $X=33900 $Y=25070
X3144 1 DigitalLDOLogic_VIA1 $T=34150 29380 0 0 $X=33900 $Y=29150
X3145 1 DigitalLDOLogic_VIA1 $T=34150 33460 0 0 $X=33900 $Y=33230
X3146 1 DigitalLDOLogic_VIA1 $T=34150 37540 0 0 $X=33900 $Y=37310
X3147 1 DigitalLDOLogic_VIA1 $T=34150 41620 0 0 $X=33900 $Y=41390
X3148 1 DigitalLDOLogic_VIA1 $T=34150 45700 0 0 $X=33900 $Y=45470
X3149 1 DigitalLDOLogic_VIA1 $T=34150 49780 0 0 $X=33900 $Y=49550
X3150 1 DigitalLDOLogic_VIA1 $T=34150 53860 0 0 $X=33900 $Y=53630
X3151 1 DigitalLDOLogic_VIA1 $T=34150 57940 0 0 $X=33900 $Y=57710
X3152 3 DigitalLDOLogic_VIA1 $T=35990 11700 0 0 $X=35740 $Y=11470
X3153 3 DigitalLDOLogic_VIA1 $T=35990 15780 0 0 $X=35740 $Y=15550
X3154 3 DigitalLDOLogic_VIA1 $T=35990 19860 0 0 $X=35740 $Y=19630
X3155 3 DigitalLDOLogic_VIA1 $T=35990 23940 0 0 $X=35740 $Y=23710
X3156 3 DigitalLDOLogic_VIA1 $T=35990 28020 0 0 $X=35740 $Y=27790
X3157 3 DigitalLDOLogic_VIA1 $T=35990 32100 0 0 $X=35740 $Y=31870
X3158 3 DigitalLDOLogic_VIA1 $T=35990 36180 0 0 $X=35740 $Y=35950
X3159 3 DigitalLDOLogic_VIA1 $T=35990 40260 0 0 $X=35740 $Y=40030
X3160 3 DigitalLDOLogic_VIA1 $T=35990 44340 0 0 $X=35740 $Y=44110
X3161 3 DigitalLDOLogic_VIA1 $T=35990 48420 0 0 $X=35740 $Y=48190
X3162 3 DigitalLDOLogic_VIA1 $T=35990 52500 0 0 $X=35740 $Y=52270
X3163 3 DigitalLDOLogic_VIA1 $T=35990 56580 0 0 $X=35740 $Y=56350
X3164 1 DigitalLDOLogic_VIA1 $T=36910 13060 0 0 $X=36660 $Y=12830
X3165 1 DigitalLDOLogic_VIA1 $T=36910 17140 0 0 $X=36660 $Y=16910
X3166 1 DigitalLDOLogic_VIA1 $T=36910 21220 0 0 $X=36660 $Y=20990
X3167 1 DigitalLDOLogic_VIA1 $T=36910 25300 0 0 $X=36660 $Y=25070
X3168 1 DigitalLDOLogic_VIA1 $T=36910 29380 0 0 $X=36660 $Y=29150
X3169 1 DigitalLDOLogic_VIA1 $T=36910 33460 0 0 $X=36660 $Y=33230
X3170 1 DigitalLDOLogic_VIA1 $T=36910 37540 0 0 $X=36660 $Y=37310
X3171 1 DigitalLDOLogic_VIA1 $T=36910 41620 0 0 $X=36660 $Y=41390
X3172 1 DigitalLDOLogic_VIA1 $T=36910 45700 0 0 $X=36660 $Y=45470
X3173 1 DigitalLDOLogic_VIA1 $T=36910 49780 0 0 $X=36660 $Y=49550
X3174 1 DigitalLDOLogic_VIA1 $T=36910 53860 0 0 $X=36660 $Y=53630
X3175 1 DigitalLDOLogic_VIA1 $T=36910 57940 0 0 $X=36660 $Y=57710
X3176 3 DigitalLDOLogic_VIA1 $T=38750 11700 0 0 $X=38500 $Y=11470
X3177 3 DigitalLDOLogic_VIA1 $T=38750 15780 0 0 $X=38500 $Y=15550
X3178 3 DigitalLDOLogic_VIA1 $T=38750 19860 0 0 $X=38500 $Y=19630
X3179 3 DigitalLDOLogic_VIA1 $T=38750 23940 0 0 $X=38500 $Y=23710
X3180 3 DigitalLDOLogic_VIA1 $T=38750 28020 0 0 $X=38500 $Y=27790
X3181 3 DigitalLDOLogic_VIA1 $T=38750 32100 0 0 $X=38500 $Y=31870
X3182 3 DigitalLDOLogic_VIA1 $T=38750 36180 0 0 $X=38500 $Y=35950
X3183 3 DigitalLDOLogic_VIA1 $T=38750 40260 0 0 $X=38500 $Y=40030
X3184 3 DigitalLDOLogic_VIA1 $T=38750 44340 0 0 $X=38500 $Y=44110
X3185 3 DigitalLDOLogic_VIA1 $T=38750 48420 0 0 $X=38500 $Y=48190
X3186 3 DigitalLDOLogic_VIA1 $T=38750 52500 0 0 $X=38500 $Y=52270
X3187 3 DigitalLDOLogic_VIA1 $T=38750 56580 0 0 $X=38500 $Y=56350
X3188 1 DigitalLDOLogic_VIA1 $T=39670 13060 0 0 $X=39420 $Y=12830
X3189 1 DigitalLDOLogic_VIA1 $T=39670 17140 0 0 $X=39420 $Y=16910
X3190 1 DigitalLDOLogic_VIA1 $T=39670 21220 0 0 $X=39420 $Y=20990
X3191 1 DigitalLDOLogic_VIA1 $T=39670 25300 0 0 $X=39420 $Y=25070
X3192 1 DigitalLDOLogic_VIA1 $T=39670 29380 0 0 $X=39420 $Y=29150
X3193 1 DigitalLDOLogic_VIA1 $T=39670 33460 0 0 $X=39420 $Y=33230
X3194 1 DigitalLDOLogic_VIA1 $T=39670 37540 0 0 $X=39420 $Y=37310
X3195 1 DigitalLDOLogic_VIA1 $T=39670 41620 0 0 $X=39420 $Y=41390
X3196 1 DigitalLDOLogic_VIA1 $T=39670 45700 0 0 $X=39420 $Y=45470
X3197 1 DigitalLDOLogic_VIA1 $T=39670 49780 0 0 $X=39420 $Y=49550
X3198 1 DigitalLDOLogic_VIA1 $T=39670 53860 0 0 $X=39420 $Y=53630
X3199 1 DigitalLDOLogic_VIA1 $T=39670 57940 0 0 $X=39420 $Y=57710
X3200 3 DigitalLDOLogic_VIA1 $T=41510 11700 0 0 $X=41260 $Y=11470
X3201 3 DigitalLDOLogic_VIA1 $T=41510 15780 0 0 $X=41260 $Y=15550
X3202 3 DigitalLDOLogic_VIA1 $T=41510 19860 0 0 $X=41260 $Y=19630
X3203 3 DigitalLDOLogic_VIA1 $T=41510 23940 0 0 $X=41260 $Y=23710
X3204 3 DigitalLDOLogic_VIA1 $T=41510 28020 0 0 $X=41260 $Y=27790
X3205 3 DigitalLDOLogic_VIA1 $T=41510 32100 0 0 $X=41260 $Y=31870
X3206 3 DigitalLDOLogic_VIA1 $T=41510 36180 0 0 $X=41260 $Y=35950
X3207 3 DigitalLDOLogic_VIA1 $T=41510 40260 0 0 $X=41260 $Y=40030
X3208 3 DigitalLDOLogic_VIA1 $T=41510 44340 0 0 $X=41260 $Y=44110
X3209 3 DigitalLDOLogic_VIA1 $T=41510 48420 0 0 $X=41260 $Y=48190
X3210 3 DigitalLDOLogic_VIA1 $T=41510 52500 0 0 $X=41260 $Y=52270
X3211 3 DigitalLDOLogic_VIA1 $T=41510 56580 0 0 $X=41260 $Y=56350
X3212 1 DigitalLDOLogic_VIA1 $T=42430 13060 0 0 $X=42180 $Y=12830
X3213 1 DigitalLDOLogic_VIA1 $T=42430 17140 0 0 $X=42180 $Y=16910
X3214 1 DigitalLDOLogic_VIA1 $T=42430 21220 0 0 $X=42180 $Y=20990
X3215 1 DigitalLDOLogic_VIA1 $T=42430 25300 0 0 $X=42180 $Y=25070
X3216 1 DigitalLDOLogic_VIA1 $T=42430 29380 0 0 $X=42180 $Y=29150
X3217 1 DigitalLDOLogic_VIA1 $T=42430 33460 0 0 $X=42180 $Y=33230
X3218 1 DigitalLDOLogic_VIA1 $T=42430 37540 0 0 $X=42180 $Y=37310
X3219 1 DigitalLDOLogic_VIA1 $T=42430 41620 0 0 $X=42180 $Y=41390
X3220 1 DigitalLDOLogic_VIA1 $T=42430 45700 0 0 $X=42180 $Y=45470
X3221 1 DigitalLDOLogic_VIA1 $T=42430 49780 0 0 $X=42180 $Y=49550
X3222 1 DigitalLDOLogic_VIA1 $T=42430 53860 0 0 $X=42180 $Y=53630
X3223 1 DigitalLDOLogic_VIA1 $T=42430 57940 0 0 $X=42180 $Y=57710
X3224 3 DigitalLDOLogic_VIA1 $T=44270 11700 0 0 $X=44020 $Y=11470
X3225 3 DigitalLDOLogic_VIA1 $T=44270 15780 0 0 $X=44020 $Y=15550
X3226 3 DigitalLDOLogic_VIA1 $T=44270 19860 0 0 $X=44020 $Y=19630
X3227 3 DigitalLDOLogic_VIA1 $T=44270 23940 0 0 $X=44020 $Y=23710
X3228 3 DigitalLDOLogic_VIA1 $T=44270 28020 0 0 $X=44020 $Y=27790
X3229 3 DigitalLDOLogic_VIA1 $T=44270 32100 0 0 $X=44020 $Y=31870
X3230 3 DigitalLDOLogic_VIA1 $T=44270 36180 0 0 $X=44020 $Y=35950
X3231 3 DigitalLDOLogic_VIA1 $T=44270 40260 0 0 $X=44020 $Y=40030
X3232 3 DigitalLDOLogic_VIA1 $T=44270 44340 0 0 $X=44020 $Y=44110
X3233 3 DigitalLDOLogic_VIA1 $T=44270 48420 0 0 $X=44020 $Y=48190
X3234 3 DigitalLDOLogic_VIA1 $T=44270 52500 0 0 $X=44020 $Y=52270
X3235 3 DigitalLDOLogic_VIA1 $T=44270 56580 0 0 $X=44020 $Y=56350
X3236 1 DigitalLDOLogic_VIA1 $T=45190 13060 0 0 $X=44940 $Y=12830
X3237 1 DigitalLDOLogic_VIA1 $T=45190 17140 0 0 $X=44940 $Y=16910
X3238 1 DigitalLDOLogic_VIA1 $T=45190 21220 0 0 $X=44940 $Y=20990
X3239 1 DigitalLDOLogic_VIA1 $T=45190 25300 0 0 $X=44940 $Y=25070
X3240 1 DigitalLDOLogic_VIA1 $T=45190 29380 0 0 $X=44940 $Y=29150
X3241 1 DigitalLDOLogic_VIA1 $T=45190 33460 0 0 $X=44940 $Y=33230
X3242 1 DigitalLDOLogic_VIA1 $T=45190 37540 0 0 $X=44940 $Y=37310
X3243 1 DigitalLDOLogic_VIA1 $T=45190 41620 0 0 $X=44940 $Y=41390
X3244 1 DigitalLDOLogic_VIA1 $T=45190 45700 0 0 $X=44940 $Y=45470
X3245 1 DigitalLDOLogic_VIA1 $T=45190 49780 0 0 $X=44940 $Y=49550
X3246 1 DigitalLDOLogic_VIA1 $T=45190 53860 0 0 $X=44940 $Y=53630
X3247 1 DigitalLDOLogic_VIA1 $T=45190 57940 0 0 $X=44940 $Y=57710
X3248 3 DigitalLDOLogic_VIA1 $T=47030 11700 0 0 $X=46780 $Y=11470
X3249 3 DigitalLDOLogic_VIA1 $T=47030 15780 0 0 $X=46780 $Y=15550
X3250 3 DigitalLDOLogic_VIA1 $T=47030 19860 0 0 $X=46780 $Y=19630
X3251 3 DigitalLDOLogic_VIA1 $T=47030 23940 0 0 $X=46780 $Y=23710
X3252 3 DigitalLDOLogic_VIA1 $T=47030 28020 0 0 $X=46780 $Y=27790
X3253 3 DigitalLDOLogic_VIA1 $T=47030 32100 0 0 $X=46780 $Y=31870
X3254 3 DigitalLDOLogic_VIA1 $T=47030 36180 0 0 $X=46780 $Y=35950
X3255 3 DigitalLDOLogic_VIA1 $T=47030 40260 0 0 $X=46780 $Y=40030
X3256 3 DigitalLDOLogic_VIA1 $T=47030 44340 0 0 $X=46780 $Y=44110
X3257 3 DigitalLDOLogic_VIA1 $T=47030 48420 0 0 $X=46780 $Y=48190
X3258 3 DigitalLDOLogic_VIA1 $T=47030 52500 0 0 $X=46780 $Y=52270
X3259 3 DigitalLDOLogic_VIA1 $T=47030 56580 0 0 $X=46780 $Y=56350
X3260 1 DigitalLDOLogic_VIA1 $T=47950 13060 0 0 $X=47700 $Y=12830
X3261 1 DigitalLDOLogic_VIA1 $T=47950 17140 0 0 $X=47700 $Y=16910
X3262 1 DigitalLDOLogic_VIA1 $T=47950 21220 0 0 $X=47700 $Y=20990
X3263 1 DigitalLDOLogic_VIA1 $T=47950 25300 0 0 $X=47700 $Y=25070
X3264 1 DigitalLDOLogic_VIA1 $T=47950 29380 0 0 $X=47700 $Y=29150
X3265 1 DigitalLDOLogic_VIA1 $T=47950 33460 0 0 $X=47700 $Y=33230
X3266 1 DigitalLDOLogic_VIA1 $T=47950 37540 0 0 $X=47700 $Y=37310
X3267 1 DigitalLDOLogic_VIA1 $T=47950 41620 0 0 $X=47700 $Y=41390
X3268 1 DigitalLDOLogic_VIA1 $T=47950 45700 0 0 $X=47700 $Y=45470
X3269 1 DigitalLDOLogic_VIA1 $T=47950 49780 0 0 $X=47700 $Y=49550
X3270 1 DigitalLDOLogic_VIA1 $T=47950 53860 0 0 $X=47700 $Y=53630
X3271 1 DigitalLDOLogic_VIA1 $T=47950 57940 0 0 $X=47700 $Y=57710
X3272 3 DigitalLDOLogic_VIA1 $T=49790 11700 0 0 $X=49540 $Y=11470
X3273 3 DigitalLDOLogic_VIA1 $T=49790 15780 0 0 $X=49540 $Y=15550
X3274 3 DigitalLDOLogic_VIA1 $T=49790 19860 0 0 $X=49540 $Y=19630
X3275 3 DigitalLDOLogic_VIA1 $T=49790 23940 0 0 $X=49540 $Y=23710
X3276 3 DigitalLDOLogic_VIA1 $T=49790 28020 0 0 $X=49540 $Y=27790
X3277 3 DigitalLDOLogic_VIA1 $T=49790 32100 0 0 $X=49540 $Y=31870
X3278 3 DigitalLDOLogic_VIA1 $T=49790 36180 0 0 $X=49540 $Y=35950
X3279 3 DigitalLDOLogic_VIA1 $T=49790 40260 0 0 $X=49540 $Y=40030
X3280 3 DigitalLDOLogic_VIA1 $T=49790 44340 0 0 $X=49540 $Y=44110
X3281 3 DigitalLDOLogic_VIA1 $T=49790 48420 0 0 $X=49540 $Y=48190
X3282 3 DigitalLDOLogic_VIA1 $T=49790 52500 0 0 $X=49540 $Y=52270
X3283 3 DigitalLDOLogic_VIA1 $T=49790 56580 0 0 $X=49540 $Y=56350
X3284 1 DigitalLDOLogic_VIA1 $T=50710 13060 0 0 $X=50460 $Y=12830
X3285 1 DigitalLDOLogic_VIA1 $T=50710 17140 0 0 $X=50460 $Y=16910
X3286 1 DigitalLDOLogic_VIA1 $T=50710 21220 0 0 $X=50460 $Y=20990
X3287 1 DigitalLDOLogic_VIA1 $T=50710 25300 0 0 $X=50460 $Y=25070
X3288 1 DigitalLDOLogic_VIA1 $T=50710 29380 0 0 $X=50460 $Y=29150
X3289 1 DigitalLDOLogic_VIA1 $T=50710 33460 0 0 $X=50460 $Y=33230
X3290 1 DigitalLDOLogic_VIA1 $T=50710 37540 0 0 $X=50460 $Y=37310
X3291 1 DigitalLDOLogic_VIA1 $T=50710 41620 0 0 $X=50460 $Y=41390
X3292 1 DigitalLDOLogic_VIA1 $T=50710 45700 0 0 $X=50460 $Y=45470
X3293 1 DigitalLDOLogic_VIA1 $T=50710 49780 0 0 $X=50460 $Y=49550
X3294 1 DigitalLDOLogic_VIA1 $T=50710 53860 0 0 $X=50460 $Y=53630
X3295 1 DigitalLDOLogic_VIA1 $T=50710 57940 0 0 $X=50460 $Y=57710
X3296 3 DigitalLDOLogic_VIA1 $T=52550 11700 0 0 $X=52300 $Y=11470
X3297 3 DigitalLDOLogic_VIA1 $T=52550 15780 0 0 $X=52300 $Y=15550
X3298 3 DigitalLDOLogic_VIA1 $T=52550 19860 0 0 $X=52300 $Y=19630
X3299 3 DigitalLDOLogic_VIA1 $T=52550 23940 0 0 $X=52300 $Y=23710
X3300 3 DigitalLDOLogic_VIA1 $T=52550 28020 0 0 $X=52300 $Y=27790
X3301 3 DigitalLDOLogic_VIA1 $T=52550 32100 0 0 $X=52300 $Y=31870
X3302 3 DigitalLDOLogic_VIA1 $T=52550 36180 0 0 $X=52300 $Y=35950
X3303 3 DigitalLDOLogic_VIA1 $T=52550 40260 0 0 $X=52300 $Y=40030
X3304 3 DigitalLDOLogic_VIA1 $T=52550 44340 0 0 $X=52300 $Y=44110
X3305 3 DigitalLDOLogic_VIA1 $T=52550 48420 0 0 $X=52300 $Y=48190
X3306 3 DigitalLDOLogic_VIA1 $T=52550 52500 0 0 $X=52300 $Y=52270
X3307 3 DigitalLDOLogic_VIA1 $T=52550 56580 0 0 $X=52300 $Y=56350
X3308 1 DigitalLDOLogic_VIA1 $T=53470 13060 0 0 $X=53220 $Y=12830
X3309 1 DigitalLDOLogic_VIA1 $T=53470 17140 0 0 $X=53220 $Y=16910
X3310 1 DigitalLDOLogic_VIA1 $T=53470 21220 0 0 $X=53220 $Y=20990
X3311 1 DigitalLDOLogic_VIA1 $T=53470 25300 0 0 $X=53220 $Y=25070
X3312 1 DigitalLDOLogic_VIA1 $T=53470 29380 0 0 $X=53220 $Y=29150
X3313 1 DigitalLDOLogic_VIA1 $T=53470 33460 0 0 $X=53220 $Y=33230
X3314 1 DigitalLDOLogic_VIA1 $T=53470 37540 0 0 $X=53220 $Y=37310
X3315 1 DigitalLDOLogic_VIA1 $T=53470 41620 0 0 $X=53220 $Y=41390
X3316 1 DigitalLDOLogic_VIA1 $T=53470 45700 0 0 $X=53220 $Y=45470
X3317 1 DigitalLDOLogic_VIA1 $T=53470 49780 0 0 $X=53220 $Y=49550
X3318 1 DigitalLDOLogic_VIA1 $T=53470 53860 0 0 $X=53220 $Y=53630
X3319 1 DigitalLDOLogic_VIA1 $T=53470 57940 0 0 $X=53220 $Y=57710
X3320 3 DigitalLDOLogic_VIA1 $T=55310 11700 0 0 $X=55060 $Y=11470
X3321 3 DigitalLDOLogic_VIA1 $T=55310 15780 0 0 $X=55060 $Y=15550
X3322 3 DigitalLDOLogic_VIA1 $T=55310 19860 0 0 $X=55060 $Y=19630
X3323 3 DigitalLDOLogic_VIA1 $T=55310 23940 0 0 $X=55060 $Y=23710
X3324 3 DigitalLDOLogic_VIA1 $T=55310 28020 0 0 $X=55060 $Y=27790
X3325 3 DigitalLDOLogic_VIA1 $T=55310 32100 0 0 $X=55060 $Y=31870
X3326 3 DigitalLDOLogic_VIA1 $T=55310 36180 0 0 $X=55060 $Y=35950
X3327 3 DigitalLDOLogic_VIA1 $T=55310 40260 0 0 $X=55060 $Y=40030
X3328 3 DigitalLDOLogic_VIA1 $T=55310 44340 0 0 $X=55060 $Y=44110
X3329 3 DigitalLDOLogic_VIA1 $T=55310 48420 0 0 $X=55060 $Y=48190
X3330 3 DigitalLDOLogic_VIA1 $T=55310 52500 0 0 $X=55060 $Y=52270
X3331 3 DigitalLDOLogic_VIA1 $T=55310 56580 0 0 $X=55060 $Y=56350
X3332 1 DigitalLDOLogic_VIA1 $T=56230 13060 0 0 $X=55980 $Y=12830
X3333 1 DigitalLDOLogic_VIA1 $T=56230 17140 0 0 $X=55980 $Y=16910
X3334 1 DigitalLDOLogic_VIA1 $T=56230 21220 0 0 $X=55980 $Y=20990
X3335 1 DigitalLDOLogic_VIA1 $T=56230 25300 0 0 $X=55980 $Y=25070
X3336 1 DigitalLDOLogic_VIA1 $T=56230 29380 0 0 $X=55980 $Y=29150
X3337 1 DigitalLDOLogic_VIA1 $T=56230 33460 0 0 $X=55980 $Y=33230
X3338 1 DigitalLDOLogic_VIA1 $T=56230 37540 0 0 $X=55980 $Y=37310
X3339 1 DigitalLDOLogic_VIA1 $T=56230 41620 0 0 $X=55980 $Y=41390
X3340 1 DigitalLDOLogic_VIA1 $T=56230 45700 0 0 $X=55980 $Y=45470
X3341 1 DigitalLDOLogic_VIA1 $T=56230 49780 0 0 $X=55980 $Y=49550
X3342 1 DigitalLDOLogic_VIA1 $T=56230 53860 0 0 $X=55980 $Y=53630
X3343 1 DigitalLDOLogic_VIA1 $T=56230 57940 0 0 $X=55980 $Y=57710
X3344 3 DigitalLDOLogic_VIA1 $T=58070 11700 0 0 $X=57820 $Y=11470
X3345 3 DigitalLDOLogic_VIA1 $T=58070 15780 0 0 $X=57820 $Y=15550
X3346 3 DigitalLDOLogic_VIA1 $T=58070 19860 0 0 $X=57820 $Y=19630
X3347 3 DigitalLDOLogic_VIA1 $T=58070 23940 0 0 $X=57820 $Y=23710
X3348 3 DigitalLDOLogic_VIA1 $T=58070 28020 0 0 $X=57820 $Y=27790
X3349 3 DigitalLDOLogic_VIA1 $T=58070 32100 0 0 $X=57820 $Y=31870
X3350 3 DigitalLDOLogic_VIA1 $T=58070 36180 0 0 $X=57820 $Y=35950
X3351 3 DigitalLDOLogic_VIA1 $T=58070 40260 0 0 $X=57820 $Y=40030
X3352 3 DigitalLDOLogic_VIA1 $T=58070 44340 0 0 $X=57820 $Y=44110
X3353 3 DigitalLDOLogic_VIA1 $T=58070 48420 0 0 $X=57820 $Y=48190
X3354 3 DigitalLDOLogic_VIA1 $T=58070 52500 0 0 $X=57820 $Y=52270
X3355 3 DigitalLDOLogic_VIA1 $T=58070 56580 0 0 $X=57820 $Y=56350
X3356 1 DigitalLDOLogic_VIA1 $T=58990 13060 0 0 $X=58740 $Y=12830
X3357 1 DigitalLDOLogic_VIA1 $T=58990 17140 0 0 $X=58740 $Y=16910
X3358 1 DigitalLDOLogic_VIA1 $T=58990 21220 0 0 $X=58740 $Y=20990
X3359 1 DigitalLDOLogic_VIA1 $T=58990 25300 0 0 $X=58740 $Y=25070
X3360 1 DigitalLDOLogic_VIA1 $T=58990 29380 0 0 $X=58740 $Y=29150
X3361 1 DigitalLDOLogic_VIA1 $T=58990 33460 0 0 $X=58740 $Y=33230
X3362 1 DigitalLDOLogic_VIA1 $T=58990 37540 0 0 $X=58740 $Y=37310
X3363 1 DigitalLDOLogic_VIA1 $T=58990 41620 0 0 $X=58740 $Y=41390
X3364 1 DigitalLDOLogic_VIA1 $T=58990 45700 0 0 $X=58740 $Y=45470
X3365 1 DigitalLDOLogic_VIA1 $T=58990 49780 0 0 $X=58740 $Y=49550
X3366 1 DigitalLDOLogic_VIA1 $T=58990 53860 0 0 $X=58740 $Y=53630
X3367 1 DigitalLDOLogic_VIA1 $T=58990 57940 0 0 $X=58740 $Y=57710
X3368 3 DigitalLDOLogic_VIA1 $T=60830 11700 0 0 $X=60580 $Y=11470
X3369 3 DigitalLDOLogic_VIA1 $T=60830 15780 0 0 $X=60580 $Y=15550
X3370 3 DigitalLDOLogic_VIA1 $T=60830 19860 0 0 $X=60580 $Y=19630
X3371 3 DigitalLDOLogic_VIA1 $T=60830 23940 0 0 $X=60580 $Y=23710
X3372 3 DigitalLDOLogic_VIA1 $T=60830 28020 0 0 $X=60580 $Y=27790
X3373 3 DigitalLDOLogic_VIA1 $T=60830 32100 0 0 $X=60580 $Y=31870
X3374 3 DigitalLDOLogic_VIA1 $T=60830 36180 0 0 $X=60580 $Y=35950
X3375 3 DigitalLDOLogic_VIA1 $T=60830 40260 0 0 $X=60580 $Y=40030
X3376 3 DigitalLDOLogic_VIA1 $T=60830 44340 0 0 $X=60580 $Y=44110
X3377 3 DigitalLDOLogic_VIA1 $T=60830 48420 0 0 $X=60580 $Y=48190
X3378 3 DigitalLDOLogic_VIA1 $T=60830 52500 0 0 $X=60580 $Y=52270
X3379 3 DigitalLDOLogic_VIA1 $T=60830 56580 0 0 $X=60580 $Y=56350
X3380 1 DigitalLDOLogic_VIA1 $T=61750 13060 0 0 $X=61500 $Y=12830
X3381 1 DigitalLDOLogic_VIA1 $T=61750 17140 0 0 $X=61500 $Y=16910
X3382 1 DigitalLDOLogic_VIA1 $T=61750 21220 0 0 $X=61500 $Y=20990
X3383 1 DigitalLDOLogic_VIA1 $T=61750 25300 0 0 $X=61500 $Y=25070
X3384 1 DigitalLDOLogic_VIA1 $T=61750 29380 0 0 $X=61500 $Y=29150
X3385 1 DigitalLDOLogic_VIA1 $T=61750 33460 0 0 $X=61500 $Y=33230
X3386 1 DigitalLDOLogic_VIA1 $T=61750 37540 0 0 $X=61500 $Y=37310
X3387 1 DigitalLDOLogic_VIA1 $T=61750 41620 0 0 $X=61500 $Y=41390
X3388 1 DigitalLDOLogic_VIA1 $T=61750 45700 0 0 $X=61500 $Y=45470
X3389 1 DigitalLDOLogic_VIA1 $T=61750 49780 0 0 $X=61500 $Y=49550
X3390 1 DigitalLDOLogic_VIA1 $T=61750 53860 0 0 $X=61500 $Y=53630
X3391 1 DigitalLDOLogic_VIA1 $T=61750 57940 0 0 $X=61500 $Y=57710
X3392 3 DigitalLDOLogic_VIA1 $T=63590 11700 0 0 $X=63340 $Y=11470
X3393 3 DigitalLDOLogic_VIA1 $T=63590 15780 0 0 $X=63340 $Y=15550
X3394 3 DigitalLDOLogic_VIA1 $T=63590 19860 0 0 $X=63340 $Y=19630
X3395 3 DigitalLDOLogic_VIA1 $T=63590 23940 0 0 $X=63340 $Y=23710
X3396 3 DigitalLDOLogic_VIA1 $T=63590 28020 0 0 $X=63340 $Y=27790
X3397 3 DigitalLDOLogic_VIA1 $T=63590 32100 0 0 $X=63340 $Y=31870
X3398 3 DigitalLDOLogic_VIA1 $T=63590 36180 0 0 $X=63340 $Y=35950
X3399 3 DigitalLDOLogic_VIA1 $T=63590 40260 0 0 $X=63340 $Y=40030
X3400 3 DigitalLDOLogic_VIA1 $T=63590 44340 0 0 $X=63340 $Y=44110
X3401 3 DigitalLDOLogic_VIA1 $T=63590 48420 0 0 $X=63340 $Y=48190
X3402 3 DigitalLDOLogic_VIA1 $T=63590 52500 0 0 $X=63340 $Y=52270
X3403 3 DigitalLDOLogic_VIA1 $T=63590 56580 0 0 $X=63340 $Y=56350
X3404 1 DigitalLDOLogic_VIA1 $T=64510 13060 0 0 $X=64260 $Y=12830
X3405 1 DigitalLDOLogic_VIA1 $T=64510 17140 0 0 $X=64260 $Y=16910
X3406 1 DigitalLDOLogic_VIA1 $T=64510 21220 0 0 $X=64260 $Y=20990
X3407 1 DigitalLDOLogic_VIA1 $T=64510 25300 0 0 $X=64260 $Y=25070
X3408 1 DigitalLDOLogic_VIA1 $T=64510 29380 0 0 $X=64260 $Y=29150
X3409 1 DigitalLDOLogic_VIA1 $T=64510 33460 0 0 $X=64260 $Y=33230
X3410 1 DigitalLDOLogic_VIA1 $T=64510 37540 0 0 $X=64260 $Y=37310
X3411 1 DigitalLDOLogic_VIA1 $T=64510 41620 0 0 $X=64260 $Y=41390
X3412 1 DigitalLDOLogic_VIA1 $T=64510 45700 0 0 $X=64260 $Y=45470
X3413 1 DigitalLDOLogic_VIA1 $T=64510 49780 0 0 $X=64260 $Y=49550
X3414 1 DigitalLDOLogic_VIA1 $T=64510 53860 0 0 $X=64260 $Y=53630
X3415 1 DigitalLDOLogic_VIA1 $T=64510 57940 0 0 $X=64260 $Y=57710
X3416 3 DigitalLDOLogic_VIA1 $T=66350 11700 0 0 $X=66100 $Y=11470
X3417 3 DigitalLDOLogic_VIA1 $T=66350 15780 0 0 $X=66100 $Y=15550
X3418 3 DigitalLDOLogic_VIA1 $T=66350 19860 0 0 $X=66100 $Y=19630
X3419 3 DigitalLDOLogic_VIA1 $T=66350 23940 0 0 $X=66100 $Y=23710
X3420 3 DigitalLDOLogic_VIA1 $T=66350 28020 0 0 $X=66100 $Y=27790
X3421 3 DigitalLDOLogic_VIA1 $T=66350 32100 0 0 $X=66100 $Y=31870
X3422 3 DigitalLDOLogic_VIA1 $T=66350 36180 0 0 $X=66100 $Y=35950
X3423 3 DigitalLDOLogic_VIA1 $T=66350 40260 0 0 $X=66100 $Y=40030
X3424 3 DigitalLDOLogic_VIA1 $T=66350 44340 0 0 $X=66100 $Y=44110
X3425 3 DigitalLDOLogic_VIA1 $T=66350 48420 0 0 $X=66100 $Y=48190
X3426 3 DigitalLDOLogic_VIA1 $T=66350 52500 0 0 $X=66100 $Y=52270
X3427 3 DigitalLDOLogic_VIA1 $T=66350 56580 0 0 $X=66100 $Y=56350
X3428 1 DigitalLDOLogic_VIA1 $T=67270 13060 0 0 $X=67020 $Y=12830
X3429 1 DigitalLDOLogic_VIA1 $T=67270 17140 0 0 $X=67020 $Y=16910
X3430 1 DigitalLDOLogic_VIA1 $T=67270 21220 0 0 $X=67020 $Y=20990
X3431 1 DigitalLDOLogic_VIA1 $T=67270 25300 0 0 $X=67020 $Y=25070
X3432 1 DigitalLDOLogic_VIA1 $T=67270 29380 0 0 $X=67020 $Y=29150
X3433 1 DigitalLDOLogic_VIA1 $T=67270 33460 0 0 $X=67020 $Y=33230
X3434 1 DigitalLDOLogic_VIA1 $T=67270 37540 0 0 $X=67020 $Y=37310
X3435 1 DigitalLDOLogic_VIA1 $T=67270 41620 0 0 $X=67020 $Y=41390
X3436 1 DigitalLDOLogic_VIA1 $T=67270 45700 0 0 $X=67020 $Y=45470
X3437 1 DigitalLDOLogic_VIA1 $T=67270 49780 0 0 $X=67020 $Y=49550
X3438 1 DigitalLDOLogic_VIA1 $T=67270 53860 0 0 $X=67020 $Y=53630
X3439 1 DigitalLDOLogic_VIA1 $T=67270 57940 0 0 $X=67020 $Y=57710
X3440 3 DigitalLDOLogic_VIA1 $T=69110 11700 0 0 $X=68860 $Y=11470
X3441 3 DigitalLDOLogic_VIA1 $T=69110 15780 0 0 $X=68860 $Y=15550
X3442 3 DigitalLDOLogic_VIA1 $T=69110 19860 0 0 $X=68860 $Y=19630
X3443 3 DigitalLDOLogic_VIA1 $T=69110 23940 0 0 $X=68860 $Y=23710
X3444 3 DigitalLDOLogic_VIA1 $T=69110 28020 0 0 $X=68860 $Y=27790
X3445 3 DigitalLDOLogic_VIA1 $T=69110 32100 0 0 $X=68860 $Y=31870
X3446 3 DigitalLDOLogic_VIA1 $T=69110 36180 0 0 $X=68860 $Y=35950
X3447 3 DigitalLDOLogic_VIA1 $T=69110 40260 0 0 $X=68860 $Y=40030
X3448 3 DigitalLDOLogic_VIA1 $T=69110 44340 0 0 $X=68860 $Y=44110
X3449 3 DigitalLDOLogic_VIA1 $T=69110 48420 0 0 $X=68860 $Y=48190
X3450 3 DigitalLDOLogic_VIA1 $T=69110 52500 0 0 $X=68860 $Y=52270
X3451 3 DigitalLDOLogic_VIA1 $T=69110 56580 0 0 $X=68860 $Y=56350
X3452 1 DigitalLDOLogic_VIA1 $T=70030 13060 0 0 $X=69780 $Y=12830
X3453 1 DigitalLDOLogic_VIA1 $T=70030 17140 0 0 $X=69780 $Y=16910
X3454 1 DigitalLDOLogic_VIA1 $T=70030 21220 0 0 $X=69780 $Y=20990
X3455 1 DigitalLDOLogic_VIA1 $T=70030 25300 0 0 $X=69780 $Y=25070
X3456 1 DigitalLDOLogic_VIA1 $T=70030 29380 0 0 $X=69780 $Y=29150
X3457 1 DigitalLDOLogic_VIA1 $T=70030 33460 0 0 $X=69780 $Y=33230
X3458 1 DigitalLDOLogic_VIA1 $T=70030 37540 0 0 $X=69780 $Y=37310
X3459 1 DigitalLDOLogic_VIA1 $T=70030 41620 0 0 $X=69780 $Y=41390
X3460 1 DigitalLDOLogic_VIA1 $T=70030 45700 0 0 $X=69780 $Y=45470
X3461 1 DigitalLDOLogic_VIA1 $T=70030 49780 0 0 $X=69780 $Y=49550
X3462 1 DigitalLDOLogic_VIA1 $T=70030 53860 0 0 $X=69780 $Y=53630
X3463 1 DigitalLDOLogic_VIA1 $T=70030 57940 0 0 $X=69780 $Y=57710
X3464 3 DigitalLDOLogic_VIA1 $T=71870 11700 0 0 $X=71620 $Y=11470
X3465 3 DigitalLDOLogic_VIA1 $T=71870 15780 0 0 $X=71620 $Y=15550
X3466 3 DigitalLDOLogic_VIA1 $T=71870 19860 0 0 $X=71620 $Y=19630
X3467 3 DigitalLDOLogic_VIA1 $T=71870 23940 0 0 $X=71620 $Y=23710
X3468 3 DigitalLDOLogic_VIA1 $T=71870 28020 0 0 $X=71620 $Y=27790
X3469 3 DigitalLDOLogic_VIA1 $T=71870 32100 0 0 $X=71620 $Y=31870
X3470 3 DigitalLDOLogic_VIA1 $T=71870 36180 0 0 $X=71620 $Y=35950
X3471 3 DigitalLDOLogic_VIA1 $T=71870 40260 0 0 $X=71620 $Y=40030
X3472 3 DigitalLDOLogic_VIA1 $T=71870 44340 0 0 $X=71620 $Y=44110
X3473 3 DigitalLDOLogic_VIA1 $T=71870 48420 0 0 $X=71620 $Y=48190
X3474 3 DigitalLDOLogic_VIA1 $T=71870 52500 0 0 $X=71620 $Y=52270
X3475 3 DigitalLDOLogic_VIA1 $T=71870 56580 0 0 $X=71620 $Y=56350
X3476 1 DigitalLDOLogic_VIA1 $T=72790 13060 0 0 $X=72540 $Y=12830
X3477 1 DigitalLDOLogic_VIA1 $T=72790 17140 0 0 $X=72540 $Y=16910
X3478 1 DigitalLDOLogic_VIA1 $T=72790 21220 0 0 $X=72540 $Y=20990
X3479 1 DigitalLDOLogic_VIA1 $T=72790 25300 0 0 $X=72540 $Y=25070
X3480 1 DigitalLDOLogic_VIA1 $T=72790 29380 0 0 $X=72540 $Y=29150
X3481 1 DigitalLDOLogic_VIA1 $T=72790 33460 0 0 $X=72540 $Y=33230
X3482 1 DigitalLDOLogic_VIA1 $T=72790 37540 0 0 $X=72540 $Y=37310
X3483 1 DigitalLDOLogic_VIA1 $T=72790 41620 0 0 $X=72540 $Y=41390
X3484 1 DigitalLDOLogic_VIA1 $T=72790 45700 0 0 $X=72540 $Y=45470
X3485 1 DigitalLDOLogic_VIA1 $T=72790 49780 0 0 $X=72540 $Y=49550
X3486 1 DigitalLDOLogic_VIA1 $T=72790 53860 0 0 $X=72540 $Y=53630
X3487 1 DigitalLDOLogic_VIA1 $T=72790 57940 0 0 $X=72540 $Y=57710
X3488 3 DigitalLDOLogic_VIA1 $T=74630 11700 0 0 $X=74380 $Y=11470
X3489 3 DigitalLDOLogic_VIA1 $T=74630 15780 0 0 $X=74380 $Y=15550
X3490 3 DigitalLDOLogic_VIA1 $T=74630 19860 0 0 $X=74380 $Y=19630
X3491 3 DigitalLDOLogic_VIA1 $T=74630 23940 0 0 $X=74380 $Y=23710
X3492 3 DigitalLDOLogic_VIA1 $T=74630 28020 0 0 $X=74380 $Y=27790
X3493 3 DigitalLDOLogic_VIA1 $T=74630 32100 0 0 $X=74380 $Y=31870
X3494 3 DigitalLDOLogic_VIA1 $T=74630 36180 0 0 $X=74380 $Y=35950
X3495 3 DigitalLDOLogic_VIA1 $T=74630 40260 0 0 $X=74380 $Y=40030
X3496 3 DigitalLDOLogic_VIA1 $T=74630 44340 0 0 $X=74380 $Y=44110
X3497 3 DigitalLDOLogic_VIA1 $T=74630 48420 0 0 $X=74380 $Y=48190
X3498 3 DigitalLDOLogic_VIA1 $T=74630 52500 0 0 $X=74380 $Y=52270
X3499 3 DigitalLDOLogic_VIA1 $T=74630 56580 0 0 $X=74380 $Y=56350
X3500 1 DigitalLDOLogic_VIA1 $T=75550 13060 0 0 $X=75300 $Y=12830
X3501 1 DigitalLDOLogic_VIA1 $T=75550 17140 0 0 $X=75300 $Y=16910
X3502 1 DigitalLDOLogic_VIA1 $T=75550 21220 0 0 $X=75300 $Y=20990
X3503 1 DigitalLDOLogic_VIA1 $T=75550 25300 0 0 $X=75300 $Y=25070
X3504 1 DigitalLDOLogic_VIA1 $T=75550 29380 0 0 $X=75300 $Y=29150
X3505 1 DigitalLDOLogic_VIA1 $T=75550 33460 0 0 $X=75300 $Y=33230
X3506 1 DigitalLDOLogic_VIA1 $T=75550 37540 0 0 $X=75300 $Y=37310
X3507 1 DigitalLDOLogic_VIA1 $T=75550 41620 0 0 $X=75300 $Y=41390
X3508 1 DigitalLDOLogic_VIA1 $T=75550 45700 0 0 $X=75300 $Y=45470
X3509 1 DigitalLDOLogic_VIA1 $T=75550 49780 0 0 $X=75300 $Y=49550
X3510 1 DigitalLDOLogic_VIA1 $T=75550 53860 0 0 $X=75300 $Y=53630
X3511 1 DigitalLDOLogic_VIA1 $T=75550 57940 0 0 $X=75300 $Y=57710
X3512 3 DigitalLDOLogic_VIA1 $T=77390 11700 0 0 $X=77140 $Y=11470
X3513 3 DigitalLDOLogic_VIA1 $T=77390 15780 0 0 $X=77140 $Y=15550
X3514 3 DigitalLDOLogic_VIA1 $T=77390 19860 0 0 $X=77140 $Y=19630
X3515 3 DigitalLDOLogic_VIA1 $T=77390 23940 0 0 $X=77140 $Y=23710
X3516 3 DigitalLDOLogic_VIA1 $T=77390 28020 0 0 $X=77140 $Y=27790
X3517 3 DigitalLDOLogic_VIA1 $T=77390 32100 0 0 $X=77140 $Y=31870
X3518 3 DigitalLDOLogic_VIA1 $T=77390 36180 0 0 $X=77140 $Y=35950
X3519 3 DigitalLDOLogic_VIA1 $T=77390 40260 0 0 $X=77140 $Y=40030
X3520 3 DigitalLDOLogic_VIA1 $T=77390 44340 0 0 $X=77140 $Y=44110
X3521 3 DigitalLDOLogic_VIA1 $T=77390 48420 0 0 $X=77140 $Y=48190
X3522 3 DigitalLDOLogic_VIA1 $T=77390 52500 0 0 $X=77140 $Y=52270
X3523 3 DigitalLDOLogic_VIA1 $T=77390 56580 0 0 $X=77140 $Y=56350
X3524 1 DigitalLDOLogic_VIA1 $T=78310 13060 0 0 $X=78060 $Y=12830
X3525 1 DigitalLDOLogic_VIA1 $T=78310 17140 0 0 $X=78060 $Y=16910
X3526 1 DigitalLDOLogic_VIA1 $T=78310 21220 0 0 $X=78060 $Y=20990
X3527 1 DigitalLDOLogic_VIA1 $T=78310 25300 0 0 $X=78060 $Y=25070
X3528 1 DigitalLDOLogic_VIA1 $T=78310 29380 0 0 $X=78060 $Y=29150
X3529 1 DigitalLDOLogic_VIA1 $T=78310 33460 0 0 $X=78060 $Y=33230
X3530 1 DigitalLDOLogic_VIA1 $T=78310 37540 0 0 $X=78060 $Y=37310
X3531 1 DigitalLDOLogic_VIA1 $T=78310 41620 0 0 $X=78060 $Y=41390
X3532 1 DigitalLDOLogic_VIA1 $T=78310 45700 0 0 $X=78060 $Y=45470
X3533 1 DigitalLDOLogic_VIA1 $T=78310 49780 0 0 $X=78060 $Y=49550
X3534 1 DigitalLDOLogic_VIA1 $T=78310 53860 0 0 $X=78060 $Y=53630
X3535 1 DigitalLDOLogic_VIA1 $T=78310 57940 0 0 $X=78060 $Y=57710
X3536 3 DigitalLDOLogic_VIA1 $T=80150 11700 0 0 $X=79900 $Y=11470
X3537 3 DigitalLDOLogic_VIA1 $T=80150 15780 0 0 $X=79900 $Y=15550
X3538 3 DigitalLDOLogic_VIA1 $T=80150 19860 0 0 $X=79900 $Y=19630
X3539 3 DigitalLDOLogic_VIA1 $T=80150 23940 0 0 $X=79900 $Y=23710
X3540 3 DigitalLDOLogic_VIA1 $T=80150 28020 0 0 $X=79900 $Y=27790
X3541 3 DigitalLDOLogic_VIA1 $T=80150 32100 0 0 $X=79900 $Y=31870
X3542 3 DigitalLDOLogic_VIA1 $T=80150 36180 0 0 $X=79900 $Y=35950
X3543 3 DigitalLDOLogic_VIA1 $T=80150 40260 0 0 $X=79900 $Y=40030
X3544 3 DigitalLDOLogic_VIA1 $T=80150 44340 0 0 $X=79900 $Y=44110
X3545 3 DigitalLDOLogic_VIA1 $T=80150 48420 0 0 $X=79900 $Y=48190
X3546 3 DigitalLDOLogic_VIA1 $T=80150 52500 0 0 $X=79900 $Y=52270
X3547 3 DigitalLDOLogic_VIA1 $T=80150 56580 0 0 $X=79900 $Y=56350
X3548 1 DigitalLDOLogic_VIA1 $T=81070 13060 0 0 $X=80820 $Y=12830
X3549 1 DigitalLDOLogic_VIA1 $T=81070 17140 0 0 $X=80820 $Y=16910
X3550 1 DigitalLDOLogic_VIA1 $T=81070 21220 0 0 $X=80820 $Y=20990
X3551 1 DigitalLDOLogic_VIA1 $T=81070 25300 0 0 $X=80820 $Y=25070
X3552 1 DigitalLDOLogic_VIA1 $T=81070 29380 0 0 $X=80820 $Y=29150
X3553 1 DigitalLDOLogic_VIA1 $T=81070 33460 0 0 $X=80820 $Y=33230
X3554 1 DigitalLDOLogic_VIA1 $T=81070 37540 0 0 $X=80820 $Y=37310
X3555 1 DigitalLDOLogic_VIA1 $T=81070 41620 0 0 $X=80820 $Y=41390
X3556 1 DigitalLDOLogic_VIA1 $T=81070 45700 0 0 $X=80820 $Y=45470
X3557 1 DigitalLDOLogic_VIA1 $T=81070 49780 0 0 $X=80820 $Y=49550
X3558 1 DigitalLDOLogic_VIA1 $T=81070 53860 0 0 $X=80820 $Y=53630
X3559 1 DigitalLDOLogic_VIA1 $T=81070 57940 0 0 $X=80820 $Y=57710
X3560 3 DigitalLDOLogic_VIA1 $T=82910 11700 0 0 $X=82660 $Y=11470
X3561 3 DigitalLDOLogic_VIA1 $T=82910 15780 0 0 $X=82660 $Y=15550
X3562 3 DigitalLDOLogic_VIA1 $T=82910 19860 0 0 $X=82660 $Y=19630
X3563 3 DigitalLDOLogic_VIA1 $T=82910 23940 0 0 $X=82660 $Y=23710
X3564 3 DigitalLDOLogic_VIA1 $T=82910 28020 0 0 $X=82660 $Y=27790
X3565 3 DigitalLDOLogic_VIA1 $T=82910 32100 0 0 $X=82660 $Y=31870
X3566 3 DigitalLDOLogic_VIA1 $T=82910 36180 0 0 $X=82660 $Y=35950
X3567 3 DigitalLDOLogic_VIA1 $T=82910 40260 0 0 $X=82660 $Y=40030
X3568 3 DigitalLDOLogic_VIA1 $T=82910 44340 0 0 $X=82660 $Y=44110
X3569 3 DigitalLDOLogic_VIA1 $T=82910 48420 0 0 $X=82660 $Y=48190
X3570 3 DigitalLDOLogic_VIA1 $T=82910 52500 0 0 $X=82660 $Y=52270
X3571 3 DigitalLDOLogic_VIA1 $T=82910 56580 0 0 $X=82660 $Y=56350
X3572 1 DigitalLDOLogic_VIA1 $T=83830 13060 0 0 $X=83580 $Y=12830
X3573 1 DigitalLDOLogic_VIA1 $T=83830 17140 0 0 $X=83580 $Y=16910
X3574 1 DigitalLDOLogic_VIA1 $T=83830 21220 0 0 $X=83580 $Y=20990
X3575 1 DigitalLDOLogic_VIA1 $T=83830 25300 0 0 $X=83580 $Y=25070
X3576 1 DigitalLDOLogic_VIA1 $T=83830 29380 0 0 $X=83580 $Y=29150
X3577 1 DigitalLDOLogic_VIA1 $T=83830 33460 0 0 $X=83580 $Y=33230
X3578 1 DigitalLDOLogic_VIA1 $T=83830 37540 0 0 $X=83580 $Y=37310
X3579 1 DigitalLDOLogic_VIA1 $T=83830 41620 0 0 $X=83580 $Y=41390
X3580 1 DigitalLDOLogic_VIA1 $T=83830 45700 0 0 $X=83580 $Y=45470
X3581 1 DigitalLDOLogic_VIA1 $T=83830 49780 0 0 $X=83580 $Y=49550
X3582 1 DigitalLDOLogic_VIA1 $T=83830 53860 0 0 $X=83580 $Y=53630
X3583 1 DigitalLDOLogic_VIA1 $T=83830 57940 0 0 $X=83580 $Y=57710
X3584 3 DigitalLDOLogic_VIA1 $T=85670 11700 0 0 $X=85420 $Y=11470
X3585 3 DigitalLDOLogic_VIA1 $T=85670 15780 0 0 $X=85420 $Y=15550
X3586 3 DigitalLDOLogic_VIA1 $T=85670 19860 0 0 $X=85420 $Y=19630
X3587 3 DigitalLDOLogic_VIA1 $T=85670 23940 0 0 $X=85420 $Y=23710
X3588 3 DigitalLDOLogic_VIA1 $T=85670 28020 0 0 $X=85420 $Y=27790
X3589 3 DigitalLDOLogic_VIA1 $T=85670 32100 0 0 $X=85420 $Y=31870
X3590 3 DigitalLDOLogic_VIA1 $T=85670 36180 0 0 $X=85420 $Y=35950
X3591 3 DigitalLDOLogic_VIA1 $T=85670 40260 0 0 $X=85420 $Y=40030
X3592 3 DigitalLDOLogic_VIA1 $T=85670 44340 0 0 $X=85420 $Y=44110
X3593 3 DigitalLDOLogic_VIA1 $T=85670 48420 0 0 $X=85420 $Y=48190
X3594 3 DigitalLDOLogic_VIA1 $T=85670 52500 0 0 $X=85420 $Y=52270
X3595 3 DigitalLDOLogic_VIA1 $T=85670 56580 0 0 $X=85420 $Y=56350
X3596 1 DigitalLDOLogic_VIA1 $T=86590 13060 0 0 $X=86340 $Y=12830
X3597 1 DigitalLDOLogic_VIA1 $T=86590 17140 0 0 $X=86340 $Y=16910
X3598 1 DigitalLDOLogic_VIA1 $T=86590 21220 0 0 $X=86340 $Y=20990
X3599 1 DigitalLDOLogic_VIA1 $T=86590 25300 0 0 $X=86340 $Y=25070
X3600 1 DigitalLDOLogic_VIA1 $T=86590 29380 0 0 $X=86340 $Y=29150
X3601 1 DigitalLDOLogic_VIA1 $T=86590 33460 0 0 $X=86340 $Y=33230
X3602 1 DigitalLDOLogic_VIA1 $T=86590 37540 0 0 $X=86340 $Y=37310
X3603 1 DigitalLDOLogic_VIA1 $T=86590 41620 0 0 $X=86340 $Y=41390
X3604 1 DigitalLDOLogic_VIA1 $T=86590 45700 0 0 $X=86340 $Y=45470
X3605 1 DigitalLDOLogic_VIA1 $T=86590 49780 0 0 $X=86340 $Y=49550
X3606 1 DigitalLDOLogic_VIA1 $T=86590 53860 0 0 $X=86340 $Y=53630
X3607 1 DigitalLDOLogic_VIA1 $T=86590 57940 0 0 $X=86340 $Y=57710
X3608 3 DigitalLDOLogic_VIA1 $T=88430 11700 0 0 $X=88180 $Y=11470
X3609 3 DigitalLDOLogic_VIA1 $T=88430 15780 0 0 $X=88180 $Y=15550
X3610 3 DigitalLDOLogic_VIA1 $T=88430 19860 0 0 $X=88180 $Y=19630
X3611 3 DigitalLDOLogic_VIA1 $T=88430 23940 0 0 $X=88180 $Y=23710
X3612 3 DigitalLDOLogic_VIA1 $T=88430 28020 0 0 $X=88180 $Y=27790
X3613 3 DigitalLDOLogic_VIA1 $T=88430 32100 0 0 $X=88180 $Y=31870
X3614 3 DigitalLDOLogic_VIA1 $T=88430 36180 0 0 $X=88180 $Y=35950
X3615 3 DigitalLDOLogic_VIA1 $T=88430 40260 0 0 $X=88180 $Y=40030
X3616 3 DigitalLDOLogic_VIA1 $T=88430 44340 0 0 $X=88180 $Y=44110
X3617 3 DigitalLDOLogic_VIA1 $T=88430 48420 0 0 $X=88180 $Y=48190
X3618 3 DigitalLDOLogic_VIA1 $T=88430 52500 0 0 $X=88180 $Y=52270
X3619 3 DigitalLDOLogic_VIA1 $T=88430 56580 0 0 $X=88180 $Y=56350
X3620 1 DigitalLDOLogic_VIA1 $T=89350 13060 0 0 $X=89100 $Y=12830
X3621 1 DigitalLDOLogic_VIA1 $T=89350 17140 0 0 $X=89100 $Y=16910
X3622 1 DigitalLDOLogic_VIA1 $T=89350 21220 0 0 $X=89100 $Y=20990
X3623 1 DigitalLDOLogic_VIA1 $T=89350 25300 0 0 $X=89100 $Y=25070
X3624 1 DigitalLDOLogic_VIA1 $T=89350 29380 0 0 $X=89100 $Y=29150
X3625 1 DigitalLDOLogic_VIA1 $T=89350 33460 0 0 $X=89100 $Y=33230
X3626 1 DigitalLDOLogic_VIA1 $T=89350 37540 0 0 $X=89100 $Y=37310
X3627 1 DigitalLDOLogic_VIA1 $T=89350 41620 0 0 $X=89100 $Y=41390
X3628 1 DigitalLDOLogic_VIA1 $T=89350 45700 0 0 $X=89100 $Y=45470
X3629 1 DigitalLDOLogic_VIA1 $T=89350 49780 0 0 $X=89100 $Y=49550
X3630 1 DigitalLDOLogic_VIA1 $T=89350 53860 0 0 $X=89100 $Y=53630
X3631 1 DigitalLDOLogic_VIA1 $T=89350 57940 0 0 $X=89100 $Y=57710
X3632 3 DigitalLDOLogic_VIA1 $T=91190 11700 0 0 $X=90940 $Y=11470
X3633 3 DigitalLDOLogic_VIA1 $T=91190 15780 0 0 $X=90940 $Y=15550
X3634 3 DigitalLDOLogic_VIA1 $T=91190 19860 0 0 $X=90940 $Y=19630
X3635 3 DigitalLDOLogic_VIA1 $T=91190 23940 0 0 $X=90940 $Y=23710
X3636 3 DigitalLDOLogic_VIA1 $T=91190 28020 0 0 $X=90940 $Y=27790
X3637 3 DigitalLDOLogic_VIA1 $T=91190 32100 0 0 $X=90940 $Y=31870
X3638 3 DigitalLDOLogic_VIA1 $T=91190 36180 0 0 $X=90940 $Y=35950
X3639 3 DigitalLDOLogic_VIA1 $T=91190 40260 0 0 $X=90940 $Y=40030
X3640 3 DigitalLDOLogic_VIA1 $T=91190 44340 0 0 $X=90940 $Y=44110
X3641 3 DigitalLDOLogic_VIA1 $T=91190 48420 0 0 $X=90940 $Y=48190
X3642 3 DigitalLDOLogic_VIA1 $T=91190 52500 0 0 $X=90940 $Y=52270
X3643 3 DigitalLDOLogic_VIA1 $T=91190 56580 0 0 $X=90940 $Y=56350
X3644 1 DigitalLDOLogic_VIA1 $T=92110 13060 0 0 $X=91860 $Y=12830
X3645 1 DigitalLDOLogic_VIA1 $T=92110 17140 0 0 $X=91860 $Y=16910
X3646 1 DigitalLDOLogic_VIA1 $T=92110 21220 0 0 $X=91860 $Y=20990
X3647 1 DigitalLDOLogic_VIA1 $T=92110 25300 0 0 $X=91860 $Y=25070
X3648 1 DigitalLDOLogic_VIA1 $T=92110 29380 0 0 $X=91860 $Y=29150
X3649 1 DigitalLDOLogic_VIA1 $T=92110 33460 0 0 $X=91860 $Y=33230
X3650 1 DigitalLDOLogic_VIA1 $T=92110 37540 0 0 $X=91860 $Y=37310
X3651 1 DigitalLDOLogic_VIA1 $T=92110 41620 0 0 $X=91860 $Y=41390
X3652 1 DigitalLDOLogic_VIA1 $T=92110 45700 0 0 $X=91860 $Y=45470
X3653 1 DigitalLDOLogic_VIA1 $T=92110 49780 0 0 $X=91860 $Y=49550
X3654 1 DigitalLDOLogic_VIA1 $T=92110 53860 0 0 $X=91860 $Y=53630
X3655 1 DigitalLDOLogic_VIA1 $T=92110 57940 0 0 $X=91860 $Y=57710
X3656 3 DigitalLDOLogic_VIA1 $T=93950 11700 0 0 $X=93700 $Y=11470
X3657 3 DigitalLDOLogic_VIA1 $T=93950 15780 0 0 $X=93700 $Y=15550
X3658 3 DigitalLDOLogic_VIA1 $T=93950 19860 0 0 $X=93700 $Y=19630
X3659 3 DigitalLDOLogic_VIA1 $T=93950 23940 0 0 $X=93700 $Y=23710
X3660 3 DigitalLDOLogic_VIA1 $T=93950 28020 0 0 $X=93700 $Y=27790
X3661 3 DigitalLDOLogic_VIA1 $T=93950 32100 0 0 $X=93700 $Y=31870
X3662 3 DigitalLDOLogic_VIA1 $T=93950 36180 0 0 $X=93700 $Y=35950
X3663 3 DigitalLDOLogic_VIA1 $T=93950 40260 0 0 $X=93700 $Y=40030
X3664 3 DigitalLDOLogic_VIA1 $T=93950 44340 0 0 $X=93700 $Y=44110
X3665 3 DigitalLDOLogic_VIA1 $T=93950 48420 0 0 $X=93700 $Y=48190
X3666 3 DigitalLDOLogic_VIA1 $T=93950 52500 0 0 $X=93700 $Y=52270
X3667 3 DigitalLDOLogic_VIA1 $T=93950 56580 0 0 $X=93700 $Y=56350
X3668 1 DigitalLDOLogic_VIA1 $T=94870 13060 0 0 $X=94620 $Y=12830
X3669 1 DigitalLDOLogic_VIA1 $T=94870 17140 0 0 $X=94620 $Y=16910
X3670 1 DigitalLDOLogic_VIA1 $T=94870 21220 0 0 $X=94620 $Y=20990
X3671 1 DigitalLDOLogic_VIA1 $T=94870 25300 0 0 $X=94620 $Y=25070
X3672 1 DigitalLDOLogic_VIA1 $T=94870 29380 0 0 $X=94620 $Y=29150
X3673 1 DigitalLDOLogic_VIA1 $T=94870 33460 0 0 $X=94620 $Y=33230
X3674 1 DigitalLDOLogic_VIA1 $T=94870 37540 0 0 $X=94620 $Y=37310
X3675 1 DigitalLDOLogic_VIA1 $T=94870 41620 0 0 $X=94620 $Y=41390
X3676 1 DigitalLDOLogic_VIA1 $T=94870 45700 0 0 $X=94620 $Y=45470
X3677 1 DigitalLDOLogic_VIA1 $T=94870 49780 0 0 $X=94620 $Y=49550
X3678 1 DigitalLDOLogic_VIA1 $T=94870 53860 0 0 $X=94620 $Y=53630
X3679 1 DigitalLDOLogic_VIA1 $T=94870 57940 0 0 $X=94620 $Y=57710
X3680 3 DigitalLDOLogic_VIA1 $T=96710 11700 0 0 $X=96460 $Y=11470
X3681 3 DigitalLDOLogic_VIA1 $T=96710 15780 0 0 $X=96460 $Y=15550
X3682 3 DigitalLDOLogic_VIA1 $T=96710 19860 0 0 $X=96460 $Y=19630
X3683 3 DigitalLDOLogic_VIA1 $T=96710 23940 0 0 $X=96460 $Y=23710
X3684 3 DigitalLDOLogic_VIA1 $T=96710 28020 0 0 $X=96460 $Y=27790
X3685 3 DigitalLDOLogic_VIA1 $T=96710 32100 0 0 $X=96460 $Y=31870
X3686 3 DigitalLDOLogic_VIA1 $T=96710 36180 0 0 $X=96460 $Y=35950
X3687 3 DigitalLDOLogic_VIA1 $T=96710 40260 0 0 $X=96460 $Y=40030
X3688 3 DigitalLDOLogic_VIA1 $T=96710 44340 0 0 $X=96460 $Y=44110
X3689 3 DigitalLDOLogic_VIA1 $T=96710 48420 0 0 $X=96460 $Y=48190
X3690 3 DigitalLDOLogic_VIA1 $T=96710 52500 0 0 $X=96460 $Y=52270
X3691 3 DigitalLDOLogic_VIA1 $T=96710 56580 0 0 $X=96460 $Y=56350
X3692 1 DigitalLDOLogic_VIA1 $T=97630 13060 0 0 $X=97380 $Y=12830
X3693 1 DigitalLDOLogic_VIA1 $T=97630 17140 0 0 $X=97380 $Y=16910
X3694 1 DigitalLDOLogic_VIA1 $T=97630 21220 0 0 $X=97380 $Y=20990
X3695 1 DigitalLDOLogic_VIA1 $T=97630 25300 0 0 $X=97380 $Y=25070
X3696 1 DigitalLDOLogic_VIA1 $T=97630 29380 0 0 $X=97380 $Y=29150
X3697 1 DigitalLDOLogic_VIA1 $T=97630 33460 0 0 $X=97380 $Y=33230
X3698 1 DigitalLDOLogic_VIA1 $T=97630 37540 0 0 $X=97380 $Y=37310
X3699 1 DigitalLDOLogic_VIA1 $T=97630 41620 0 0 $X=97380 $Y=41390
X3700 1 DigitalLDOLogic_VIA1 $T=97630 45700 0 0 $X=97380 $Y=45470
X3701 1 DigitalLDOLogic_VIA1 $T=97630 49780 0 0 $X=97380 $Y=49550
X3702 1 DigitalLDOLogic_VIA1 $T=97630 53860 0 0 $X=97380 $Y=53630
X3703 1 DigitalLDOLogic_VIA1 $T=97630 57940 0 0 $X=97380 $Y=57710
X3704 3 DigitalLDOLogic_VIA1 $T=99470 11700 0 0 $X=99220 $Y=11470
X3705 3 DigitalLDOLogic_VIA1 $T=99470 15780 0 0 $X=99220 $Y=15550
X3706 3 DigitalLDOLogic_VIA1 $T=99470 19860 0 0 $X=99220 $Y=19630
X3707 3 DigitalLDOLogic_VIA1 $T=99470 23940 0 0 $X=99220 $Y=23710
X3708 3 DigitalLDOLogic_VIA1 $T=99470 28020 0 0 $X=99220 $Y=27790
X3709 3 DigitalLDOLogic_VIA1 $T=99470 32100 0 0 $X=99220 $Y=31870
X3710 3 DigitalLDOLogic_VIA1 $T=99470 36180 0 0 $X=99220 $Y=35950
X3711 3 DigitalLDOLogic_VIA1 $T=99470 40260 0 0 $X=99220 $Y=40030
X3712 3 DigitalLDOLogic_VIA1 $T=99470 44340 0 0 $X=99220 $Y=44110
X3713 3 DigitalLDOLogic_VIA1 $T=99470 48420 0 0 $X=99220 $Y=48190
X3714 3 DigitalLDOLogic_VIA1 $T=99470 52500 0 0 $X=99220 $Y=52270
X3715 3 DigitalLDOLogic_VIA1 $T=99470 56580 0 0 $X=99220 $Y=56350
X3716 1 DigitalLDOLogic_VIA1 $T=100390 13060 0 0 $X=100140 $Y=12830
X3717 1 DigitalLDOLogic_VIA1 $T=100390 17140 0 0 $X=100140 $Y=16910
X3718 1 DigitalLDOLogic_VIA1 $T=100390 21220 0 0 $X=100140 $Y=20990
X3719 1 DigitalLDOLogic_VIA1 $T=100390 25300 0 0 $X=100140 $Y=25070
X3720 1 DigitalLDOLogic_VIA1 $T=100390 29380 0 0 $X=100140 $Y=29150
X3721 1 DigitalLDOLogic_VIA1 $T=100390 33460 0 0 $X=100140 $Y=33230
X3722 1 DigitalLDOLogic_VIA1 $T=100390 37540 0 0 $X=100140 $Y=37310
X3723 1 DigitalLDOLogic_VIA1 $T=100390 41620 0 0 $X=100140 $Y=41390
X3724 1 DigitalLDOLogic_VIA1 $T=100390 45700 0 0 $X=100140 $Y=45470
X3725 1 DigitalLDOLogic_VIA1 $T=100390 49780 0 0 $X=100140 $Y=49550
X3726 1 DigitalLDOLogic_VIA1 $T=100390 53860 0 0 $X=100140 $Y=53630
X3727 1 DigitalLDOLogic_VIA1 $T=100390 57940 0 0 $X=100140 $Y=57710
X3728 3 DigitalLDOLogic_VIA1 $T=102230 11700 0 0 $X=101980 $Y=11470
X3729 3 DigitalLDOLogic_VIA1 $T=102230 15780 0 0 $X=101980 $Y=15550
X3730 3 DigitalLDOLogic_VIA1 $T=102230 19860 0 0 $X=101980 $Y=19630
X3731 3 DigitalLDOLogic_VIA1 $T=102230 23940 0 0 $X=101980 $Y=23710
X3732 3 DigitalLDOLogic_VIA1 $T=102230 28020 0 0 $X=101980 $Y=27790
X3733 3 DigitalLDOLogic_VIA1 $T=102230 32100 0 0 $X=101980 $Y=31870
X3734 3 DigitalLDOLogic_VIA1 $T=102230 36180 0 0 $X=101980 $Y=35950
X3735 3 DigitalLDOLogic_VIA1 $T=102230 40260 0 0 $X=101980 $Y=40030
X3736 3 DigitalLDOLogic_VIA1 $T=102230 44340 0 0 $X=101980 $Y=44110
X3737 3 DigitalLDOLogic_VIA1 $T=102230 48420 0 0 $X=101980 $Y=48190
X3738 3 DigitalLDOLogic_VIA1 $T=102230 52500 0 0 $X=101980 $Y=52270
X3739 3 DigitalLDOLogic_VIA1 $T=102230 56580 0 0 $X=101980 $Y=56350
X3740 1 DigitalLDOLogic_VIA1 $T=103150 13060 0 0 $X=102900 $Y=12830
X3741 1 DigitalLDOLogic_VIA1 $T=103150 17140 0 0 $X=102900 $Y=16910
X3742 1 DigitalLDOLogic_VIA1 $T=103150 21220 0 0 $X=102900 $Y=20990
X3743 1 DigitalLDOLogic_VIA1 $T=103150 25300 0 0 $X=102900 $Y=25070
X3744 1 DigitalLDOLogic_VIA1 $T=103150 29380 0 0 $X=102900 $Y=29150
X3745 1 DigitalLDOLogic_VIA1 $T=103150 33460 0 0 $X=102900 $Y=33230
X3746 1 DigitalLDOLogic_VIA1 $T=103150 37540 0 0 $X=102900 $Y=37310
X3747 1 DigitalLDOLogic_VIA1 $T=103150 41620 0 0 $X=102900 $Y=41390
X3748 1 DigitalLDOLogic_VIA1 $T=103150 45700 0 0 $X=102900 $Y=45470
X3749 1 DigitalLDOLogic_VIA1 $T=103150 49780 0 0 $X=102900 $Y=49550
X3750 1 DigitalLDOLogic_VIA1 $T=103150 53860 0 0 $X=102900 $Y=53630
X3751 1 DigitalLDOLogic_VIA1 $T=103150 57940 0 0 $X=102900 $Y=57710
X3752 3 DigitalLDOLogic_VIA1 $T=104990 11700 0 0 $X=104740 $Y=11470
X3753 3 DigitalLDOLogic_VIA1 $T=104990 15780 0 0 $X=104740 $Y=15550
X3754 3 DigitalLDOLogic_VIA1 $T=104990 19860 0 0 $X=104740 $Y=19630
X3755 3 DigitalLDOLogic_VIA1 $T=104990 23940 0 0 $X=104740 $Y=23710
X3756 3 DigitalLDOLogic_VIA1 $T=104990 28020 0 0 $X=104740 $Y=27790
X3757 3 DigitalLDOLogic_VIA1 $T=104990 32100 0 0 $X=104740 $Y=31870
X3758 3 DigitalLDOLogic_VIA1 $T=104990 36180 0 0 $X=104740 $Y=35950
X3759 3 DigitalLDOLogic_VIA1 $T=104990 40260 0 0 $X=104740 $Y=40030
X3760 3 DigitalLDOLogic_VIA1 $T=104990 44340 0 0 $X=104740 $Y=44110
X3761 3 DigitalLDOLogic_VIA1 $T=104990 48420 0 0 $X=104740 $Y=48190
X3762 3 DigitalLDOLogic_VIA1 $T=104990 52500 0 0 $X=104740 $Y=52270
X3763 3 DigitalLDOLogic_VIA1 $T=104990 56580 0 0 $X=104740 $Y=56350
X3764 1 DigitalLDOLogic_VIA1 $T=105910 13060 0 0 $X=105660 $Y=12830
X3765 1 DigitalLDOLogic_VIA1 $T=105910 17140 0 0 $X=105660 $Y=16910
X3766 1 DigitalLDOLogic_VIA1 $T=105910 21220 0 0 $X=105660 $Y=20990
X3767 1 DigitalLDOLogic_VIA1 $T=105910 25300 0 0 $X=105660 $Y=25070
X3768 1 DigitalLDOLogic_VIA1 $T=105910 29380 0 0 $X=105660 $Y=29150
X3769 1 DigitalLDOLogic_VIA1 $T=105910 33460 0 0 $X=105660 $Y=33230
X3770 1 DigitalLDOLogic_VIA1 $T=105910 37540 0 0 $X=105660 $Y=37310
X3771 1 DigitalLDOLogic_VIA1 $T=105910 41620 0 0 $X=105660 $Y=41390
X3772 1 DigitalLDOLogic_VIA1 $T=105910 45700 0 0 $X=105660 $Y=45470
X3773 1 DigitalLDOLogic_VIA1 $T=105910 49780 0 0 $X=105660 $Y=49550
X3774 1 DigitalLDOLogic_VIA1 $T=105910 53860 0 0 $X=105660 $Y=53630
X3775 1 DigitalLDOLogic_VIA1 $T=105910 57940 0 0 $X=105660 $Y=57710
X3776 3 DigitalLDOLogic_VIA1 $T=107750 11700 0 0 $X=107500 $Y=11470
X3777 3 DigitalLDOLogic_VIA1 $T=107750 15780 0 0 $X=107500 $Y=15550
X3778 3 DigitalLDOLogic_VIA1 $T=107750 19860 0 0 $X=107500 $Y=19630
X3779 3 DigitalLDOLogic_VIA1 $T=107750 23940 0 0 $X=107500 $Y=23710
X3780 3 DigitalLDOLogic_VIA1 $T=107750 28020 0 0 $X=107500 $Y=27790
X3781 3 DigitalLDOLogic_VIA1 $T=107750 32100 0 0 $X=107500 $Y=31870
X3782 3 DigitalLDOLogic_VIA1 $T=107750 36180 0 0 $X=107500 $Y=35950
X3783 3 DigitalLDOLogic_VIA1 $T=107750 40260 0 0 $X=107500 $Y=40030
X3784 3 DigitalLDOLogic_VIA1 $T=107750 44340 0 0 $X=107500 $Y=44110
X3785 3 DigitalLDOLogic_VIA1 $T=107750 48420 0 0 $X=107500 $Y=48190
X3786 3 DigitalLDOLogic_VIA1 $T=107750 52500 0 0 $X=107500 $Y=52270
X3787 3 DigitalLDOLogic_VIA1 $T=107750 56580 0 0 $X=107500 $Y=56350
X3788 1 DigitalLDOLogic_VIA1 $T=108670 13060 0 0 $X=108420 $Y=12830
X3789 1 DigitalLDOLogic_VIA1 $T=108670 17140 0 0 $X=108420 $Y=16910
X3790 1 DigitalLDOLogic_VIA1 $T=108670 21220 0 0 $X=108420 $Y=20990
X3791 1 DigitalLDOLogic_VIA1 $T=108670 25300 0 0 $X=108420 $Y=25070
X3792 1 DigitalLDOLogic_VIA1 $T=108670 29380 0 0 $X=108420 $Y=29150
X3793 1 DigitalLDOLogic_VIA1 $T=108670 33460 0 0 $X=108420 $Y=33230
X3794 1 DigitalLDOLogic_VIA1 $T=108670 37540 0 0 $X=108420 $Y=37310
X3795 1 DigitalLDOLogic_VIA1 $T=108670 41620 0 0 $X=108420 $Y=41390
X3796 1 DigitalLDOLogic_VIA1 $T=108670 45700 0 0 $X=108420 $Y=45470
X3797 1 DigitalLDOLogic_VIA1 $T=108670 49780 0 0 $X=108420 $Y=49550
X3798 1 DigitalLDOLogic_VIA1 $T=108670 53860 0 0 $X=108420 $Y=53630
X3799 1 DigitalLDOLogic_VIA1 $T=108670 57940 0 0 $X=108420 $Y=57710
X3800 3 DigitalLDOLogic_VIA1 $T=110510 11700 0 0 $X=110260 $Y=11470
X3801 3 DigitalLDOLogic_VIA1 $T=110510 15780 0 0 $X=110260 $Y=15550
X3802 3 DigitalLDOLogic_VIA1 $T=110510 19860 0 0 $X=110260 $Y=19630
X3803 3 DigitalLDOLogic_VIA1 $T=110510 23940 0 0 $X=110260 $Y=23710
X3804 3 DigitalLDOLogic_VIA1 $T=110510 28020 0 0 $X=110260 $Y=27790
X3805 3 DigitalLDOLogic_VIA1 $T=110510 32100 0 0 $X=110260 $Y=31870
X3806 3 DigitalLDOLogic_VIA1 $T=110510 36180 0 0 $X=110260 $Y=35950
X3807 3 DigitalLDOLogic_VIA1 $T=110510 40260 0 0 $X=110260 $Y=40030
X3808 3 DigitalLDOLogic_VIA1 $T=110510 44340 0 0 $X=110260 $Y=44110
X3809 3 DigitalLDOLogic_VIA1 $T=110510 48420 0 0 $X=110260 $Y=48190
X3810 3 DigitalLDOLogic_VIA1 $T=110510 52500 0 0 $X=110260 $Y=52270
X3811 3 DigitalLDOLogic_VIA1 $T=110510 56580 0 0 $X=110260 $Y=56350
X3812 1 DigitalLDOLogic_VIA1 $T=111430 13060 0 0 $X=111180 $Y=12830
X3813 1 DigitalLDOLogic_VIA1 $T=111430 17140 0 0 $X=111180 $Y=16910
X3814 1 DigitalLDOLogic_VIA1 $T=111430 21220 0 0 $X=111180 $Y=20990
X3815 1 DigitalLDOLogic_VIA1 $T=111430 25300 0 0 $X=111180 $Y=25070
X3816 1 DigitalLDOLogic_VIA1 $T=111430 29380 0 0 $X=111180 $Y=29150
X3817 1 DigitalLDOLogic_VIA1 $T=111430 33460 0 0 $X=111180 $Y=33230
X3818 1 DigitalLDOLogic_VIA1 $T=111430 37540 0 0 $X=111180 $Y=37310
X3819 1 DigitalLDOLogic_VIA1 $T=111430 41620 0 0 $X=111180 $Y=41390
X3820 1 DigitalLDOLogic_VIA1 $T=111430 45700 0 0 $X=111180 $Y=45470
X3821 1 DigitalLDOLogic_VIA1 $T=111430 49780 0 0 $X=111180 $Y=49550
X3822 1 DigitalLDOLogic_VIA1 $T=111430 53860 0 0 $X=111180 $Y=53630
X3823 1 DigitalLDOLogic_VIA1 $T=111430 57940 0 0 $X=111180 $Y=57710
X3824 3 DigitalLDOLogic_VIA1 $T=113270 11700 0 0 $X=113020 $Y=11470
X3825 3 DigitalLDOLogic_VIA1 $T=113270 15780 0 0 $X=113020 $Y=15550
X3826 3 DigitalLDOLogic_VIA1 $T=113270 19860 0 0 $X=113020 $Y=19630
X3827 3 DigitalLDOLogic_VIA1 $T=113270 23940 0 0 $X=113020 $Y=23710
X3828 3 DigitalLDOLogic_VIA1 $T=113270 28020 0 0 $X=113020 $Y=27790
X3829 3 DigitalLDOLogic_VIA1 $T=113270 32100 0 0 $X=113020 $Y=31870
X3830 3 DigitalLDOLogic_VIA1 $T=113270 36180 0 0 $X=113020 $Y=35950
X3831 3 DigitalLDOLogic_VIA1 $T=113270 40260 0 0 $X=113020 $Y=40030
X3832 3 DigitalLDOLogic_VIA1 $T=113270 44340 0 0 $X=113020 $Y=44110
X3833 3 DigitalLDOLogic_VIA1 $T=113270 48420 0 0 $X=113020 $Y=48190
X3834 3 DigitalLDOLogic_VIA1 $T=113270 52500 0 0 $X=113020 $Y=52270
X3835 3 DigitalLDOLogic_VIA1 $T=113270 56580 0 0 $X=113020 $Y=56350
X3836 1 DigitalLDOLogic_VIA1 $T=114190 13060 0 0 $X=113940 $Y=12830
X3837 1 DigitalLDOLogic_VIA1 $T=114190 17140 0 0 $X=113940 $Y=16910
X3838 1 DigitalLDOLogic_VIA1 $T=114190 21220 0 0 $X=113940 $Y=20990
X3839 1 DigitalLDOLogic_VIA1 $T=114190 25300 0 0 $X=113940 $Y=25070
X3840 1 DigitalLDOLogic_VIA1 $T=114190 29380 0 0 $X=113940 $Y=29150
X3841 1 DigitalLDOLogic_VIA1 $T=114190 33460 0 0 $X=113940 $Y=33230
X3842 1 DigitalLDOLogic_VIA1 $T=114190 37540 0 0 $X=113940 $Y=37310
X3843 1 DigitalLDOLogic_VIA1 $T=114190 41620 0 0 $X=113940 $Y=41390
X3844 1 DigitalLDOLogic_VIA1 $T=114190 45700 0 0 $X=113940 $Y=45470
X3845 1 DigitalLDOLogic_VIA1 $T=114190 49780 0 0 $X=113940 $Y=49550
X3846 1 DigitalLDOLogic_VIA1 $T=114190 53860 0 0 $X=113940 $Y=53630
X3847 1 DigitalLDOLogic_VIA1 $T=114190 57940 0 0 $X=113940 $Y=57710
X3848 3 DigitalLDOLogic_VIA1 $T=116030 11700 0 0 $X=115780 $Y=11470
X3849 3 DigitalLDOLogic_VIA1 $T=116030 15780 0 0 $X=115780 $Y=15550
X3850 3 DigitalLDOLogic_VIA1 $T=116030 19860 0 0 $X=115780 $Y=19630
X3851 3 DigitalLDOLogic_VIA1 $T=116030 23940 0 0 $X=115780 $Y=23710
X3852 3 DigitalLDOLogic_VIA1 $T=116030 28020 0 0 $X=115780 $Y=27790
X3853 3 DigitalLDOLogic_VIA1 $T=116030 32100 0 0 $X=115780 $Y=31870
X3854 3 DigitalLDOLogic_VIA1 $T=116030 36180 0 0 $X=115780 $Y=35950
X3855 3 DigitalLDOLogic_VIA1 $T=116030 40260 0 0 $X=115780 $Y=40030
X3856 3 DigitalLDOLogic_VIA1 $T=116030 44340 0 0 $X=115780 $Y=44110
X3857 3 DigitalLDOLogic_VIA1 $T=116030 48420 0 0 $X=115780 $Y=48190
X3858 3 DigitalLDOLogic_VIA1 $T=116030 52500 0 0 $X=115780 $Y=52270
X3859 3 DigitalLDOLogic_VIA1 $T=116030 56580 0 0 $X=115780 $Y=56350
X3860 1 DigitalLDOLogic_VIA1 $T=116950 13060 0 0 $X=116700 $Y=12830
X3861 1 DigitalLDOLogic_VIA1 $T=116950 17140 0 0 $X=116700 $Y=16910
X3862 1 DigitalLDOLogic_VIA1 $T=116950 21220 0 0 $X=116700 $Y=20990
X3863 1 DigitalLDOLogic_VIA1 $T=116950 25300 0 0 $X=116700 $Y=25070
X3864 1 DigitalLDOLogic_VIA1 $T=116950 29380 0 0 $X=116700 $Y=29150
X3865 1 DigitalLDOLogic_VIA1 $T=116950 33460 0 0 $X=116700 $Y=33230
X3866 1 DigitalLDOLogic_VIA1 $T=116950 37540 0 0 $X=116700 $Y=37310
X3867 1 DigitalLDOLogic_VIA1 $T=116950 41620 0 0 $X=116700 $Y=41390
X3868 1 DigitalLDOLogic_VIA1 $T=116950 45700 0 0 $X=116700 $Y=45470
X3869 1 DigitalLDOLogic_VIA1 $T=116950 49780 0 0 $X=116700 $Y=49550
X3870 1 DigitalLDOLogic_VIA1 $T=116950 53860 0 0 $X=116700 $Y=53630
X3871 1 DigitalLDOLogic_VIA1 $T=116950 57940 0 0 $X=116700 $Y=57710
X3872 3 DigitalLDOLogic_VIA1 $T=118790 11700 0 0 $X=118540 $Y=11470
X3873 3 DigitalLDOLogic_VIA1 $T=118790 15780 0 0 $X=118540 $Y=15550
X3874 3 DigitalLDOLogic_VIA1 $T=118790 19860 0 0 $X=118540 $Y=19630
X3875 3 DigitalLDOLogic_VIA1 $T=118790 23940 0 0 $X=118540 $Y=23710
X3876 3 DigitalLDOLogic_VIA1 $T=118790 28020 0 0 $X=118540 $Y=27790
X3877 3 DigitalLDOLogic_VIA1 $T=118790 32100 0 0 $X=118540 $Y=31870
X3878 3 DigitalLDOLogic_VIA1 $T=118790 36180 0 0 $X=118540 $Y=35950
X3879 3 DigitalLDOLogic_VIA1 $T=118790 40260 0 0 $X=118540 $Y=40030
X3880 3 DigitalLDOLogic_VIA1 $T=118790 44340 0 0 $X=118540 $Y=44110
X3881 3 DigitalLDOLogic_VIA1 $T=118790 48420 0 0 $X=118540 $Y=48190
X3882 3 DigitalLDOLogic_VIA1 $T=118790 52500 0 0 $X=118540 $Y=52270
X3883 3 DigitalLDOLogic_VIA1 $T=118790 56580 0 0 $X=118540 $Y=56350
X3884 1 DigitalLDOLogic_VIA1 $T=119710 13060 0 0 $X=119460 $Y=12830
X3885 1 DigitalLDOLogic_VIA1 $T=119710 17140 0 0 $X=119460 $Y=16910
X3886 1 DigitalLDOLogic_VIA1 $T=119710 21220 0 0 $X=119460 $Y=20990
X3887 1 DigitalLDOLogic_VIA1 $T=119710 25300 0 0 $X=119460 $Y=25070
X3888 1 DigitalLDOLogic_VIA1 $T=119710 29380 0 0 $X=119460 $Y=29150
X3889 1 DigitalLDOLogic_VIA1 $T=119710 33460 0 0 $X=119460 $Y=33230
X3890 1 DigitalLDOLogic_VIA1 $T=119710 37540 0 0 $X=119460 $Y=37310
X3891 1 DigitalLDOLogic_VIA1 $T=119710 41620 0 0 $X=119460 $Y=41390
X3892 1 DigitalLDOLogic_VIA1 $T=119710 45700 0 0 $X=119460 $Y=45470
X3893 1 DigitalLDOLogic_VIA1 $T=119710 49780 0 0 $X=119460 $Y=49550
X3894 1 DigitalLDOLogic_VIA1 $T=119710 53860 0 0 $X=119460 $Y=53630
X3895 1 DigitalLDOLogic_VIA1 $T=119710 57940 0 0 $X=119460 $Y=57710
X3896 3 DigitalLDOLogic_VIA1 $T=121550 11700 0 0 $X=121300 $Y=11470
X3897 3 DigitalLDOLogic_VIA1 $T=121550 15780 0 0 $X=121300 $Y=15550
X3898 3 DigitalLDOLogic_VIA1 $T=121550 19860 0 0 $X=121300 $Y=19630
X3899 3 DigitalLDOLogic_VIA1 $T=121550 23940 0 0 $X=121300 $Y=23710
X3900 3 DigitalLDOLogic_VIA1 $T=121550 28020 0 0 $X=121300 $Y=27790
X3901 3 DigitalLDOLogic_VIA1 $T=121550 32100 0 0 $X=121300 $Y=31870
X3902 3 DigitalLDOLogic_VIA1 $T=121550 36180 0 0 $X=121300 $Y=35950
X3903 3 DigitalLDOLogic_VIA1 $T=121550 40260 0 0 $X=121300 $Y=40030
X3904 3 DigitalLDOLogic_VIA1 $T=121550 44340 0 0 $X=121300 $Y=44110
X3905 3 DigitalLDOLogic_VIA1 $T=121550 48420 0 0 $X=121300 $Y=48190
X3906 3 DigitalLDOLogic_VIA1 $T=121550 52500 0 0 $X=121300 $Y=52270
X3907 3 DigitalLDOLogic_VIA1 $T=121550 56580 0 0 $X=121300 $Y=56350
X3908 1 DigitalLDOLogic_VIA1 $T=122470 13060 0 0 $X=122220 $Y=12830
X3909 1 DigitalLDOLogic_VIA1 $T=122470 17140 0 0 $X=122220 $Y=16910
X3910 1 DigitalLDOLogic_VIA1 $T=122470 21220 0 0 $X=122220 $Y=20990
X3911 1 DigitalLDOLogic_VIA1 $T=122470 25300 0 0 $X=122220 $Y=25070
X3912 1 DigitalLDOLogic_VIA1 $T=122470 29380 0 0 $X=122220 $Y=29150
X3913 1 DigitalLDOLogic_VIA1 $T=122470 33460 0 0 $X=122220 $Y=33230
X3914 1 DigitalLDOLogic_VIA1 $T=122470 37540 0 0 $X=122220 $Y=37310
X3915 1 DigitalLDOLogic_VIA1 $T=122470 41620 0 0 $X=122220 $Y=41390
X3916 1 DigitalLDOLogic_VIA1 $T=122470 45700 0 0 $X=122220 $Y=45470
X3917 1 DigitalLDOLogic_VIA1 $T=122470 49780 0 0 $X=122220 $Y=49550
X3918 1 DigitalLDOLogic_VIA1 $T=122470 53860 0 0 $X=122220 $Y=53630
X3919 1 DigitalLDOLogic_VIA1 $T=122470 57940 0 0 $X=122220 $Y=57710
X3920 3 DigitalLDOLogic_VIA1 $T=124310 11700 0 0 $X=124060 $Y=11470
X3921 3 DigitalLDOLogic_VIA1 $T=124310 15780 0 0 $X=124060 $Y=15550
X3922 3 DigitalLDOLogic_VIA1 $T=124310 19860 0 0 $X=124060 $Y=19630
X3923 3 DigitalLDOLogic_VIA1 $T=124310 23940 0 0 $X=124060 $Y=23710
X3924 3 DigitalLDOLogic_VIA1 $T=124310 28020 0 0 $X=124060 $Y=27790
X3925 3 DigitalLDOLogic_VIA1 $T=124310 32100 0 0 $X=124060 $Y=31870
X3926 3 DigitalLDOLogic_VIA1 $T=124310 36180 0 0 $X=124060 $Y=35950
X3927 3 DigitalLDOLogic_VIA1 $T=124310 40260 0 0 $X=124060 $Y=40030
X3928 3 DigitalLDOLogic_VIA1 $T=124310 44340 0 0 $X=124060 $Y=44110
X3929 3 DigitalLDOLogic_VIA1 $T=124310 48420 0 0 $X=124060 $Y=48190
X3930 3 DigitalLDOLogic_VIA1 $T=124310 52500 0 0 $X=124060 $Y=52270
X3931 3 DigitalLDOLogic_VIA1 $T=124310 56580 0 0 $X=124060 $Y=56350
X3932 1 DigitalLDOLogic_VIA1 $T=125230 13060 0 0 $X=124980 $Y=12830
X3933 1 DigitalLDOLogic_VIA1 $T=125230 17140 0 0 $X=124980 $Y=16910
X3934 1 DigitalLDOLogic_VIA1 $T=125230 21220 0 0 $X=124980 $Y=20990
X3935 1 DigitalLDOLogic_VIA1 $T=125230 25300 0 0 $X=124980 $Y=25070
X3936 1 DigitalLDOLogic_VIA1 $T=125230 29380 0 0 $X=124980 $Y=29150
X3937 1 DigitalLDOLogic_VIA1 $T=125230 33460 0 0 $X=124980 $Y=33230
X3938 1 DigitalLDOLogic_VIA1 $T=125230 37540 0 0 $X=124980 $Y=37310
X3939 1 DigitalLDOLogic_VIA1 $T=125230 41620 0 0 $X=124980 $Y=41390
X3940 1 DigitalLDOLogic_VIA1 $T=125230 45700 0 0 $X=124980 $Y=45470
X3941 1 DigitalLDOLogic_VIA1 $T=125230 49780 0 0 $X=124980 $Y=49550
X3942 1 DigitalLDOLogic_VIA1 $T=125230 53860 0 0 $X=124980 $Y=53630
X3943 1 DigitalLDOLogic_VIA1 $T=125230 57940 0 0 $X=124980 $Y=57710
X3944 3 DigitalLDOLogic_VIA1 $T=127070 11700 0 0 $X=126820 $Y=11470
X3945 3 DigitalLDOLogic_VIA1 $T=127070 15780 0 0 $X=126820 $Y=15550
X3946 3 DigitalLDOLogic_VIA1 $T=127070 19860 0 0 $X=126820 $Y=19630
X3947 3 DigitalLDOLogic_VIA1 $T=127070 23940 0 0 $X=126820 $Y=23710
X3948 3 DigitalLDOLogic_VIA1 $T=127070 28020 0 0 $X=126820 $Y=27790
X3949 3 DigitalLDOLogic_VIA1 $T=127070 32100 0 0 $X=126820 $Y=31870
X3950 3 DigitalLDOLogic_VIA1 $T=127070 36180 0 0 $X=126820 $Y=35950
X3951 3 DigitalLDOLogic_VIA1 $T=127070 40260 0 0 $X=126820 $Y=40030
X3952 3 DigitalLDOLogic_VIA1 $T=127070 44340 0 0 $X=126820 $Y=44110
X3953 3 DigitalLDOLogic_VIA1 $T=127070 48420 0 0 $X=126820 $Y=48190
X3954 3 DigitalLDOLogic_VIA1 $T=127070 52500 0 0 $X=126820 $Y=52270
X3955 3 DigitalLDOLogic_VIA1 $T=127070 56580 0 0 $X=126820 $Y=56350
X3956 1 DigitalLDOLogic_VIA1 $T=127990 13060 0 0 $X=127740 $Y=12830
X3957 1 DigitalLDOLogic_VIA1 $T=127990 17140 0 0 $X=127740 $Y=16910
X3958 1 DigitalLDOLogic_VIA1 $T=127990 21220 0 0 $X=127740 $Y=20990
X3959 1 DigitalLDOLogic_VIA1 $T=127990 25300 0 0 $X=127740 $Y=25070
X3960 1 DigitalLDOLogic_VIA1 $T=127990 29380 0 0 $X=127740 $Y=29150
X3961 1 DigitalLDOLogic_VIA1 $T=127990 33460 0 0 $X=127740 $Y=33230
X3962 1 DigitalLDOLogic_VIA1 $T=127990 37540 0 0 $X=127740 $Y=37310
X3963 1 DigitalLDOLogic_VIA1 $T=127990 41620 0 0 $X=127740 $Y=41390
X3964 1 DigitalLDOLogic_VIA1 $T=127990 45700 0 0 $X=127740 $Y=45470
X3965 1 DigitalLDOLogic_VIA1 $T=127990 49780 0 0 $X=127740 $Y=49550
X3966 1 DigitalLDOLogic_VIA1 $T=127990 53860 0 0 $X=127740 $Y=53630
X3967 1 DigitalLDOLogic_VIA1 $T=127990 57940 0 0 $X=127740 $Y=57710
X3968 3 DigitalLDOLogic_VIA1 $T=129830 11700 0 0 $X=129580 $Y=11470
X3969 3 DigitalLDOLogic_VIA1 $T=129830 15780 0 0 $X=129580 $Y=15550
X3970 3 DigitalLDOLogic_VIA1 $T=129830 19860 0 0 $X=129580 $Y=19630
X3971 3 DigitalLDOLogic_VIA1 $T=129830 23940 0 0 $X=129580 $Y=23710
X3972 3 DigitalLDOLogic_VIA1 $T=129830 28020 0 0 $X=129580 $Y=27790
X3973 3 DigitalLDOLogic_VIA1 $T=129830 32100 0 0 $X=129580 $Y=31870
X3974 3 DigitalLDOLogic_VIA1 $T=129830 36180 0 0 $X=129580 $Y=35950
X3975 3 DigitalLDOLogic_VIA1 $T=129830 40260 0 0 $X=129580 $Y=40030
X3976 3 DigitalLDOLogic_VIA1 $T=129830 44340 0 0 $X=129580 $Y=44110
X3977 3 DigitalLDOLogic_VIA1 $T=129830 48420 0 0 $X=129580 $Y=48190
X3978 3 DigitalLDOLogic_VIA1 $T=129830 52500 0 0 $X=129580 $Y=52270
X3979 3 DigitalLDOLogic_VIA1 $T=129830 56580 0 0 $X=129580 $Y=56350
X3980 1 DigitalLDOLogic_VIA1 $T=130750 13060 0 0 $X=130500 $Y=12830
X3981 1 DigitalLDOLogic_VIA1 $T=130750 17140 0 0 $X=130500 $Y=16910
X3982 1 DigitalLDOLogic_VIA1 $T=130750 21220 0 0 $X=130500 $Y=20990
X3983 1 DigitalLDOLogic_VIA1 $T=130750 25300 0 0 $X=130500 $Y=25070
X3984 1 DigitalLDOLogic_VIA1 $T=130750 29380 0 0 $X=130500 $Y=29150
X3985 1 DigitalLDOLogic_VIA1 $T=130750 33460 0 0 $X=130500 $Y=33230
X3986 1 DigitalLDOLogic_VIA1 $T=130750 37540 0 0 $X=130500 $Y=37310
X3987 1 DigitalLDOLogic_VIA1 $T=130750 41620 0 0 $X=130500 $Y=41390
X3988 1 DigitalLDOLogic_VIA1 $T=130750 45700 0 0 $X=130500 $Y=45470
X3989 1 DigitalLDOLogic_VIA1 $T=130750 49780 0 0 $X=130500 $Y=49550
X3990 1 DigitalLDOLogic_VIA1 $T=130750 53860 0 0 $X=130500 $Y=53630
X3991 1 DigitalLDOLogic_VIA1 $T=130750 57940 0 0 $X=130500 $Y=57710
X3992 3 DigitalLDOLogic_VIA1 $T=132590 11700 0 0 $X=132340 $Y=11470
X3993 3 DigitalLDOLogic_VIA1 $T=132590 15780 0 0 $X=132340 $Y=15550
X3994 3 DigitalLDOLogic_VIA1 $T=132590 19860 0 0 $X=132340 $Y=19630
X3995 3 DigitalLDOLogic_VIA1 $T=132590 23940 0 0 $X=132340 $Y=23710
X3996 3 DigitalLDOLogic_VIA1 $T=132590 28020 0 0 $X=132340 $Y=27790
X3997 3 DigitalLDOLogic_VIA1 $T=132590 32100 0 0 $X=132340 $Y=31870
X3998 3 DigitalLDOLogic_VIA1 $T=132590 36180 0 0 $X=132340 $Y=35950
X3999 3 DigitalLDOLogic_VIA1 $T=132590 40260 0 0 $X=132340 $Y=40030
X4000 3 DigitalLDOLogic_VIA1 $T=132590 44340 0 0 $X=132340 $Y=44110
X4001 3 DigitalLDOLogic_VIA1 $T=132590 48420 0 0 $X=132340 $Y=48190
X4002 3 DigitalLDOLogic_VIA1 $T=132590 52500 0 0 $X=132340 $Y=52270
X4003 3 DigitalLDOLogic_VIA1 $T=132590 56580 0 0 $X=132340 $Y=56350
X4004 1 DigitalLDOLogic_VIA1 $T=133510 13060 0 0 $X=133260 $Y=12830
X4005 1 DigitalLDOLogic_VIA1 $T=133510 17140 0 0 $X=133260 $Y=16910
X4006 1 DigitalLDOLogic_VIA1 $T=133510 21220 0 0 $X=133260 $Y=20990
X4007 1 DigitalLDOLogic_VIA1 $T=133510 25300 0 0 $X=133260 $Y=25070
X4008 1 DigitalLDOLogic_VIA1 $T=133510 29380 0 0 $X=133260 $Y=29150
X4009 1 DigitalLDOLogic_VIA1 $T=133510 33460 0 0 $X=133260 $Y=33230
X4010 1 DigitalLDOLogic_VIA1 $T=133510 37540 0 0 $X=133260 $Y=37310
X4011 1 DigitalLDOLogic_VIA1 $T=133510 41620 0 0 $X=133260 $Y=41390
X4012 1 DigitalLDOLogic_VIA1 $T=133510 45700 0 0 $X=133260 $Y=45470
X4013 1 DigitalLDOLogic_VIA1 $T=133510 49780 0 0 $X=133260 $Y=49550
X4014 1 DigitalLDOLogic_VIA1 $T=133510 53860 0 0 $X=133260 $Y=53630
X4015 1 DigitalLDOLogic_VIA1 $T=133510 57940 0 0 $X=133260 $Y=57710
X4016 3 DigitalLDOLogic_VIA1 $T=135350 11700 0 0 $X=135100 $Y=11470
X4017 3 DigitalLDOLogic_VIA1 $T=135350 15780 0 0 $X=135100 $Y=15550
X4018 3 DigitalLDOLogic_VIA1 $T=135350 19860 0 0 $X=135100 $Y=19630
X4019 3 DigitalLDOLogic_VIA1 $T=135350 23940 0 0 $X=135100 $Y=23710
X4020 3 DigitalLDOLogic_VIA1 $T=135350 28020 0 0 $X=135100 $Y=27790
X4021 3 DigitalLDOLogic_VIA1 $T=135350 32100 0 0 $X=135100 $Y=31870
X4022 3 DigitalLDOLogic_VIA1 $T=135350 36180 0 0 $X=135100 $Y=35950
X4023 3 DigitalLDOLogic_VIA1 $T=135350 40260 0 0 $X=135100 $Y=40030
X4024 3 DigitalLDOLogic_VIA1 $T=135350 44340 0 0 $X=135100 $Y=44110
X4025 3 DigitalLDOLogic_VIA1 $T=135350 48420 0 0 $X=135100 $Y=48190
X4026 3 DigitalLDOLogic_VIA1 $T=135350 52500 0 0 $X=135100 $Y=52270
X4027 3 DigitalLDOLogic_VIA1 $T=135350 56580 0 0 $X=135100 $Y=56350
X4028 1 DigitalLDOLogic_VIA1 $T=136270 13060 0 0 $X=136020 $Y=12830
X4029 1 DigitalLDOLogic_VIA1 $T=136270 17140 0 0 $X=136020 $Y=16910
X4030 1 DigitalLDOLogic_VIA1 $T=136270 21220 0 0 $X=136020 $Y=20990
X4031 1 DigitalLDOLogic_VIA1 $T=136270 25300 0 0 $X=136020 $Y=25070
X4032 1 DigitalLDOLogic_VIA1 $T=136270 29380 0 0 $X=136020 $Y=29150
X4033 1 DigitalLDOLogic_VIA1 $T=136270 33460 0 0 $X=136020 $Y=33230
X4034 1 DigitalLDOLogic_VIA1 $T=136270 37540 0 0 $X=136020 $Y=37310
X4035 1 DigitalLDOLogic_VIA1 $T=136270 41620 0 0 $X=136020 $Y=41390
X4036 1 DigitalLDOLogic_VIA1 $T=136270 45700 0 0 $X=136020 $Y=45470
X4037 1 DigitalLDOLogic_VIA1 $T=136270 49780 0 0 $X=136020 $Y=49550
X4038 1 DigitalLDOLogic_VIA1 $T=136270 53860 0 0 $X=136020 $Y=53630
X4039 1 DigitalLDOLogic_VIA1 $T=136270 57940 0 0 $X=136020 $Y=57710
X4040 3 DigitalLDOLogic_VIA1 $T=138110 11700 0 0 $X=137860 $Y=11470
X4041 3 DigitalLDOLogic_VIA1 $T=138110 15780 0 0 $X=137860 $Y=15550
X4042 3 DigitalLDOLogic_VIA1 $T=138110 19860 0 0 $X=137860 $Y=19630
X4043 3 DigitalLDOLogic_VIA1 $T=138110 23940 0 0 $X=137860 $Y=23710
X4044 3 DigitalLDOLogic_VIA1 $T=138110 28020 0 0 $X=137860 $Y=27790
X4045 3 DigitalLDOLogic_VIA1 $T=138110 32100 0 0 $X=137860 $Y=31870
X4046 3 DigitalLDOLogic_VIA1 $T=138110 36180 0 0 $X=137860 $Y=35950
X4047 3 DigitalLDOLogic_VIA1 $T=138110 40260 0 0 $X=137860 $Y=40030
X4048 3 DigitalLDOLogic_VIA1 $T=138110 44340 0 0 $X=137860 $Y=44110
X4049 3 DigitalLDOLogic_VIA1 $T=138110 48420 0 0 $X=137860 $Y=48190
X4050 3 DigitalLDOLogic_VIA1 $T=138110 52500 0 0 $X=137860 $Y=52270
X4051 3 DigitalLDOLogic_VIA1 $T=138110 56580 0 0 $X=137860 $Y=56350
X4052 1 DigitalLDOLogic_VIA1 $T=139030 13060 0 0 $X=138780 $Y=12830
X4053 1 DigitalLDOLogic_VIA1 $T=139030 17140 0 0 $X=138780 $Y=16910
X4054 1 DigitalLDOLogic_VIA1 $T=139030 21220 0 0 $X=138780 $Y=20990
X4055 1 DigitalLDOLogic_VIA1 $T=139030 25300 0 0 $X=138780 $Y=25070
X4056 1 DigitalLDOLogic_VIA1 $T=139030 29380 0 0 $X=138780 $Y=29150
X4057 1 DigitalLDOLogic_VIA1 $T=139030 33460 0 0 $X=138780 $Y=33230
X4058 1 DigitalLDOLogic_VIA1 $T=139030 37540 0 0 $X=138780 $Y=37310
X4059 1 DigitalLDOLogic_VIA1 $T=139030 41620 0 0 $X=138780 $Y=41390
X4060 1 DigitalLDOLogic_VIA1 $T=139030 45700 0 0 $X=138780 $Y=45470
X4061 1 DigitalLDOLogic_VIA1 $T=139030 49780 0 0 $X=138780 $Y=49550
X4062 1 DigitalLDOLogic_VIA1 $T=139030 53860 0 0 $X=138780 $Y=53630
X4063 1 DigitalLDOLogic_VIA1 $T=139030 57940 0 0 $X=138780 $Y=57710
X4064 3 DigitalLDOLogic_VIA1 $T=140870 11700 0 0 $X=140620 $Y=11470
X4065 3 DigitalLDOLogic_VIA1 $T=140870 15780 0 0 $X=140620 $Y=15550
X4066 3 DigitalLDOLogic_VIA1 $T=140870 19860 0 0 $X=140620 $Y=19630
X4067 3 DigitalLDOLogic_VIA1 $T=140870 23940 0 0 $X=140620 $Y=23710
X4068 3 DigitalLDOLogic_VIA1 $T=140870 28020 0 0 $X=140620 $Y=27790
X4069 3 DigitalLDOLogic_VIA1 $T=140870 32100 0 0 $X=140620 $Y=31870
X4070 3 DigitalLDOLogic_VIA1 $T=140870 36180 0 0 $X=140620 $Y=35950
X4071 3 DigitalLDOLogic_VIA1 $T=140870 40260 0 0 $X=140620 $Y=40030
X4072 3 DigitalLDOLogic_VIA1 $T=140870 44340 0 0 $X=140620 $Y=44110
X4073 3 DigitalLDOLogic_VIA1 $T=140870 48420 0 0 $X=140620 $Y=48190
X4074 3 DigitalLDOLogic_VIA1 $T=140870 52500 0 0 $X=140620 $Y=52270
X4075 3 DigitalLDOLogic_VIA1 $T=140870 56580 0 0 $X=140620 $Y=56350
X4076 1 DigitalLDOLogic_VIA1 $T=141790 13060 0 0 $X=141540 $Y=12830
X4077 1 DigitalLDOLogic_VIA1 $T=141790 17140 0 0 $X=141540 $Y=16910
X4078 1 DigitalLDOLogic_VIA1 $T=141790 21220 0 0 $X=141540 $Y=20990
X4079 1 DigitalLDOLogic_VIA1 $T=141790 25300 0 0 $X=141540 $Y=25070
X4080 1 DigitalLDOLogic_VIA1 $T=141790 29380 0 0 $X=141540 $Y=29150
X4081 1 DigitalLDOLogic_VIA1 $T=141790 33460 0 0 $X=141540 $Y=33230
X4082 1 DigitalLDOLogic_VIA1 $T=141790 37540 0 0 $X=141540 $Y=37310
X4083 1 DigitalLDOLogic_VIA1 $T=141790 41620 0 0 $X=141540 $Y=41390
X4084 1 DigitalLDOLogic_VIA1 $T=141790 45700 0 0 $X=141540 $Y=45470
X4085 1 DigitalLDOLogic_VIA1 $T=141790 49780 0 0 $X=141540 $Y=49550
X4086 1 DigitalLDOLogic_VIA1 $T=141790 53860 0 0 $X=141540 $Y=53630
X4087 1 DigitalLDOLogic_VIA1 $T=141790 57940 0 0 $X=141540 $Y=57710
X4088 3 DigitalLDOLogic_VIA1 $T=143630 11700 0 0 $X=143380 $Y=11470
X4089 3 DigitalLDOLogic_VIA1 $T=143630 15780 0 0 $X=143380 $Y=15550
X4090 3 DigitalLDOLogic_VIA1 $T=143630 19860 0 0 $X=143380 $Y=19630
X4091 3 DigitalLDOLogic_VIA1 $T=143630 23940 0 0 $X=143380 $Y=23710
X4092 3 DigitalLDOLogic_VIA1 $T=143630 28020 0 0 $X=143380 $Y=27790
X4093 3 DigitalLDOLogic_VIA1 $T=143630 32100 0 0 $X=143380 $Y=31870
X4094 3 DigitalLDOLogic_VIA1 $T=143630 36180 0 0 $X=143380 $Y=35950
X4095 3 DigitalLDOLogic_VIA1 $T=143630 40260 0 0 $X=143380 $Y=40030
X4096 3 DigitalLDOLogic_VIA1 $T=143630 44340 0 0 $X=143380 $Y=44110
X4097 3 DigitalLDOLogic_VIA1 $T=143630 48420 0 0 $X=143380 $Y=48190
X4098 3 DigitalLDOLogic_VIA1 $T=143630 52500 0 0 $X=143380 $Y=52270
X4099 3 DigitalLDOLogic_VIA1 $T=143630 56580 0 0 $X=143380 $Y=56350
X4100 1 DigitalLDOLogic_VIA1 $T=144550 13060 0 0 $X=144300 $Y=12830
X4101 1 DigitalLDOLogic_VIA1 $T=144550 17140 0 0 $X=144300 $Y=16910
X4102 1 DigitalLDOLogic_VIA1 $T=144550 21220 0 0 $X=144300 $Y=20990
X4103 1 DigitalLDOLogic_VIA1 $T=144550 25300 0 0 $X=144300 $Y=25070
X4104 1 DigitalLDOLogic_VIA1 $T=144550 29380 0 0 $X=144300 $Y=29150
X4105 1 DigitalLDOLogic_VIA1 $T=144550 33460 0 0 $X=144300 $Y=33230
X4106 1 DigitalLDOLogic_VIA1 $T=144550 37540 0 0 $X=144300 $Y=37310
X4107 1 DigitalLDOLogic_VIA1 $T=144550 41620 0 0 $X=144300 $Y=41390
X4108 1 DigitalLDOLogic_VIA1 $T=144550 45700 0 0 $X=144300 $Y=45470
X4109 1 DigitalLDOLogic_VIA1 $T=144550 49780 0 0 $X=144300 $Y=49550
X4110 1 DigitalLDOLogic_VIA1 $T=144550 53860 0 0 $X=144300 $Y=53630
X4111 1 DigitalLDOLogic_VIA1 $T=144550 57940 0 0 $X=144300 $Y=57710
X4112 3 DigitalLDOLogic_VIA1 $T=146390 11700 0 0 $X=146140 $Y=11470
X4113 3 DigitalLDOLogic_VIA1 $T=146390 15780 0 0 $X=146140 $Y=15550
X4114 3 DigitalLDOLogic_VIA1 $T=146390 19860 0 0 $X=146140 $Y=19630
X4115 3 DigitalLDOLogic_VIA1 $T=146390 23940 0 0 $X=146140 $Y=23710
X4116 3 DigitalLDOLogic_VIA1 $T=146390 28020 0 0 $X=146140 $Y=27790
X4117 3 DigitalLDOLogic_VIA1 $T=146390 32100 0 0 $X=146140 $Y=31870
X4118 3 DigitalLDOLogic_VIA1 $T=146390 36180 0 0 $X=146140 $Y=35950
X4119 3 DigitalLDOLogic_VIA1 $T=146390 40260 0 0 $X=146140 $Y=40030
X4120 3 DigitalLDOLogic_VIA1 $T=146390 44340 0 0 $X=146140 $Y=44110
X4121 3 DigitalLDOLogic_VIA1 $T=146390 48420 0 0 $X=146140 $Y=48190
X4122 3 DigitalLDOLogic_VIA1 $T=146390 52500 0 0 $X=146140 $Y=52270
X4123 3 DigitalLDOLogic_VIA1 $T=146390 56580 0 0 $X=146140 $Y=56350
X4124 1 DigitalLDOLogic_VIA1 $T=147310 13060 0 0 $X=147060 $Y=12830
X4125 1 DigitalLDOLogic_VIA1 $T=147310 17140 0 0 $X=147060 $Y=16910
X4126 1 DigitalLDOLogic_VIA1 $T=147310 21220 0 0 $X=147060 $Y=20990
X4127 1 DigitalLDOLogic_VIA1 $T=147310 25300 0 0 $X=147060 $Y=25070
X4128 1 DigitalLDOLogic_VIA1 $T=147310 29380 0 0 $X=147060 $Y=29150
X4129 1 DigitalLDOLogic_VIA1 $T=147310 33460 0 0 $X=147060 $Y=33230
X4130 1 DigitalLDOLogic_VIA1 $T=147310 37540 0 0 $X=147060 $Y=37310
X4131 1 DigitalLDOLogic_VIA1 $T=147310 41620 0 0 $X=147060 $Y=41390
X4132 1 DigitalLDOLogic_VIA1 $T=147310 45700 0 0 $X=147060 $Y=45470
X4133 1 DigitalLDOLogic_VIA1 $T=147310 49780 0 0 $X=147060 $Y=49550
X4134 1 DigitalLDOLogic_VIA1 $T=147310 53860 0 0 $X=147060 $Y=53630
X4135 1 DigitalLDOLogic_VIA1 $T=147310 57940 0 0 $X=147060 $Y=57710
X4136 3 DigitalLDOLogic_VIA1 $T=149150 11700 0 0 $X=148900 $Y=11470
X4137 3 DigitalLDOLogic_VIA1 $T=149150 15780 0 0 $X=148900 $Y=15550
X4138 3 DigitalLDOLogic_VIA1 $T=149150 19860 0 0 $X=148900 $Y=19630
X4139 3 DigitalLDOLogic_VIA1 $T=149150 23940 0 0 $X=148900 $Y=23710
X4140 3 DigitalLDOLogic_VIA1 $T=149150 28020 0 0 $X=148900 $Y=27790
X4141 3 DigitalLDOLogic_VIA1 $T=149150 32100 0 0 $X=148900 $Y=31870
X4142 3 DigitalLDOLogic_VIA1 $T=149150 36180 0 0 $X=148900 $Y=35950
X4143 3 DigitalLDOLogic_VIA1 $T=149150 40260 0 0 $X=148900 $Y=40030
X4144 3 DigitalLDOLogic_VIA1 $T=149150 44340 0 0 $X=148900 $Y=44110
X4145 3 DigitalLDOLogic_VIA1 $T=149150 48420 0 0 $X=148900 $Y=48190
X4146 3 DigitalLDOLogic_VIA1 $T=149150 52500 0 0 $X=148900 $Y=52270
X4147 3 DigitalLDOLogic_VIA1 $T=149150 56580 0 0 $X=148900 $Y=56350
X4148 1 DigitalLDOLogic_VIA1 $T=150070 13060 0 0 $X=149820 $Y=12830
X4149 1 DigitalLDOLogic_VIA1 $T=150070 17140 0 0 $X=149820 $Y=16910
X4150 1 DigitalLDOLogic_VIA1 $T=150070 21220 0 0 $X=149820 $Y=20990
X4151 1 DigitalLDOLogic_VIA1 $T=150070 25300 0 0 $X=149820 $Y=25070
X4152 1 DigitalLDOLogic_VIA1 $T=150070 29380 0 0 $X=149820 $Y=29150
X4153 1 DigitalLDOLogic_VIA1 $T=150070 33460 0 0 $X=149820 $Y=33230
X4154 1 DigitalLDOLogic_VIA1 $T=150070 37540 0 0 $X=149820 $Y=37310
X4155 1 DigitalLDOLogic_VIA1 $T=150070 41620 0 0 $X=149820 $Y=41390
X4156 1 DigitalLDOLogic_VIA1 $T=150070 45700 0 0 $X=149820 $Y=45470
X4157 1 DigitalLDOLogic_VIA1 $T=150070 49780 0 0 $X=149820 $Y=49550
X4158 1 DigitalLDOLogic_VIA1 $T=150070 53860 0 0 $X=149820 $Y=53630
X4159 1 DigitalLDOLogic_VIA1 $T=150070 57940 0 0 $X=149820 $Y=57710
X4160 3 DigitalLDOLogic_VIA1 $T=151910 11700 0 0 $X=151660 $Y=11470
X4161 3 DigitalLDOLogic_VIA1 $T=151910 15780 0 0 $X=151660 $Y=15550
X4162 3 DigitalLDOLogic_VIA1 $T=151910 19860 0 0 $X=151660 $Y=19630
X4163 3 DigitalLDOLogic_VIA1 $T=151910 23940 0 0 $X=151660 $Y=23710
X4164 3 DigitalLDOLogic_VIA1 $T=151910 28020 0 0 $X=151660 $Y=27790
X4165 3 DigitalLDOLogic_VIA1 $T=151910 32100 0 0 $X=151660 $Y=31870
X4166 3 DigitalLDOLogic_VIA1 $T=151910 36180 0 0 $X=151660 $Y=35950
X4167 3 DigitalLDOLogic_VIA1 $T=151910 40260 0 0 $X=151660 $Y=40030
X4168 3 DigitalLDOLogic_VIA1 $T=151910 44340 0 0 $X=151660 $Y=44110
X4169 3 DigitalLDOLogic_VIA1 $T=151910 48420 0 0 $X=151660 $Y=48190
X4170 3 DigitalLDOLogic_VIA1 $T=151910 52500 0 0 $X=151660 $Y=52270
X4171 3 DigitalLDOLogic_VIA1 $T=151910 56580 0 0 $X=151660 $Y=56350
X4172 1 DigitalLDOLogic_VIA1 $T=152830 13060 0 0 $X=152580 $Y=12830
X4173 1 DigitalLDOLogic_VIA1 $T=152830 17140 0 0 $X=152580 $Y=16910
X4174 1 DigitalLDOLogic_VIA1 $T=152830 21220 0 0 $X=152580 $Y=20990
X4175 1 DigitalLDOLogic_VIA1 $T=152830 25300 0 0 $X=152580 $Y=25070
X4176 1 DigitalLDOLogic_VIA1 $T=152830 29380 0 0 $X=152580 $Y=29150
X4177 1 DigitalLDOLogic_VIA1 $T=152830 33460 0 0 $X=152580 $Y=33230
X4178 1 DigitalLDOLogic_VIA1 $T=152830 37540 0 0 $X=152580 $Y=37310
X4179 1 DigitalLDOLogic_VIA1 $T=152830 41620 0 0 $X=152580 $Y=41390
X4180 1 DigitalLDOLogic_VIA1 $T=152830 45700 0 0 $X=152580 $Y=45470
X4181 1 DigitalLDOLogic_VIA1 $T=152830 49780 0 0 $X=152580 $Y=49550
X4182 1 DigitalLDOLogic_VIA1 $T=152830 53860 0 0 $X=152580 $Y=53630
X4183 1 DigitalLDOLogic_VIA1 $T=152830 57940 0 0 $X=152580 $Y=57710
X4184 3 DigitalLDOLogic_VIA1 $T=154670 11700 0 0 $X=154420 $Y=11470
X4185 3 DigitalLDOLogic_VIA1 $T=154670 15780 0 0 $X=154420 $Y=15550
X4186 3 DigitalLDOLogic_VIA1 $T=154670 19860 0 0 $X=154420 $Y=19630
X4187 3 DigitalLDOLogic_VIA1 $T=154670 23940 0 0 $X=154420 $Y=23710
X4188 3 DigitalLDOLogic_VIA1 $T=154670 28020 0 0 $X=154420 $Y=27790
X4189 3 DigitalLDOLogic_VIA1 $T=154670 32100 0 0 $X=154420 $Y=31870
X4190 3 DigitalLDOLogic_VIA1 $T=154670 36180 0 0 $X=154420 $Y=35950
X4191 3 DigitalLDOLogic_VIA1 $T=154670 40260 0 0 $X=154420 $Y=40030
X4192 3 DigitalLDOLogic_VIA1 $T=154670 44340 0 0 $X=154420 $Y=44110
X4193 3 DigitalLDOLogic_VIA1 $T=154670 48420 0 0 $X=154420 $Y=48190
X4194 3 DigitalLDOLogic_VIA1 $T=154670 52500 0 0 $X=154420 $Y=52270
X4195 3 DigitalLDOLogic_VIA1 $T=154670 56580 0 0 $X=154420 $Y=56350
X4196 1 DigitalLDOLogic_VIA1 $T=155590 13060 0 0 $X=155340 $Y=12830
X4197 1 DigitalLDOLogic_VIA1 $T=155590 17140 0 0 $X=155340 $Y=16910
X4198 1 DigitalLDOLogic_VIA1 $T=155590 21220 0 0 $X=155340 $Y=20990
X4199 1 DigitalLDOLogic_VIA1 $T=155590 25300 0 0 $X=155340 $Y=25070
X4200 1 DigitalLDOLogic_VIA1 $T=155590 29380 0 0 $X=155340 $Y=29150
X4201 1 DigitalLDOLogic_VIA1 $T=155590 33460 0 0 $X=155340 $Y=33230
X4202 1 DigitalLDOLogic_VIA1 $T=155590 37540 0 0 $X=155340 $Y=37310
X4203 1 DigitalLDOLogic_VIA1 $T=155590 41620 0 0 $X=155340 $Y=41390
X4204 1 DigitalLDOLogic_VIA1 $T=155590 45700 0 0 $X=155340 $Y=45470
X4205 1 DigitalLDOLogic_VIA1 $T=155590 49780 0 0 $X=155340 $Y=49550
X4206 1 DigitalLDOLogic_VIA1 $T=155590 53860 0 0 $X=155340 $Y=53630
X4207 1 DigitalLDOLogic_VIA1 $T=155590 57940 0 0 $X=155340 $Y=57710
X4208 3 DigitalLDOLogic_VIA1 $T=157430 11700 0 0 $X=157180 $Y=11470
X4209 3 DigitalLDOLogic_VIA1 $T=157430 15780 0 0 $X=157180 $Y=15550
X4210 3 DigitalLDOLogic_VIA1 $T=157430 19860 0 0 $X=157180 $Y=19630
X4211 3 DigitalLDOLogic_VIA1 $T=157430 23940 0 0 $X=157180 $Y=23710
X4212 3 DigitalLDOLogic_VIA1 $T=157430 28020 0 0 $X=157180 $Y=27790
X4213 3 DigitalLDOLogic_VIA1 $T=157430 32100 0 0 $X=157180 $Y=31870
X4214 3 DigitalLDOLogic_VIA1 $T=157430 36180 0 0 $X=157180 $Y=35950
X4215 3 DigitalLDOLogic_VIA1 $T=157430 40260 0 0 $X=157180 $Y=40030
X4216 3 DigitalLDOLogic_VIA1 $T=157430 44340 0 0 $X=157180 $Y=44110
X4217 3 DigitalLDOLogic_VIA1 $T=157430 48420 0 0 $X=157180 $Y=48190
X4218 3 DigitalLDOLogic_VIA1 $T=157430 52500 0 0 $X=157180 $Y=52270
X4219 3 DigitalLDOLogic_VIA1 $T=157430 56580 0 0 $X=157180 $Y=56350
X4220 1 DigitalLDOLogic_VIA1 $T=158350 13060 0 0 $X=158100 $Y=12830
X4221 1 DigitalLDOLogic_VIA1 $T=158350 17140 0 0 $X=158100 $Y=16910
X4222 1 DigitalLDOLogic_VIA1 $T=158350 21220 0 0 $X=158100 $Y=20990
X4223 1 DigitalLDOLogic_VIA1 $T=158350 25300 0 0 $X=158100 $Y=25070
X4224 1 DigitalLDOLogic_VIA1 $T=158350 29380 0 0 $X=158100 $Y=29150
X4225 1 DigitalLDOLogic_VIA1 $T=158350 33460 0 0 $X=158100 $Y=33230
X4226 1 DigitalLDOLogic_VIA1 $T=158350 37540 0 0 $X=158100 $Y=37310
X4227 1 DigitalLDOLogic_VIA1 $T=158350 41620 0 0 $X=158100 $Y=41390
X4228 1 DigitalLDOLogic_VIA1 $T=158350 45700 0 0 $X=158100 $Y=45470
X4229 1 DigitalLDOLogic_VIA1 $T=158350 49780 0 0 $X=158100 $Y=49550
X4230 1 DigitalLDOLogic_VIA1 $T=158350 53860 0 0 $X=158100 $Y=53630
X4231 1 DigitalLDOLogic_VIA1 $T=158350 57940 0 0 $X=158100 $Y=57710
X4232 3 DigitalLDOLogic_VIA1 $T=160190 11700 0 0 $X=159940 $Y=11470
X4233 3 DigitalLDOLogic_VIA1 $T=160190 15780 0 0 $X=159940 $Y=15550
X4234 3 DigitalLDOLogic_VIA1 $T=160190 19860 0 0 $X=159940 $Y=19630
X4235 3 DigitalLDOLogic_VIA1 $T=160190 23940 0 0 $X=159940 $Y=23710
X4236 3 DigitalLDOLogic_VIA1 $T=160190 28020 0 0 $X=159940 $Y=27790
X4237 3 DigitalLDOLogic_VIA1 $T=160190 32100 0 0 $X=159940 $Y=31870
X4238 3 DigitalLDOLogic_VIA1 $T=160190 36180 0 0 $X=159940 $Y=35950
X4239 3 DigitalLDOLogic_VIA1 $T=160190 40260 0 0 $X=159940 $Y=40030
X4240 3 DigitalLDOLogic_VIA1 $T=160190 44340 0 0 $X=159940 $Y=44110
X4241 3 DigitalLDOLogic_VIA1 $T=160190 48420 0 0 $X=159940 $Y=48190
X4242 3 DigitalLDOLogic_VIA1 $T=160190 52500 0 0 $X=159940 $Y=52270
X4243 3 DigitalLDOLogic_VIA1 $T=160190 56580 0 0 $X=159940 $Y=56350
X4244 1 DigitalLDOLogic_VIA1 $T=161110 13060 0 0 $X=160860 $Y=12830
X4245 1 DigitalLDOLogic_VIA1 $T=161110 17140 0 0 $X=160860 $Y=16910
X4246 1 DigitalLDOLogic_VIA1 $T=161110 21220 0 0 $X=160860 $Y=20990
X4247 1 DigitalLDOLogic_VIA1 $T=161110 25300 0 0 $X=160860 $Y=25070
X4248 1 DigitalLDOLogic_VIA1 $T=161110 29380 0 0 $X=160860 $Y=29150
X4249 1 DigitalLDOLogic_VIA1 $T=161110 33460 0 0 $X=160860 $Y=33230
X4250 1 DigitalLDOLogic_VIA1 $T=161110 37540 0 0 $X=160860 $Y=37310
X4251 1 DigitalLDOLogic_VIA1 $T=161110 41620 0 0 $X=160860 $Y=41390
X4252 1 DigitalLDOLogic_VIA1 $T=161110 45700 0 0 $X=160860 $Y=45470
X4253 1 DigitalLDOLogic_VIA1 $T=161110 49780 0 0 $X=160860 $Y=49550
X4254 1 DigitalLDOLogic_VIA1 $T=161110 53860 0 0 $X=160860 $Y=53630
X4255 1 DigitalLDOLogic_VIA1 $T=161110 57940 0 0 $X=160860 $Y=57710
X4256 3 DigitalLDOLogic_VIA1 $T=162950 11700 0 0 $X=162700 $Y=11470
X4257 3 DigitalLDOLogic_VIA1 $T=162950 15780 0 0 $X=162700 $Y=15550
X4258 3 DigitalLDOLogic_VIA1 $T=162950 19860 0 0 $X=162700 $Y=19630
X4259 3 DigitalLDOLogic_VIA1 $T=162950 23940 0 0 $X=162700 $Y=23710
X4260 3 DigitalLDOLogic_VIA1 $T=162950 28020 0 0 $X=162700 $Y=27790
X4261 3 DigitalLDOLogic_VIA1 $T=162950 32100 0 0 $X=162700 $Y=31870
X4262 3 DigitalLDOLogic_VIA1 $T=162950 36180 0 0 $X=162700 $Y=35950
X4263 3 DigitalLDOLogic_VIA1 $T=162950 40260 0 0 $X=162700 $Y=40030
X4264 3 DigitalLDOLogic_VIA1 $T=162950 44340 0 0 $X=162700 $Y=44110
X4265 3 DigitalLDOLogic_VIA1 $T=162950 48420 0 0 $X=162700 $Y=48190
X4266 3 DigitalLDOLogic_VIA1 $T=162950 52500 0 0 $X=162700 $Y=52270
X4267 3 DigitalLDOLogic_VIA1 $T=162950 56580 0 0 $X=162700 $Y=56350
X4268 1 DigitalLDOLogic_VIA1 $T=163870 13060 0 0 $X=163620 $Y=12830
X4269 1 DigitalLDOLogic_VIA1 $T=163870 17140 0 0 $X=163620 $Y=16910
X4270 1 DigitalLDOLogic_VIA1 $T=163870 21220 0 0 $X=163620 $Y=20990
X4271 1 DigitalLDOLogic_VIA1 $T=163870 25300 0 0 $X=163620 $Y=25070
X4272 1 DigitalLDOLogic_VIA1 $T=163870 29380 0 0 $X=163620 $Y=29150
X4273 1 DigitalLDOLogic_VIA1 $T=163870 33460 0 0 $X=163620 $Y=33230
X4274 1 DigitalLDOLogic_VIA1 $T=163870 37540 0 0 $X=163620 $Y=37310
X4275 1 DigitalLDOLogic_VIA1 $T=163870 41620 0 0 $X=163620 $Y=41390
X4276 1 DigitalLDOLogic_VIA1 $T=163870 45700 0 0 $X=163620 $Y=45470
X4277 1 DigitalLDOLogic_VIA1 $T=163870 49780 0 0 $X=163620 $Y=49550
X4278 1 DigitalLDOLogic_VIA1 $T=163870 53860 0 0 $X=163620 $Y=53630
X4279 1 DigitalLDOLogic_VIA1 $T=163870 57940 0 0 $X=163620 $Y=57710
X4280 3 DigitalLDOLogic_VIA1 $T=165710 11700 0 0 $X=165460 $Y=11470
X4281 3 DigitalLDOLogic_VIA1 $T=165710 15780 0 0 $X=165460 $Y=15550
X4282 3 DigitalLDOLogic_VIA1 $T=165710 19860 0 0 $X=165460 $Y=19630
X4283 3 DigitalLDOLogic_VIA1 $T=165710 23940 0 0 $X=165460 $Y=23710
X4284 3 DigitalLDOLogic_VIA1 $T=165710 28020 0 0 $X=165460 $Y=27790
X4285 3 DigitalLDOLogic_VIA1 $T=165710 32100 0 0 $X=165460 $Y=31870
X4286 3 DigitalLDOLogic_VIA1 $T=165710 36180 0 0 $X=165460 $Y=35950
X4287 3 DigitalLDOLogic_VIA1 $T=165710 40260 0 0 $X=165460 $Y=40030
X4288 3 DigitalLDOLogic_VIA1 $T=165710 44340 0 0 $X=165460 $Y=44110
X4289 3 DigitalLDOLogic_VIA1 $T=165710 48420 0 0 $X=165460 $Y=48190
X4290 3 DigitalLDOLogic_VIA1 $T=165710 52500 0 0 $X=165460 $Y=52270
X4291 3 DigitalLDOLogic_VIA1 $T=165710 56580 0 0 $X=165460 $Y=56350
X4292 1 DigitalLDOLogic_VIA1 $T=166630 13060 0 0 $X=166380 $Y=12830
X4293 1 DigitalLDOLogic_VIA1 $T=166630 17140 0 0 $X=166380 $Y=16910
X4294 1 DigitalLDOLogic_VIA1 $T=166630 21220 0 0 $X=166380 $Y=20990
X4295 1 DigitalLDOLogic_VIA1 $T=166630 25300 0 0 $X=166380 $Y=25070
X4296 1 DigitalLDOLogic_VIA1 $T=166630 29380 0 0 $X=166380 $Y=29150
X4297 1 DigitalLDOLogic_VIA1 $T=166630 33460 0 0 $X=166380 $Y=33230
X4298 1 DigitalLDOLogic_VIA1 $T=166630 37540 0 0 $X=166380 $Y=37310
X4299 1 DigitalLDOLogic_VIA1 $T=166630 41620 0 0 $X=166380 $Y=41390
X4300 1 DigitalLDOLogic_VIA1 $T=166630 45700 0 0 $X=166380 $Y=45470
X4301 1 DigitalLDOLogic_VIA1 $T=166630 49780 0 0 $X=166380 $Y=49550
X4302 1 DigitalLDOLogic_VIA1 $T=166630 53860 0 0 $X=166380 $Y=53630
X4303 1 DigitalLDOLogic_VIA1 $T=166630 57940 0 0 $X=166380 $Y=57710
X4304 3 DigitalLDOLogic_VIA1 $T=168470 11700 0 0 $X=168220 $Y=11470
X4305 3 DigitalLDOLogic_VIA1 $T=168470 15780 0 0 $X=168220 $Y=15550
X4306 3 DigitalLDOLogic_VIA1 $T=168470 19860 0 0 $X=168220 $Y=19630
X4307 3 DigitalLDOLogic_VIA1 $T=168470 23940 0 0 $X=168220 $Y=23710
X4308 3 DigitalLDOLogic_VIA1 $T=168470 28020 0 0 $X=168220 $Y=27790
X4309 3 DigitalLDOLogic_VIA1 $T=168470 32100 0 0 $X=168220 $Y=31870
X4310 3 DigitalLDOLogic_VIA1 $T=168470 36180 0 0 $X=168220 $Y=35950
X4311 3 DigitalLDOLogic_VIA1 $T=168470 40260 0 0 $X=168220 $Y=40030
X4312 3 DigitalLDOLogic_VIA1 $T=168470 44340 0 0 $X=168220 $Y=44110
X4313 3 DigitalLDOLogic_VIA1 $T=168470 48420 0 0 $X=168220 $Y=48190
X4314 3 DigitalLDOLogic_VIA1 $T=168470 52500 0 0 $X=168220 $Y=52270
X4315 3 DigitalLDOLogic_VIA1 $T=168470 56580 0 0 $X=168220 $Y=56350
X4316 1 DigitalLDOLogic_VIA1 $T=169390 13060 0 0 $X=169140 $Y=12830
X4317 1 DigitalLDOLogic_VIA1 $T=169390 17140 0 0 $X=169140 $Y=16910
X4318 1 DigitalLDOLogic_VIA1 $T=169390 21220 0 0 $X=169140 $Y=20990
X4319 1 DigitalLDOLogic_VIA1 $T=169390 25300 0 0 $X=169140 $Y=25070
X4320 1 DigitalLDOLogic_VIA1 $T=169390 29380 0 0 $X=169140 $Y=29150
X4321 1 DigitalLDOLogic_VIA1 $T=169390 33460 0 0 $X=169140 $Y=33230
X4322 1 DigitalLDOLogic_VIA1 $T=169390 37540 0 0 $X=169140 $Y=37310
X4323 1 DigitalLDOLogic_VIA1 $T=169390 41620 0 0 $X=169140 $Y=41390
X4324 1 DigitalLDOLogic_VIA1 $T=169390 45700 0 0 $X=169140 $Y=45470
X4325 1 DigitalLDOLogic_VIA1 $T=169390 49780 0 0 $X=169140 $Y=49550
X4326 1 DigitalLDOLogic_VIA1 $T=169390 53860 0 0 $X=169140 $Y=53630
X4327 1 DigitalLDOLogic_VIA1 $T=169390 57940 0 0 $X=169140 $Y=57710
X4328 3 DigitalLDOLogic_VIA1 $T=171230 11700 0 0 $X=170980 $Y=11470
X4329 3 DigitalLDOLogic_VIA1 $T=171230 15780 0 0 $X=170980 $Y=15550
X4330 3 DigitalLDOLogic_VIA1 $T=171230 19860 0 0 $X=170980 $Y=19630
X4331 3 DigitalLDOLogic_VIA1 $T=171230 23940 0 0 $X=170980 $Y=23710
X4332 3 DigitalLDOLogic_VIA1 $T=171230 28020 0 0 $X=170980 $Y=27790
X4333 3 DigitalLDOLogic_VIA1 $T=171230 32100 0 0 $X=170980 $Y=31870
X4334 3 DigitalLDOLogic_VIA1 $T=171230 36180 0 0 $X=170980 $Y=35950
X4335 3 DigitalLDOLogic_VIA1 $T=171230 40260 0 0 $X=170980 $Y=40030
X4336 3 DigitalLDOLogic_VIA1 $T=171230 44340 0 0 $X=170980 $Y=44110
X4337 3 DigitalLDOLogic_VIA1 $T=171230 48420 0 0 $X=170980 $Y=48190
X4338 3 DigitalLDOLogic_VIA1 $T=171230 52500 0 0 $X=170980 $Y=52270
X4339 3 DigitalLDOLogic_VIA1 $T=171230 56580 0 0 $X=170980 $Y=56350
X4340 1 DigitalLDOLogic_VIA1 $T=172150 13060 0 0 $X=171900 $Y=12830
X4341 1 DigitalLDOLogic_VIA1 $T=172150 17140 0 0 $X=171900 $Y=16910
X4342 1 DigitalLDOLogic_VIA1 $T=172150 21220 0 0 $X=171900 $Y=20990
X4343 1 DigitalLDOLogic_VIA1 $T=172150 25300 0 0 $X=171900 $Y=25070
X4344 1 DigitalLDOLogic_VIA1 $T=172150 29380 0 0 $X=171900 $Y=29150
X4345 1 DigitalLDOLogic_VIA1 $T=172150 33460 0 0 $X=171900 $Y=33230
X4346 1 DigitalLDOLogic_VIA1 $T=172150 37540 0 0 $X=171900 $Y=37310
X4347 1 DigitalLDOLogic_VIA1 $T=172150 41620 0 0 $X=171900 $Y=41390
X4348 1 DigitalLDOLogic_VIA1 $T=172150 45700 0 0 $X=171900 $Y=45470
X4349 1 DigitalLDOLogic_VIA1 $T=172150 49780 0 0 $X=171900 $Y=49550
X4350 1 DigitalLDOLogic_VIA1 $T=172150 53860 0 0 $X=171900 $Y=53630
X4351 1 DigitalLDOLogic_VIA1 $T=172150 57940 0 0 $X=171900 $Y=57710
X4352 3 DigitalLDOLogic_VIA1 $T=173990 11700 0 0 $X=173740 $Y=11470
X4353 3 DigitalLDOLogic_VIA1 $T=173990 15780 0 0 $X=173740 $Y=15550
X4354 3 DigitalLDOLogic_VIA1 $T=173990 19860 0 0 $X=173740 $Y=19630
X4355 3 DigitalLDOLogic_VIA1 $T=173990 23940 0 0 $X=173740 $Y=23710
X4356 3 DigitalLDOLogic_VIA1 $T=173990 28020 0 0 $X=173740 $Y=27790
X4357 3 DigitalLDOLogic_VIA1 $T=173990 32100 0 0 $X=173740 $Y=31870
X4358 3 DigitalLDOLogic_VIA1 $T=173990 36180 0 0 $X=173740 $Y=35950
X4359 3 DigitalLDOLogic_VIA1 $T=173990 40260 0 0 $X=173740 $Y=40030
X4360 3 DigitalLDOLogic_VIA1 $T=173990 44340 0 0 $X=173740 $Y=44110
X4361 3 DigitalLDOLogic_VIA1 $T=173990 48420 0 0 $X=173740 $Y=48190
X4362 3 DigitalLDOLogic_VIA1 $T=173990 52500 0 0 $X=173740 $Y=52270
X4363 3 DigitalLDOLogic_VIA1 $T=173990 56580 0 0 $X=173740 $Y=56350
X4364 1 DigitalLDOLogic_VIA1 $T=174910 13060 0 0 $X=174660 $Y=12830
X4365 1 DigitalLDOLogic_VIA1 $T=174910 17140 0 0 $X=174660 $Y=16910
X4366 1 DigitalLDOLogic_VIA1 $T=174910 21220 0 0 $X=174660 $Y=20990
X4367 1 DigitalLDOLogic_VIA1 $T=174910 25300 0 0 $X=174660 $Y=25070
X4368 1 DigitalLDOLogic_VIA1 $T=174910 29380 0 0 $X=174660 $Y=29150
X4369 1 DigitalLDOLogic_VIA1 $T=174910 33460 0 0 $X=174660 $Y=33230
X4370 1 DigitalLDOLogic_VIA1 $T=174910 37540 0 0 $X=174660 $Y=37310
X4371 1 DigitalLDOLogic_VIA1 $T=174910 41620 0 0 $X=174660 $Y=41390
X4372 1 DigitalLDOLogic_VIA1 $T=174910 45700 0 0 $X=174660 $Y=45470
X4373 1 DigitalLDOLogic_VIA1 $T=174910 49780 0 0 $X=174660 $Y=49550
X4374 1 DigitalLDOLogic_VIA1 $T=174910 53860 0 0 $X=174660 $Y=53630
X4375 1 DigitalLDOLogic_VIA1 $T=174910 57940 0 0 $X=174660 $Y=57710
X4376 3 DigitalLDOLogic_VIA1 $T=176750 11700 0 0 $X=176500 $Y=11470
X4377 3 DigitalLDOLogic_VIA1 $T=176750 15780 0 0 $X=176500 $Y=15550
X4378 3 DigitalLDOLogic_VIA1 $T=176750 19860 0 0 $X=176500 $Y=19630
X4379 3 DigitalLDOLogic_VIA1 $T=176750 23940 0 0 $X=176500 $Y=23710
X4380 3 DigitalLDOLogic_VIA1 $T=176750 28020 0 0 $X=176500 $Y=27790
X4381 3 DigitalLDOLogic_VIA1 $T=176750 32100 0 0 $X=176500 $Y=31870
X4382 3 DigitalLDOLogic_VIA1 $T=176750 36180 0 0 $X=176500 $Y=35950
X4383 3 DigitalLDOLogic_VIA1 $T=176750 40260 0 0 $X=176500 $Y=40030
X4384 3 DigitalLDOLogic_VIA1 $T=176750 44340 0 0 $X=176500 $Y=44110
X4385 3 DigitalLDOLogic_VIA1 $T=176750 48420 0 0 $X=176500 $Y=48190
X4386 3 DigitalLDOLogic_VIA1 $T=176750 52500 0 0 $X=176500 $Y=52270
X4387 3 DigitalLDOLogic_VIA1 $T=176750 56580 0 0 $X=176500 $Y=56350
X4388 1 DigitalLDOLogic_VIA1 $T=177670 13060 0 0 $X=177420 $Y=12830
X4389 1 DigitalLDOLogic_VIA1 $T=177670 17140 0 0 $X=177420 $Y=16910
X4390 1 DigitalLDOLogic_VIA1 $T=177670 21220 0 0 $X=177420 $Y=20990
X4391 1 DigitalLDOLogic_VIA1 $T=177670 25300 0 0 $X=177420 $Y=25070
X4392 1 DigitalLDOLogic_VIA1 $T=177670 29380 0 0 $X=177420 $Y=29150
X4393 1 DigitalLDOLogic_VIA1 $T=177670 33460 0 0 $X=177420 $Y=33230
X4394 1 DigitalLDOLogic_VIA1 $T=177670 37540 0 0 $X=177420 $Y=37310
X4395 1 DigitalLDOLogic_VIA1 $T=177670 41620 0 0 $X=177420 $Y=41390
X4396 1 DigitalLDOLogic_VIA1 $T=177670 45700 0 0 $X=177420 $Y=45470
X4397 1 DigitalLDOLogic_VIA1 $T=177670 49780 0 0 $X=177420 $Y=49550
X4398 1 DigitalLDOLogic_VIA1 $T=177670 53860 0 0 $X=177420 $Y=53630
X4399 1 DigitalLDOLogic_VIA1 $T=177670 57940 0 0 $X=177420 $Y=57710
X4400 3 DigitalLDOLogic_VIA1 $T=179510 11700 0 0 $X=179260 $Y=11470
X4401 3 DigitalLDOLogic_VIA1 $T=179510 15780 0 0 $X=179260 $Y=15550
X4402 3 DigitalLDOLogic_VIA1 $T=179510 19860 0 0 $X=179260 $Y=19630
X4403 3 DigitalLDOLogic_VIA1 $T=179510 23940 0 0 $X=179260 $Y=23710
X4404 3 DigitalLDOLogic_VIA1 $T=179510 28020 0 0 $X=179260 $Y=27790
X4405 3 DigitalLDOLogic_VIA1 $T=179510 32100 0 0 $X=179260 $Y=31870
X4406 3 DigitalLDOLogic_VIA1 $T=179510 36180 0 0 $X=179260 $Y=35950
X4407 3 DigitalLDOLogic_VIA1 $T=179510 40260 0 0 $X=179260 $Y=40030
X4408 3 DigitalLDOLogic_VIA1 $T=179510 44340 0 0 $X=179260 $Y=44110
X4409 3 DigitalLDOLogic_VIA1 $T=179510 48420 0 0 $X=179260 $Y=48190
X4410 3 DigitalLDOLogic_VIA1 $T=179510 52500 0 0 $X=179260 $Y=52270
X4411 3 DigitalLDOLogic_VIA1 $T=179510 56580 0 0 $X=179260 $Y=56350
X4412 1 DigitalLDOLogic_VIA1 $T=180430 13060 0 0 $X=180180 $Y=12830
X4413 1 DigitalLDOLogic_VIA1 $T=180430 17140 0 0 $X=180180 $Y=16910
X4414 1 DigitalLDOLogic_VIA1 $T=180430 21220 0 0 $X=180180 $Y=20990
X4415 1 DigitalLDOLogic_VIA1 $T=180430 25300 0 0 $X=180180 $Y=25070
X4416 1 DigitalLDOLogic_VIA1 $T=180430 29380 0 0 $X=180180 $Y=29150
X4417 1 DigitalLDOLogic_VIA1 $T=180430 33460 0 0 $X=180180 $Y=33230
X4418 1 DigitalLDOLogic_VIA1 $T=180430 37540 0 0 $X=180180 $Y=37310
X4419 1 DigitalLDOLogic_VIA1 $T=180430 41620 0 0 $X=180180 $Y=41390
X4420 1 DigitalLDOLogic_VIA1 $T=180430 45700 0 0 $X=180180 $Y=45470
X4421 1 DigitalLDOLogic_VIA1 $T=180430 49780 0 0 $X=180180 $Y=49550
X4422 1 DigitalLDOLogic_VIA1 $T=180430 53860 0 0 $X=180180 $Y=53630
X4423 1 DigitalLDOLogic_VIA1 $T=180430 57940 0 0 $X=180180 $Y=57710
X4424 3 DigitalLDOLogic_VIA1 $T=182270 11700 0 0 $X=182020 $Y=11470
X4425 3 DigitalLDOLogic_VIA1 $T=182270 15780 0 0 $X=182020 $Y=15550
X4426 3 DigitalLDOLogic_VIA1 $T=182270 19860 0 0 $X=182020 $Y=19630
X4427 3 DigitalLDOLogic_VIA1 $T=182270 23940 0 0 $X=182020 $Y=23710
X4428 3 DigitalLDOLogic_VIA1 $T=182270 28020 0 0 $X=182020 $Y=27790
X4429 3 DigitalLDOLogic_VIA1 $T=182270 32100 0 0 $X=182020 $Y=31870
X4430 3 DigitalLDOLogic_VIA1 $T=182270 36180 0 0 $X=182020 $Y=35950
X4431 3 DigitalLDOLogic_VIA1 $T=182270 40260 0 0 $X=182020 $Y=40030
X4432 3 DigitalLDOLogic_VIA1 $T=182270 44340 0 0 $X=182020 $Y=44110
X4433 3 DigitalLDOLogic_VIA1 $T=182270 48420 0 0 $X=182020 $Y=48190
X4434 3 DigitalLDOLogic_VIA1 $T=182270 52500 0 0 $X=182020 $Y=52270
X4435 3 DigitalLDOLogic_VIA1 $T=182270 56580 0 0 $X=182020 $Y=56350
X4436 1 DigitalLDOLogic_VIA1 $T=183190 13060 0 0 $X=182940 $Y=12830
X4437 1 DigitalLDOLogic_VIA1 $T=183190 17140 0 0 $X=182940 $Y=16910
X4438 1 DigitalLDOLogic_VIA1 $T=183190 21220 0 0 $X=182940 $Y=20990
X4439 1 DigitalLDOLogic_VIA1 $T=183190 25300 0 0 $X=182940 $Y=25070
X4440 1 DigitalLDOLogic_VIA1 $T=183190 29380 0 0 $X=182940 $Y=29150
X4441 1 DigitalLDOLogic_VIA1 $T=183190 33460 0 0 $X=182940 $Y=33230
X4442 1 DigitalLDOLogic_VIA1 $T=183190 37540 0 0 $X=182940 $Y=37310
X4443 1 DigitalLDOLogic_VIA1 $T=183190 41620 0 0 $X=182940 $Y=41390
X4444 1 DigitalLDOLogic_VIA1 $T=183190 45700 0 0 $X=182940 $Y=45470
X4445 1 DigitalLDOLogic_VIA1 $T=183190 49780 0 0 $X=182940 $Y=49550
X4446 1 DigitalLDOLogic_VIA1 $T=183190 53860 0 0 $X=182940 $Y=53630
X4447 1 DigitalLDOLogic_VIA1 $T=183190 57940 0 0 $X=182940 $Y=57710
X4448 3 DigitalLDOLogic_VIA1 $T=185030 11700 0 0 $X=184780 $Y=11470
X4449 3 DigitalLDOLogic_VIA1 $T=185030 15780 0 0 $X=184780 $Y=15550
X4450 3 DigitalLDOLogic_VIA1 $T=185030 19860 0 0 $X=184780 $Y=19630
X4451 3 DigitalLDOLogic_VIA1 $T=185030 23940 0 0 $X=184780 $Y=23710
X4452 3 DigitalLDOLogic_VIA1 $T=185030 28020 0 0 $X=184780 $Y=27790
X4453 3 DigitalLDOLogic_VIA1 $T=185030 32100 0 0 $X=184780 $Y=31870
X4454 3 DigitalLDOLogic_VIA1 $T=185030 36180 0 0 $X=184780 $Y=35950
X4455 3 DigitalLDOLogic_VIA1 $T=185030 40260 0 0 $X=184780 $Y=40030
X4456 3 DigitalLDOLogic_VIA1 $T=185030 44340 0 0 $X=184780 $Y=44110
X4457 3 DigitalLDOLogic_VIA1 $T=185030 48420 0 0 $X=184780 $Y=48190
X4458 3 DigitalLDOLogic_VIA1 $T=185030 52500 0 0 $X=184780 $Y=52270
X4459 3 DigitalLDOLogic_VIA1 $T=185030 56580 0 0 $X=184780 $Y=56350
X4460 1 DigitalLDOLogic_VIA1 $T=185950 13060 0 0 $X=185700 $Y=12830
X4461 1 DigitalLDOLogic_VIA1 $T=185950 17140 0 0 $X=185700 $Y=16910
X4462 1 DigitalLDOLogic_VIA1 $T=185950 21220 0 0 $X=185700 $Y=20990
X4463 1 DigitalLDOLogic_VIA1 $T=185950 25300 0 0 $X=185700 $Y=25070
X4464 1 DigitalLDOLogic_VIA1 $T=185950 29380 0 0 $X=185700 $Y=29150
X4465 1 DigitalLDOLogic_VIA1 $T=185950 33460 0 0 $X=185700 $Y=33230
X4466 1 DigitalLDOLogic_VIA1 $T=185950 37540 0 0 $X=185700 $Y=37310
X4467 1 DigitalLDOLogic_VIA1 $T=185950 41620 0 0 $X=185700 $Y=41390
X4468 1 DigitalLDOLogic_VIA1 $T=185950 45700 0 0 $X=185700 $Y=45470
X4469 1 DigitalLDOLogic_VIA1 $T=185950 49780 0 0 $X=185700 $Y=49550
X4470 1 DigitalLDOLogic_VIA1 $T=185950 53860 0 0 $X=185700 $Y=53630
X4471 1 DigitalLDOLogic_VIA1 $T=185950 57940 0 0 $X=185700 $Y=57710
X4472 3 DigitalLDOLogic_VIA1 $T=187790 11700 0 0 $X=187540 $Y=11470
X4473 3 DigitalLDOLogic_VIA1 $T=187790 15780 0 0 $X=187540 $Y=15550
X4474 3 DigitalLDOLogic_VIA1 $T=187790 19860 0 0 $X=187540 $Y=19630
X4475 3 DigitalLDOLogic_VIA1 $T=187790 23940 0 0 $X=187540 $Y=23710
X4476 3 DigitalLDOLogic_VIA1 $T=187790 28020 0 0 $X=187540 $Y=27790
X4477 3 DigitalLDOLogic_VIA1 $T=187790 32100 0 0 $X=187540 $Y=31870
X4478 3 DigitalLDOLogic_VIA1 $T=187790 36180 0 0 $X=187540 $Y=35950
X4479 3 DigitalLDOLogic_VIA1 $T=187790 40260 0 0 $X=187540 $Y=40030
X4480 3 DigitalLDOLogic_VIA1 $T=187790 44340 0 0 $X=187540 $Y=44110
X4481 3 DigitalLDOLogic_VIA1 $T=187790 48420 0 0 $X=187540 $Y=48190
X4482 3 DigitalLDOLogic_VIA1 $T=187790 52500 0 0 $X=187540 $Y=52270
X4483 3 DigitalLDOLogic_VIA1 $T=187790 56580 0 0 $X=187540 $Y=56350
X4484 1 DigitalLDOLogic_VIA1 $T=188710 13060 0 0 $X=188460 $Y=12830
X4485 1 DigitalLDOLogic_VIA1 $T=188710 17140 0 0 $X=188460 $Y=16910
X4486 1 DigitalLDOLogic_VIA1 $T=188710 21220 0 0 $X=188460 $Y=20990
X4487 1 DigitalLDOLogic_VIA1 $T=188710 25300 0 0 $X=188460 $Y=25070
X4488 1 DigitalLDOLogic_VIA1 $T=188710 29380 0 0 $X=188460 $Y=29150
X4489 1 DigitalLDOLogic_VIA1 $T=188710 33460 0 0 $X=188460 $Y=33230
X4490 1 DigitalLDOLogic_VIA1 $T=188710 37540 0 0 $X=188460 $Y=37310
X4491 1 DigitalLDOLogic_VIA1 $T=188710 41620 0 0 $X=188460 $Y=41390
X4492 1 DigitalLDOLogic_VIA1 $T=188710 45700 0 0 $X=188460 $Y=45470
X4493 1 DigitalLDOLogic_VIA1 $T=188710 49780 0 0 $X=188460 $Y=49550
X4494 1 DigitalLDOLogic_VIA1 $T=188710 53860 0 0 $X=188460 $Y=53630
X4495 1 DigitalLDOLogic_VIA1 $T=188710 57940 0 0 $X=188460 $Y=57710
X4496 3 DigitalLDOLogic_VIA2 $T=12300 11700 0 0 $X=11830 $Y=11470
X4497 3 DigitalLDOLogic_VIA2 $T=12300 15780 0 0 $X=11830 $Y=15550
X4498 3 DigitalLDOLogic_VIA2 $T=12300 19860 0 0 $X=11830 $Y=19630
X4499 3 DigitalLDOLogic_VIA2 $T=12300 23940 0 0 $X=11830 $Y=23710
X4500 3 DigitalLDOLogic_VIA2 $T=12300 28020 0 0 $X=11830 $Y=27790
X4501 3 DigitalLDOLogic_VIA2 $T=12300 32100 0 0 $X=11830 $Y=31870
X4502 3 DigitalLDOLogic_VIA2 $T=12300 36180 0 0 $X=11830 $Y=35950
X4503 3 DigitalLDOLogic_VIA2 $T=12300 40260 0 0 $X=11830 $Y=40030
X4504 3 DigitalLDOLogic_VIA2 $T=12300 44340 0 0 $X=11830 $Y=44110
X4505 3 DigitalLDOLogic_VIA2 $T=12300 48420 0 0 $X=11830 $Y=48190
X4506 3 DigitalLDOLogic_VIA2 $T=12300 52500 0 0 $X=11830 $Y=52270
X4507 3 DigitalLDOLogic_VIA2 $T=12300 56580 0 0 $X=11830 $Y=56350
X4508 1 DigitalLDOLogic_VIA2 $T=14140 13060 0 0 $X=13670 $Y=12830
X4509 1 DigitalLDOLogic_VIA2 $T=14140 17140 0 0 $X=13670 $Y=16910
X4510 1 DigitalLDOLogic_VIA2 $T=14140 21220 0 0 $X=13670 $Y=20990
X4511 1 DigitalLDOLogic_VIA2 $T=14140 25300 0 0 $X=13670 $Y=25070
X4512 1 DigitalLDOLogic_VIA2 $T=14140 29380 0 0 $X=13670 $Y=29150
X4513 1 DigitalLDOLogic_VIA2 $T=14140 33460 0 0 $X=13670 $Y=33230
X4514 1 DigitalLDOLogic_VIA2 $T=14140 37540 0 0 $X=13670 $Y=37310
X4515 1 DigitalLDOLogic_VIA2 $T=14140 41620 0 0 $X=13670 $Y=41390
X4516 1 DigitalLDOLogic_VIA2 $T=14140 45700 0 0 $X=13670 $Y=45470
X4517 1 DigitalLDOLogic_VIA2 $T=14140 49780 0 0 $X=13670 $Y=49550
X4518 1 DigitalLDOLogic_VIA2 $T=14140 53860 0 0 $X=13670 $Y=53630
X4519 1 DigitalLDOLogic_VIA2 $T=14140 57940 0 0 $X=13670 $Y=57710
X4520 3 DigitalLDOLogic_VIA2 $T=17820 11700 0 0 $X=17350 $Y=11470
X4521 3 DigitalLDOLogic_VIA2 $T=17820 15780 0 0 $X=17350 $Y=15550
X4522 3 DigitalLDOLogic_VIA2 $T=17820 19860 0 0 $X=17350 $Y=19630
X4523 3 DigitalLDOLogic_VIA2 $T=17820 23940 0 0 $X=17350 $Y=23710
X4524 3 DigitalLDOLogic_VIA2 $T=17820 28020 0 0 $X=17350 $Y=27790
X4525 3 DigitalLDOLogic_VIA2 $T=17820 32100 0 0 $X=17350 $Y=31870
X4526 3 DigitalLDOLogic_VIA2 $T=17820 36180 0 0 $X=17350 $Y=35950
X4527 3 DigitalLDOLogic_VIA2 $T=17820 40260 0 0 $X=17350 $Y=40030
X4528 3 DigitalLDOLogic_VIA2 $T=17820 44340 0 0 $X=17350 $Y=44110
X4529 3 DigitalLDOLogic_VIA2 $T=17820 48420 0 0 $X=17350 $Y=48190
X4530 3 DigitalLDOLogic_VIA2 $T=17820 52500 0 0 $X=17350 $Y=52270
X4531 3 DigitalLDOLogic_VIA2 $T=17820 56580 0 0 $X=17350 $Y=56350
X4532 1 DigitalLDOLogic_VIA2 $T=19660 13060 0 0 $X=19190 $Y=12830
X4533 1 DigitalLDOLogic_VIA2 $T=19660 17140 0 0 $X=19190 $Y=16910
X4534 1 DigitalLDOLogic_VIA2 $T=19660 21220 0 0 $X=19190 $Y=20990
X4535 1 DigitalLDOLogic_VIA2 $T=19660 25300 0 0 $X=19190 $Y=25070
X4536 1 DigitalLDOLogic_VIA2 $T=19660 29380 0 0 $X=19190 $Y=29150
X4537 1 DigitalLDOLogic_VIA2 $T=19660 33460 0 0 $X=19190 $Y=33230
X4538 1 DigitalLDOLogic_VIA2 $T=19660 37540 0 0 $X=19190 $Y=37310
X4539 1 DigitalLDOLogic_VIA2 $T=19660 41620 0 0 $X=19190 $Y=41390
X4540 1 DigitalLDOLogic_VIA2 $T=19660 45700 0 0 $X=19190 $Y=45470
X4541 1 DigitalLDOLogic_VIA2 $T=19660 49780 0 0 $X=19190 $Y=49550
X4542 1 DigitalLDOLogic_VIA2 $T=19660 53860 0 0 $X=19190 $Y=53630
X4543 1 DigitalLDOLogic_VIA2 $T=19660 57940 0 0 $X=19190 $Y=57710
X4544 3 DigitalLDOLogic_VIA2 $T=23340 11700 0 0 $X=22870 $Y=11470
X4545 3 DigitalLDOLogic_VIA2 $T=23340 15780 0 0 $X=22870 $Y=15550
X4546 3 DigitalLDOLogic_VIA2 $T=23340 19860 0 0 $X=22870 $Y=19630
X4547 3 DigitalLDOLogic_VIA2 $T=23340 23940 0 0 $X=22870 $Y=23710
X4548 3 DigitalLDOLogic_VIA2 $T=23340 28020 0 0 $X=22870 $Y=27790
X4549 3 DigitalLDOLogic_VIA2 $T=23340 32100 0 0 $X=22870 $Y=31870
X4550 3 DigitalLDOLogic_VIA2 $T=23340 36180 0 0 $X=22870 $Y=35950
X4551 3 DigitalLDOLogic_VIA2 $T=23340 40260 0 0 $X=22870 $Y=40030
X4552 3 DigitalLDOLogic_VIA2 $T=23340 44340 0 0 $X=22870 $Y=44110
X4553 3 DigitalLDOLogic_VIA2 $T=23340 48420 0 0 $X=22870 $Y=48190
X4554 3 DigitalLDOLogic_VIA2 $T=23340 52500 0 0 $X=22870 $Y=52270
X4555 3 DigitalLDOLogic_VIA2 $T=23340 56580 0 0 $X=22870 $Y=56350
X4556 1 DigitalLDOLogic_VIA2 $T=25180 13060 0 0 $X=24710 $Y=12830
X4557 1 DigitalLDOLogic_VIA2 $T=25180 17140 0 0 $X=24710 $Y=16910
X4558 1 DigitalLDOLogic_VIA2 $T=25180 21220 0 0 $X=24710 $Y=20990
X4559 1 DigitalLDOLogic_VIA2 $T=25180 25300 0 0 $X=24710 $Y=25070
X4560 1 DigitalLDOLogic_VIA2 $T=25180 29380 0 0 $X=24710 $Y=29150
X4561 1 DigitalLDOLogic_VIA2 $T=25180 33460 0 0 $X=24710 $Y=33230
X4562 1 DigitalLDOLogic_VIA2 $T=25180 37540 0 0 $X=24710 $Y=37310
X4563 1 DigitalLDOLogic_VIA2 $T=25180 41620 0 0 $X=24710 $Y=41390
X4564 1 DigitalLDOLogic_VIA2 $T=25180 45700 0 0 $X=24710 $Y=45470
X4565 1 DigitalLDOLogic_VIA2 $T=25180 49780 0 0 $X=24710 $Y=49550
X4566 1 DigitalLDOLogic_VIA2 $T=25180 53860 0 0 $X=24710 $Y=53630
X4567 1 DigitalLDOLogic_VIA2 $T=25180 57940 0 0 $X=24710 $Y=57710
X4568 3 DigitalLDOLogic_VIA2 $T=28860 11700 0 0 $X=28390 $Y=11470
X4569 3 DigitalLDOLogic_VIA2 $T=28860 15780 0 0 $X=28390 $Y=15550
X4570 3 DigitalLDOLogic_VIA2 $T=28860 19860 0 0 $X=28390 $Y=19630
X4571 3 DigitalLDOLogic_VIA2 $T=28860 23940 0 0 $X=28390 $Y=23710
X4572 3 DigitalLDOLogic_VIA2 $T=28860 28020 0 0 $X=28390 $Y=27790
X4573 3 DigitalLDOLogic_VIA2 $T=28860 32100 0 0 $X=28390 $Y=31870
X4574 3 DigitalLDOLogic_VIA2 $T=28860 36180 0 0 $X=28390 $Y=35950
X4575 3 DigitalLDOLogic_VIA2 $T=28860 40260 0 0 $X=28390 $Y=40030
X4576 3 DigitalLDOLogic_VIA2 $T=28860 44340 0 0 $X=28390 $Y=44110
X4577 3 DigitalLDOLogic_VIA2 $T=28860 48420 0 0 $X=28390 $Y=48190
X4578 3 DigitalLDOLogic_VIA2 $T=28860 52500 0 0 $X=28390 $Y=52270
X4579 3 DigitalLDOLogic_VIA2 $T=28860 56580 0 0 $X=28390 $Y=56350
X4580 1 DigitalLDOLogic_VIA2 $T=30700 13060 0 0 $X=30230 $Y=12830
X4581 1 DigitalLDOLogic_VIA2 $T=30700 17140 0 0 $X=30230 $Y=16910
X4582 1 DigitalLDOLogic_VIA2 $T=30700 21220 0 0 $X=30230 $Y=20990
X4583 1 DigitalLDOLogic_VIA2 $T=30700 25300 0 0 $X=30230 $Y=25070
X4584 1 DigitalLDOLogic_VIA2 $T=30700 29380 0 0 $X=30230 $Y=29150
X4585 1 DigitalLDOLogic_VIA2 $T=30700 33460 0 0 $X=30230 $Y=33230
X4586 1 DigitalLDOLogic_VIA2 $T=30700 37540 0 0 $X=30230 $Y=37310
X4587 1 DigitalLDOLogic_VIA2 $T=30700 41620 0 0 $X=30230 $Y=41390
X4588 1 DigitalLDOLogic_VIA2 $T=30700 45700 0 0 $X=30230 $Y=45470
X4589 1 DigitalLDOLogic_VIA2 $T=30700 49780 0 0 $X=30230 $Y=49550
X4590 1 DigitalLDOLogic_VIA2 $T=30700 53860 0 0 $X=30230 $Y=53630
X4591 1 DigitalLDOLogic_VIA2 $T=30700 57940 0 0 $X=30230 $Y=57710
X4592 3 DigitalLDOLogic_VIA2 $T=34380 11700 0 0 $X=33910 $Y=11470
X4593 3 DigitalLDOLogic_VIA2 $T=34380 15780 0 0 $X=33910 $Y=15550
X4594 3 DigitalLDOLogic_VIA2 $T=34380 19860 0 0 $X=33910 $Y=19630
X4595 3 DigitalLDOLogic_VIA2 $T=34380 23940 0 0 $X=33910 $Y=23710
X4596 3 DigitalLDOLogic_VIA2 $T=34380 28020 0 0 $X=33910 $Y=27790
X4597 3 DigitalLDOLogic_VIA2 $T=34380 32100 0 0 $X=33910 $Y=31870
X4598 3 DigitalLDOLogic_VIA2 $T=34380 36180 0 0 $X=33910 $Y=35950
X4599 3 DigitalLDOLogic_VIA2 $T=34380 40260 0 0 $X=33910 $Y=40030
X4600 3 DigitalLDOLogic_VIA2 $T=34380 44340 0 0 $X=33910 $Y=44110
X4601 3 DigitalLDOLogic_VIA2 $T=34380 48420 0 0 $X=33910 $Y=48190
X4602 3 DigitalLDOLogic_VIA2 $T=34380 52500 0 0 $X=33910 $Y=52270
X4603 3 DigitalLDOLogic_VIA2 $T=34380 56580 0 0 $X=33910 $Y=56350
X4604 1 DigitalLDOLogic_VIA2 $T=36220 13060 0 0 $X=35750 $Y=12830
X4605 1 DigitalLDOLogic_VIA2 $T=36220 17140 0 0 $X=35750 $Y=16910
X4606 1 DigitalLDOLogic_VIA2 $T=36220 21220 0 0 $X=35750 $Y=20990
X4607 1 DigitalLDOLogic_VIA2 $T=36220 25300 0 0 $X=35750 $Y=25070
X4608 1 DigitalLDOLogic_VIA2 $T=36220 29380 0 0 $X=35750 $Y=29150
X4609 1 DigitalLDOLogic_VIA2 $T=36220 33460 0 0 $X=35750 $Y=33230
X4610 1 DigitalLDOLogic_VIA2 $T=36220 37540 0 0 $X=35750 $Y=37310
X4611 1 DigitalLDOLogic_VIA2 $T=36220 41620 0 0 $X=35750 $Y=41390
X4612 1 DigitalLDOLogic_VIA2 $T=36220 45700 0 0 $X=35750 $Y=45470
X4613 1 DigitalLDOLogic_VIA2 $T=36220 49780 0 0 $X=35750 $Y=49550
X4614 1 DigitalLDOLogic_VIA2 $T=36220 53860 0 0 $X=35750 $Y=53630
X4615 1 DigitalLDOLogic_VIA2 $T=36220 57940 0 0 $X=35750 $Y=57710
X4616 3 DigitalLDOLogic_VIA2 $T=39900 11700 0 0 $X=39430 $Y=11470
X4617 3 DigitalLDOLogic_VIA2 $T=39900 15780 0 0 $X=39430 $Y=15550
X4618 3 DigitalLDOLogic_VIA2 $T=39900 19860 0 0 $X=39430 $Y=19630
X4619 3 DigitalLDOLogic_VIA2 $T=39900 23940 0 0 $X=39430 $Y=23710
X4620 3 DigitalLDOLogic_VIA2 $T=39900 28020 0 0 $X=39430 $Y=27790
X4621 3 DigitalLDOLogic_VIA2 $T=39900 32100 0 0 $X=39430 $Y=31870
X4622 3 DigitalLDOLogic_VIA2 $T=39900 36180 0 0 $X=39430 $Y=35950
X4623 3 DigitalLDOLogic_VIA2 $T=39900 40260 0 0 $X=39430 $Y=40030
X4624 3 DigitalLDOLogic_VIA2 $T=39900 44340 0 0 $X=39430 $Y=44110
X4625 3 DigitalLDOLogic_VIA2 $T=39900 48420 0 0 $X=39430 $Y=48190
X4626 3 DigitalLDOLogic_VIA2 $T=39900 52500 0 0 $X=39430 $Y=52270
X4627 3 DigitalLDOLogic_VIA2 $T=39900 56580 0 0 $X=39430 $Y=56350
X4628 1 DigitalLDOLogic_VIA2 $T=41740 13060 0 0 $X=41270 $Y=12830
X4629 1 DigitalLDOLogic_VIA2 $T=41740 17140 0 0 $X=41270 $Y=16910
X4630 1 DigitalLDOLogic_VIA2 $T=41740 21220 0 0 $X=41270 $Y=20990
X4631 1 DigitalLDOLogic_VIA2 $T=41740 25300 0 0 $X=41270 $Y=25070
X4632 1 DigitalLDOLogic_VIA2 $T=41740 29380 0 0 $X=41270 $Y=29150
X4633 1 DigitalLDOLogic_VIA2 $T=41740 33460 0 0 $X=41270 $Y=33230
X4634 1 DigitalLDOLogic_VIA2 $T=41740 37540 0 0 $X=41270 $Y=37310
X4635 1 DigitalLDOLogic_VIA2 $T=41740 41620 0 0 $X=41270 $Y=41390
X4636 1 DigitalLDOLogic_VIA2 $T=41740 45700 0 0 $X=41270 $Y=45470
X4637 1 DigitalLDOLogic_VIA2 $T=41740 49780 0 0 $X=41270 $Y=49550
X4638 1 DigitalLDOLogic_VIA2 $T=41740 53860 0 0 $X=41270 $Y=53630
X4639 1 DigitalLDOLogic_VIA2 $T=41740 57940 0 0 $X=41270 $Y=57710
X4640 3 DigitalLDOLogic_VIA2 $T=45420 11700 0 0 $X=44950 $Y=11470
X4641 3 DigitalLDOLogic_VIA2 $T=45420 15780 0 0 $X=44950 $Y=15550
X4642 3 DigitalLDOLogic_VIA2 $T=45420 19860 0 0 $X=44950 $Y=19630
X4643 3 DigitalLDOLogic_VIA2 $T=45420 23940 0 0 $X=44950 $Y=23710
X4644 3 DigitalLDOLogic_VIA2 $T=45420 28020 0 0 $X=44950 $Y=27790
X4645 3 DigitalLDOLogic_VIA2 $T=45420 32100 0 0 $X=44950 $Y=31870
X4646 3 DigitalLDOLogic_VIA2 $T=45420 36180 0 0 $X=44950 $Y=35950
X4647 3 DigitalLDOLogic_VIA2 $T=45420 40260 0 0 $X=44950 $Y=40030
X4648 3 DigitalLDOLogic_VIA2 $T=45420 44340 0 0 $X=44950 $Y=44110
X4649 3 DigitalLDOLogic_VIA2 $T=45420 48420 0 0 $X=44950 $Y=48190
X4650 3 DigitalLDOLogic_VIA2 $T=45420 52500 0 0 $X=44950 $Y=52270
X4651 3 DigitalLDOLogic_VIA2 $T=45420 56580 0 0 $X=44950 $Y=56350
X4652 1 DigitalLDOLogic_VIA2 $T=47260 13060 0 0 $X=46790 $Y=12830
X4653 1 DigitalLDOLogic_VIA2 $T=47260 17140 0 0 $X=46790 $Y=16910
X4654 1 DigitalLDOLogic_VIA2 $T=47260 21220 0 0 $X=46790 $Y=20990
X4655 1 DigitalLDOLogic_VIA2 $T=47260 25300 0 0 $X=46790 $Y=25070
X4656 1 DigitalLDOLogic_VIA2 $T=47260 29380 0 0 $X=46790 $Y=29150
X4657 1 DigitalLDOLogic_VIA2 $T=47260 33460 0 0 $X=46790 $Y=33230
X4658 1 DigitalLDOLogic_VIA2 $T=47260 37540 0 0 $X=46790 $Y=37310
X4659 1 DigitalLDOLogic_VIA2 $T=47260 41620 0 0 $X=46790 $Y=41390
X4660 1 DigitalLDOLogic_VIA2 $T=47260 45700 0 0 $X=46790 $Y=45470
X4661 1 DigitalLDOLogic_VIA2 $T=47260 49780 0 0 $X=46790 $Y=49550
X4662 1 DigitalLDOLogic_VIA2 $T=47260 53860 0 0 $X=46790 $Y=53630
X4663 1 DigitalLDOLogic_VIA2 $T=47260 57940 0 0 $X=46790 $Y=57710
X4664 3 DigitalLDOLogic_VIA2 $T=50940 11700 0 0 $X=50470 $Y=11470
X4665 3 DigitalLDOLogic_VIA2 $T=50940 15780 0 0 $X=50470 $Y=15550
X4666 3 DigitalLDOLogic_VIA2 $T=50940 19860 0 0 $X=50470 $Y=19630
X4667 3 DigitalLDOLogic_VIA2 $T=50940 23940 0 0 $X=50470 $Y=23710
X4668 3 DigitalLDOLogic_VIA2 $T=50940 28020 0 0 $X=50470 $Y=27790
X4669 3 DigitalLDOLogic_VIA2 $T=50940 32100 0 0 $X=50470 $Y=31870
X4670 3 DigitalLDOLogic_VIA2 $T=50940 36180 0 0 $X=50470 $Y=35950
X4671 3 DigitalLDOLogic_VIA2 $T=50940 40260 0 0 $X=50470 $Y=40030
X4672 3 DigitalLDOLogic_VIA2 $T=50940 44340 0 0 $X=50470 $Y=44110
X4673 3 DigitalLDOLogic_VIA2 $T=50940 48420 0 0 $X=50470 $Y=48190
X4674 3 DigitalLDOLogic_VIA2 $T=50940 52500 0 0 $X=50470 $Y=52270
X4675 3 DigitalLDOLogic_VIA2 $T=50940 56580 0 0 $X=50470 $Y=56350
X4676 1 DigitalLDOLogic_VIA2 $T=52780 13060 0 0 $X=52310 $Y=12830
X4677 1 DigitalLDOLogic_VIA2 $T=52780 17140 0 0 $X=52310 $Y=16910
X4678 1 DigitalLDOLogic_VIA2 $T=52780 21220 0 0 $X=52310 $Y=20990
X4679 1 DigitalLDOLogic_VIA2 $T=52780 25300 0 0 $X=52310 $Y=25070
X4680 1 DigitalLDOLogic_VIA2 $T=52780 29380 0 0 $X=52310 $Y=29150
X4681 1 DigitalLDOLogic_VIA2 $T=52780 33460 0 0 $X=52310 $Y=33230
X4682 1 DigitalLDOLogic_VIA2 $T=52780 37540 0 0 $X=52310 $Y=37310
X4683 1 DigitalLDOLogic_VIA2 $T=52780 41620 0 0 $X=52310 $Y=41390
X4684 1 DigitalLDOLogic_VIA2 $T=52780 45700 0 0 $X=52310 $Y=45470
X4685 1 DigitalLDOLogic_VIA2 $T=52780 49780 0 0 $X=52310 $Y=49550
X4686 1 DigitalLDOLogic_VIA2 $T=52780 53860 0 0 $X=52310 $Y=53630
X4687 1 DigitalLDOLogic_VIA2 $T=52780 57940 0 0 $X=52310 $Y=57710
X4688 3 DigitalLDOLogic_VIA2 $T=56460 11700 0 0 $X=55990 $Y=11470
X4689 3 DigitalLDOLogic_VIA2 $T=56460 15780 0 0 $X=55990 $Y=15550
X4690 3 DigitalLDOLogic_VIA2 $T=56460 19860 0 0 $X=55990 $Y=19630
X4691 3 DigitalLDOLogic_VIA2 $T=56460 23940 0 0 $X=55990 $Y=23710
X4692 3 DigitalLDOLogic_VIA2 $T=56460 28020 0 0 $X=55990 $Y=27790
X4693 3 DigitalLDOLogic_VIA2 $T=56460 32100 0 0 $X=55990 $Y=31870
X4694 3 DigitalLDOLogic_VIA2 $T=56460 36180 0 0 $X=55990 $Y=35950
X4695 3 DigitalLDOLogic_VIA2 $T=56460 40260 0 0 $X=55990 $Y=40030
X4696 3 DigitalLDOLogic_VIA2 $T=56460 44340 0 0 $X=55990 $Y=44110
X4697 3 DigitalLDOLogic_VIA2 $T=56460 48420 0 0 $X=55990 $Y=48190
X4698 3 DigitalLDOLogic_VIA2 $T=56460 52500 0 0 $X=55990 $Y=52270
X4699 3 DigitalLDOLogic_VIA2 $T=56460 56580 0 0 $X=55990 $Y=56350
X4700 1 DigitalLDOLogic_VIA2 $T=58300 13060 0 0 $X=57830 $Y=12830
X4701 1 DigitalLDOLogic_VIA2 $T=58300 17140 0 0 $X=57830 $Y=16910
X4702 1 DigitalLDOLogic_VIA2 $T=58300 21220 0 0 $X=57830 $Y=20990
X4703 1 DigitalLDOLogic_VIA2 $T=58300 25300 0 0 $X=57830 $Y=25070
X4704 1 DigitalLDOLogic_VIA2 $T=58300 29380 0 0 $X=57830 $Y=29150
X4705 1 DigitalLDOLogic_VIA2 $T=58300 33460 0 0 $X=57830 $Y=33230
X4706 1 DigitalLDOLogic_VIA2 $T=58300 37540 0 0 $X=57830 $Y=37310
X4707 1 DigitalLDOLogic_VIA2 $T=58300 41620 0 0 $X=57830 $Y=41390
X4708 1 DigitalLDOLogic_VIA2 $T=58300 45700 0 0 $X=57830 $Y=45470
X4709 1 DigitalLDOLogic_VIA2 $T=58300 49780 0 0 $X=57830 $Y=49550
X4710 1 DigitalLDOLogic_VIA2 $T=58300 53860 0 0 $X=57830 $Y=53630
X4711 1 DigitalLDOLogic_VIA2 $T=58300 57940 0 0 $X=57830 $Y=57710
X4712 3 DigitalLDOLogic_VIA2 $T=61980 11700 0 0 $X=61510 $Y=11470
X4713 3 DigitalLDOLogic_VIA2 $T=61980 15780 0 0 $X=61510 $Y=15550
X4714 3 DigitalLDOLogic_VIA2 $T=61980 19860 0 0 $X=61510 $Y=19630
X4715 3 DigitalLDOLogic_VIA2 $T=61980 23940 0 0 $X=61510 $Y=23710
X4716 3 DigitalLDOLogic_VIA2 $T=61980 28020 0 0 $X=61510 $Y=27790
X4717 3 DigitalLDOLogic_VIA2 $T=61980 32100 0 0 $X=61510 $Y=31870
X4718 3 DigitalLDOLogic_VIA2 $T=61980 36180 0 0 $X=61510 $Y=35950
X4719 3 DigitalLDOLogic_VIA2 $T=61980 40260 0 0 $X=61510 $Y=40030
X4720 3 DigitalLDOLogic_VIA2 $T=61980 44340 0 0 $X=61510 $Y=44110
X4721 3 DigitalLDOLogic_VIA2 $T=61980 48420 0 0 $X=61510 $Y=48190
X4722 3 DigitalLDOLogic_VIA2 $T=61980 52500 0 0 $X=61510 $Y=52270
X4723 3 DigitalLDOLogic_VIA2 $T=61980 56580 0 0 $X=61510 $Y=56350
X4724 1 DigitalLDOLogic_VIA2 $T=63820 13060 0 0 $X=63350 $Y=12830
X4725 1 DigitalLDOLogic_VIA2 $T=63820 17140 0 0 $X=63350 $Y=16910
X4726 1 DigitalLDOLogic_VIA2 $T=63820 21220 0 0 $X=63350 $Y=20990
X4727 1 DigitalLDOLogic_VIA2 $T=63820 25300 0 0 $X=63350 $Y=25070
X4728 1 DigitalLDOLogic_VIA2 $T=63820 29380 0 0 $X=63350 $Y=29150
X4729 1 DigitalLDOLogic_VIA2 $T=63820 33460 0 0 $X=63350 $Y=33230
X4730 1 DigitalLDOLogic_VIA2 $T=63820 37540 0 0 $X=63350 $Y=37310
X4731 1 DigitalLDOLogic_VIA2 $T=63820 41620 0 0 $X=63350 $Y=41390
X4732 1 DigitalLDOLogic_VIA2 $T=63820 45700 0 0 $X=63350 $Y=45470
X4733 1 DigitalLDOLogic_VIA2 $T=63820 49780 0 0 $X=63350 $Y=49550
X4734 1 DigitalLDOLogic_VIA2 $T=63820 53860 0 0 $X=63350 $Y=53630
X4735 1 DigitalLDOLogic_VIA2 $T=63820 57940 0 0 $X=63350 $Y=57710
X4736 3 DigitalLDOLogic_VIA2 $T=67500 11700 0 0 $X=67030 $Y=11470
X4737 3 DigitalLDOLogic_VIA2 $T=67500 15780 0 0 $X=67030 $Y=15550
X4738 3 DigitalLDOLogic_VIA2 $T=67500 19860 0 0 $X=67030 $Y=19630
X4739 3 DigitalLDOLogic_VIA2 $T=67500 23940 0 0 $X=67030 $Y=23710
X4740 3 DigitalLDOLogic_VIA2 $T=67500 28020 0 0 $X=67030 $Y=27790
X4741 3 DigitalLDOLogic_VIA2 $T=67500 32100 0 0 $X=67030 $Y=31870
X4742 3 DigitalLDOLogic_VIA2 $T=67500 36180 0 0 $X=67030 $Y=35950
X4743 3 DigitalLDOLogic_VIA2 $T=67500 40260 0 0 $X=67030 $Y=40030
X4744 3 DigitalLDOLogic_VIA2 $T=67500 44340 0 0 $X=67030 $Y=44110
X4745 3 DigitalLDOLogic_VIA2 $T=67500 48420 0 0 $X=67030 $Y=48190
X4746 3 DigitalLDOLogic_VIA2 $T=67500 52500 0 0 $X=67030 $Y=52270
X4747 3 DigitalLDOLogic_VIA2 $T=67500 56580 0 0 $X=67030 $Y=56350
X4748 1 DigitalLDOLogic_VIA2 $T=69340 13060 0 0 $X=68870 $Y=12830
X4749 1 DigitalLDOLogic_VIA2 $T=69340 17140 0 0 $X=68870 $Y=16910
X4750 1 DigitalLDOLogic_VIA2 $T=69340 21220 0 0 $X=68870 $Y=20990
X4751 1 DigitalLDOLogic_VIA2 $T=69340 25300 0 0 $X=68870 $Y=25070
X4752 1 DigitalLDOLogic_VIA2 $T=69340 29380 0 0 $X=68870 $Y=29150
X4753 1 DigitalLDOLogic_VIA2 $T=69340 33460 0 0 $X=68870 $Y=33230
X4754 1 DigitalLDOLogic_VIA2 $T=69340 37540 0 0 $X=68870 $Y=37310
X4755 1 DigitalLDOLogic_VIA2 $T=69340 41620 0 0 $X=68870 $Y=41390
X4756 1 DigitalLDOLogic_VIA2 $T=69340 45700 0 0 $X=68870 $Y=45470
X4757 1 DigitalLDOLogic_VIA2 $T=69340 49780 0 0 $X=68870 $Y=49550
X4758 1 DigitalLDOLogic_VIA2 $T=69340 53860 0 0 $X=68870 $Y=53630
X4759 1 DigitalLDOLogic_VIA2 $T=69340 57940 0 0 $X=68870 $Y=57710
X4760 3 DigitalLDOLogic_VIA2 $T=73020 11700 0 0 $X=72550 $Y=11470
X4761 3 DigitalLDOLogic_VIA2 $T=73020 15780 0 0 $X=72550 $Y=15550
X4762 3 DigitalLDOLogic_VIA2 $T=73020 19860 0 0 $X=72550 $Y=19630
X4763 3 DigitalLDOLogic_VIA2 $T=73020 23940 0 0 $X=72550 $Y=23710
X4764 3 DigitalLDOLogic_VIA2 $T=73020 28020 0 0 $X=72550 $Y=27790
X4765 3 DigitalLDOLogic_VIA2 $T=73020 32100 0 0 $X=72550 $Y=31870
X4766 3 DigitalLDOLogic_VIA2 $T=73020 36180 0 0 $X=72550 $Y=35950
X4767 3 DigitalLDOLogic_VIA2 $T=73020 40260 0 0 $X=72550 $Y=40030
X4768 3 DigitalLDOLogic_VIA2 $T=73020 44340 0 0 $X=72550 $Y=44110
X4769 3 DigitalLDOLogic_VIA2 $T=73020 48420 0 0 $X=72550 $Y=48190
X4770 3 DigitalLDOLogic_VIA2 $T=73020 52500 0 0 $X=72550 $Y=52270
X4771 3 DigitalLDOLogic_VIA2 $T=73020 56580 0 0 $X=72550 $Y=56350
X4772 1 DigitalLDOLogic_VIA2 $T=74860 13060 0 0 $X=74390 $Y=12830
X4773 1 DigitalLDOLogic_VIA2 $T=74860 17140 0 0 $X=74390 $Y=16910
X4774 1 DigitalLDOLogic_VIA2 $T=74860 21220 0 0 $X=74390 $Y=20990
X4775 1 DigitalLDOLogic_VIA2 $T=74860 25300 0 0 $X=74390 $Y=25070
X4776 1 DigitalLDOLogic_VIA2 $T=74860 29380 0 0 $X=74390 $Y=29150
X4777 1 DigitalLDOLogic_VIA2 $T=74860 33460 0 0 $X=74390 $Y=33230
X4778 1 DigitalLDOLogic_VIA2 $T=74860 37540 0 0 $X=74390 $Y=37310
X4779 1 DigitalLDOLogic_VIA2 $T=74860 41620 0 0 $X=74390 $Y=41390
X4780 1 DigitalLDOLogic_VIA2 $T=74860 45700 0 0 $X=74390 $Y=45470
X4781 1 DigitalLDOLogic_VIA2 $T=74860 49780 0 0 $X=74390 $Y=49550
X4782 1 DigitalLDOLogic_VIA2 $T=74860 53860 0 0 $X=74390 $Y=53630
X4783 1 DigitalLDOLogic_VIA2 $T=74860 57940 0 0 $X=74390 $Y=57710
X4784 3 DigitalLDOLogic_VIA2 $T=78540 11700 0 0 $X=78070 $Y=11470
X4785 3 DigitalLDOLogic_VIA2 $T=78540 15780 0 0 $X=78070 $Y=15550
X4786 3 DigitalLDOLogic_VIA2 $T=78540 19860 0 0 $X=78070 $Y=19630
X4787 3 DigitalLDOLogic_VIA2 $T=78540 23940 0 0 $X=78070 $Y=23710
X4788 3 DigitalLDOLogic_VIA2 $T=78540 28020 0 0 $X=78070 $Y=27790
X4789 3 DigitalLDOLogic_VIA2 $T=78540 32100 0 0 $X=78070 $Y=31870
X4790 3 DigitalLDOLogic_VIA2 $T=78540 36180 0 0 $X=78070 $Y=35950
X4791 3 DigitalLDOLogic_VIA2 $T=78540 40260 0 0 $X=78070 $Y=40030
X4792 3 DigitalLDOLogic_VIA2 $T=78540 44340 0 0 $X=78070 $Y=44110
X4793 3 DigitalLDOLogic_VIA2 $T=78540 48420 0 0 $X=78070 $Y=48190
X4794 3 DigitalLDOLogic_VIA2 $T=78540 52500 0 0 $X=78070 $Y=52270
X4795 3 DigitalLDOLogic_VIA2 $T=78540 56580 0 0 $X=78070 $Y=56350
X4796 1 DigitalLDOLogic_VIA2 $T=80380 13060 0 0 $X=79910 $Y=12830
X4797 1 DigitalLDOLogic_VIA2 $T=80380 17140 0 0 $X=79910 $Y=16910
X4798 1 DigitalLDOLogic_VIA2 $T=80380 21220 0 0 $X=79910 $Y=20990
X4799 1 DigitalLDOLogic_VIA2 $T=80380 25300 0 0 $X=79910 $Y=25070
X4800 1 DigitalLDOLogic_VIA2 $T=80380 29380 0 0 $X=79910 $Y=29150
X4801 1 DigitalLDOLogic_VIA2 $T=80380 33460 0 0 $X=79910 $Y=33230
X4802 1 DigitalLDOLogic_VIA2 $T=80380 37540 0 0 $X=79910 $Y=37310
X4803 1 DigitalLDOLogic_VIA2 $T=80380 41620 0 0 $X=79910 $Y=41390
X4804 1 DigitalLDOLogic_VIA2 $T=80380 45700 0 0 $X=79910 $Y=45470
X4805 1 DigitalLDOLogic_VIA2 $T=80380 49780 0 0 $X=79910 $Y=49550
X4806 1 DigitalLDOLogic_VIA2 $T=80380 53860 0 0 $X=79910 $Y=53630
X4807 1 DigitalLDOLogic_VIA2 $T=80380 57940 0 0 $X=79910 $Y=57710
X4808 3 DigitalLDOLogic_VIA2 $T=84060 11700 0 0 $X=83590 $Y=11470
X4809 3 DigitalLDOLogic_VIA2 $T=84060 15780 0 0 $X=83590 $Y=15550
X4810 3 DigitalLDOLogic_VIA2 $T=84060 19860 0 0 $X=83590 $Y=19630
X4811 3 DigitalLDOLogic_VIA2 $T=84060 23940 0 0 $X=83590 $Y=23710
X4812 3 DigitalLDOLogic_VIA2 $T=84060 28020 0 0 $X=83590 $Y=27790
X4813 3 DigitalLDOLogic_VIA2 $T=84060 32100 0 0 $X=83590 $Y=31870
X4814 3 DigitalLDOLogic_VIA2 $T=84060 36180 0 0 $X=83590 $Y=35950
X4815 3 DigitalLDOLogic_VIA2 $T=84060 40260 0 0 $X=83590 $Y=40030
X4816 3 DigitalLDOLogic_VIA2 $T=84060 44340 0 0 $X=83590 $Y=44110
X4817 3 DigitalLDOLogic_VIA2 $T=84060 48420 0 0 $X=83590 $Y=48190
X4818 3 DigitalLDOLogic_VIA2 $T=84060 52500 0 0 $X=83590 $Y=52270
X4819 3 DigitalLDOLogic_VIA2 $T=84060 56580 0 0 $X=83590 $Y=56350
X4820 1 DigitalLDOLogic_VIA2 $T=85900 13060 0 0 $X=85430 $Y=12830
X4821 1 DigitalLDOLogic_VIA2 $T=85900 17140 0 0 $X=85430 $Y=16910
X4822 1 DigitalLDOLogic_VIA2 $T=85900 21220 0 0 $X=85430 $Y=20990
X4823 1 DigitalLDOLogic_VIA2 $T=85900 25300 0 0 $X=85430 $Y=25070
X4824 1 DigitalLDOLogic_VIA2 $T=85900 29380 0 0 $X=85430 $Y=29150
X4825 1 DigitalLDOLogic_VIA2 $T=85900 33460 0 0 $X=85430 $Y=33230
X4826 1 DigitalLDOLogic_VIA2 $T=85900 37540 0 0 $X=85430 $Y=37310
X4827 1 DigitalLDOLogic_VIA2 $T=85900 41620 0 0 $X=85430 $Y=41390
X4828 1 DigitalLDOLogic_VIA2 $T=85900 45700 0 0 $X=85430 $Y=45470
X4829 1 DigitalLDOLogic_VIA2 $T=85900 49780 0 0 $X=85430 $Y=49550
X4830 1 DigitalLDOLogic_VIA2 $T=85900 53860 0 0 $X=85430 $Y=53630
X4831 1 DigitalLDOLogic_VIA2 $T=85900 57940 0 0 $X=85430 $Y=57710
X4832 3 DigitalLDOLogic_VIA2 $T=89580 11700 0 0 $X=89110 $Y=11470
X4833 3 DigitalLDOLogic_VIA2 $T=89580 15780 0 0 $X=89110 $Y=15550
X4834 3 DigitalLDOLogic_VIA2 $T=89580 19860 0 0 $X=89110 $Y=19630
X4835 3 DigitalLDOLogic_VIA2 $T=89580 23940 0 0 $X=89110 $Y=23710
X4836 3 DigitalLDOLogic_VIA2 $T=89580 28020 0 0 $X=89110 $Y=27790
X4837 3 DigitalLDOLogic_VIA2 $T=89580 32100 0 0 $X=89110 $Y=31870
X4838 3 DigitalLDOLogic_VIA2 $T=89580 36180 0 0 $X=89110 $Y=35950
X4839 3 DigitalLDOLogic_VIA2 $T=89580 40260 0 0 $X=89110 $Y=40030
X4840 3 DigitalLDOLogic_VIA2 $T=89580 44340 0 0 $X=89110 $Y=44110
X4841 3 DigitalLDOLogic_VIA2 $T=89580 48420 0 0 $X=89110 $Y=48190
X4842 3 DigitalLDOLogic_VIA2 $T=89580 52500 0 0 $X=89110 $Y=52270
X4843 3 DigitalLDOLogic_VIA2 $T=89580 56580 0 0 $X=89110 $Y=56350
X4844 1 DigitalLDOLogic_VIA2 $T=91420 13060 0 0 $X=90950 $Y=12830
X4845 1 DigitalLDOLogic_VIA2 $T=91420 17140 0 0 $X=90950 $Y=16910
X4846 1 DigitalLDOLogic_VIA2 $T=91420 21220 0 0 $X=90950 $Y=20990
X4847 1 DigitalLDOLogic_VIA2 $T=91420 25300 0 0 $X=90950 $Y=25070
X4848 1 DigitalLDOLogic_VIA2 $T=91420 29380 0 0 $X=90950 $Y=29150
X4849 1 DigitalLDOLogic_VIA2 $T=91420 33460 0 0 $X=90950 $Y=33230
X4850 1 DigitalLDOLogic_VIA2 $T=91420 37540 0 0 $X=90950 $Y=37310
X4851 1 DigitalLDOLogic_VIA2 $T=91420 41620 0 0 $X=90950 $Y=41390
X4852 1 DigitalLDOLogic_VIA2 $T=91420 45700 0 0 $X=90950 $Y=45470
X4853 1 DigitalLDOLogic_VIA2 $T=91420 49780 0 0 $X=90950 $Y=49550
X4854 1 DigitalLDOLogic_VIA2 $T=91420 53860 0 0 $X=90950 $Y=53630
X4855 1 DigitalLDOLogic_VIA2 $T=91420 57940 0 0 $X=90950 $Y=57710
X4856 3 DigitalLDOLogic_VIA2 $T=95100 11700 0 0 $X=94630 $Y=11470
X4857 3 DigitalLDOLogic_VIA2 $T=95100 15780 0 0 $X=94630 $Y=15550
X4858 3 DigitalLDOLogic_VIA2 $T=95100 19860 0 0 $X=94630 $Y=19630
X4859 3 DigitalLDOLogic_VIA2 $T=95100 23940 0 0 $X=94630 $Y=23710
X4860 3 DigitalLDOLogic_VIA2 $T=95100 28020 0 0 $X=94630 $Y=27790
X4861 3 DigitalLDOLogic_VIA2 $T=95100 32100 0 0 $X=94630 $Y=31870
X4862 3 DigitalLDOLogic_VIA2 $T=95100 36180 0 0 $X=94630 $Y=35950
X4863 3 DigitalLDOLogic_VIA2 $T=95100 40260 0 0 $X=94630 $Y=40030
X4864 3 DigitalLDOLogic_VIA2 $T=95100 44340 0 0 $X=94630 $Y=44110
X4865 3 DigitalLDOLogic_VIA2 $T=95100 48420 0 0 $X=94630 $Y=48190
X4866 3 DigitalLDOLogic_VIA2 $T=95100 52500 0 0 $X=94630 $Y=52270
X4867 3 DigitalLDOLogic_VIA2 $T=95100 56580 0 0 $X=94630 $Y=56350
X4868 1 DigitalLDOLogic_VIA2 $T=96940 13060 0 0 $X=96470 $Y=12830
X4869 1 DigitalLDOLogic_VIA2 $T=96940 17140 0 0 $X=96470 $Y=16910
X4870 1 DigitalLDOLogic_VIA2 $T=96940 21220 0 0 $X=96470 $Y=20990
X4871 1 DigitalLDOLogic_VIA2 $T=96940 25300 0 0 $X=96470 $Y=25070
X4872 1 DigitalLDOLogic_VIA2 $T=96940 29380 0 0 $X=96470 $Y=29150
X4873 1 DigitalLDOLogic_VIA2 $T=96940 33460 0 0 $X=96470 $Y=33230
X4874 1 DigitalLDOLogic_VIA2 $T=96940 37540 0 0 $X=96470 $Y=37310
X4875 1 DigitalLDOLogic_VIA2 $T=96940 41620 0 0 $X=96470 $Y=41390
X4876 1 DigitalLDOLogic_VIA2 $T=96940 45700 0 0 $X=96470 $Y=45470
X4877 1 DigitalLDOLogic_VIA2 $T=96940 49780 0 0 $X=96470 $Y=49550
X4878 1 DigitalLDOLogic_VIA2 $T=96940 53860 0 0 $X=96470 $Y=53630
X4879 1 DigitalLDOLogic_VIA2 $T=96940 57940 0 0 $X=96470 $Y=57710
X4880 3 DigitalLDOLogic_VIA2 $T=100620 11700 0 0 $X=100150 $Y=11470
X4881 3 DigitalLDOLogic_VIA2 $T=100620 15780 0 0 $X=100150 $Y=15550
X4882 3 DigitalLDOLogic_VIA2 $T=100620 19860 0 0 $X=100150 $Y=19630
X4883 3 DigitalLDOLogic_VIA2 $T=100620 23940 0 0 $X=100150 $Y=23710
X4884 3 DigitalLDOLogic_VIA2 $T=100620 28020 0 0 $X=100150 $Y=27790
X4885 3 DigitalLDOLogic_VIA2 $T=100620 32100 0 0 $X=100150 $Y=31870
X4886 3 DigitalLDOLogic_VIA2 $T=100620 36180 0 0 $X=100150 $Y=35950
X4887 3 DigitalLDOLogic_VIA2 $T=100620 40260 0 0 $X=100150 $Y=40030
X4888 3 DigitalLDOLogic_VIA2 $T=100620 44340 0 0 $X=100150 $Y=44110
X4889 3 DigitalLDOLogic_VIA2 $T=100620 48420 0 0 $X=100150 $Y=48190
X4890 3 DigitalLDOLogic_VIA2 $T=100620 52500 0 0 $X=100150 $Y=52270
X4891 3 DigitalLDOLogic_VIA2 $T=100620 56580 0 0 $X=100150 $Y=56350
X4892 1 DigitalLDOLogic_VIA2 $T=102460 13060 0 0 $X=101990 $Y=12830
X4893 1 DigitalLDOLogic_VIA2 $T=102460 17140 0 0 $X=101990 $Y=16910
X4894 1 DigitalLDOLogic_VIA2 $T=102460 21220 0 0 $X=101990 $Y=20990
X4895 1 DigitalLDOLogic_VIA2 $T=102460 25300 0 0 $X=101990 $Y=25070
X4896 1 DigitalLDOLogic_VIA2 $T=102460 29380 0 0 $X=101990 $Y=29150
X4897 1 DigitalLDOLogic_VIA2 $T=102460 33460 0 0 $X=101990 $Y=33230
X4898 1 DigitalLDOLogic_VIA2 $T=102460 37540 0 0 $X=101990 $Y=37310
X4899 1 DigitalLDOLogic_VIA2 $T=102460 41620 0 0 $X=101990 $Y=41390
X4900 1 DigitalLDOLogic_VIA2 $T=102460 45700 0 0 $X=101990 $Y=45470
X4901 1 DigitalLDOLogic_VIA2 $T=102460 49780 0 0 $X=101990 $Y=49550
X4902 1 DigitalLDOLogic_VIA2 $T=102460 53860 0 0 $X=101990 $Y=53630
X4903 1 DigitalLDOLogic_VIA2 $T=102460 57940 0 0 $X=101990 $Y=57710
X4904 3 DigitalLDOLogic_VIA2 $T=106140 11700 0 0 $X=105670 $Y=11470
X4905 3 DigitalLDOLogic_VIA2 $T=106140 15780 0 0 $X=105670 $Y=15550
X4906 3 DigitalLDOLogic_VIA2 $T=106140 19860 0 0 $X=105670 $Y=19630
X4907 3 DigitalLDOLogic_VIA2 $T=106140 23940 0 0 $X=105670 $Y=23710
X4908 3 DigitalLDOLogic_VIA2 $T=106140 28020 0 0 $X=105670 $Y=27790
X4909 3 DigitalLDOLogic_VIA2 $T=106140 32100 0 0 $X=105670 $Y=31870
X4910 3 DigitalLDOLogic_VIA2 $T=106140 36180 0 0 $X=105670 $Y=35950
X4911 3 DigitalLDOLogic_VIA2 $T=106140 40260 0 0 $X=105670 $Y=40030
X4912 3 DigitalLDOLogic_VIA2 $T=106140 44340 0 0 $X=105670 $Y=44110
X4913 3 DigitalLDOLogic_VIA2 $T=106140 48420 0 0 $X=105670 $Y=48190
X4914 3 DigitalLDOLogic_VIA2 $T=106140 52500 0 0 $X=105670 $Y=52270
X4915 3 DigitalLDOLogic_VIA2 $T=106140 56580 0 0 $X=105670 $Y=56350
X4916 1 DigitalLDOLogic_VIA2 $T=107980 13060 0 0 $X=107510 $Y=12830
X4917 1 DigitalLDOLogic_VIA2 $T=107980 17140 0 0 $X=107510 $Y=16910
X4918 1 DigitalLDOLogic_VIA2 $T=107980 21220 0 0 $X=107510 $Y=20990
X4919 1 DigitalLDOLogic_VIA2 $T=107980 25300 0 0 $X=107510 $Y=25070
X4920 1 DigitalLDOLogic_VIA2 $T=107980 29380 0 0 $X=107510 $Y=29150
X4921 1 DigitalLDOLogic_VIA2 $T=107980 33460 0 0 $X=107510 $Y=33230
X4922 1 DigitalLDOLogic_VIA2 $T=107980 37540 0 0 $X=107510 $Y=37310
X4923 1 DigitalLDOLogic_VIA2 $T=107980 41620 0 0 $X=107510 $Y=41390
X4924 1 DigitalLDOLogic_VIA2 $T=107980 45700 0 0 $X=107510 $Y=45470
X4925 1 DigitalLDOLogic_VIA2 $T=107980 49780 0 0 $X=107510 $Y=49550
X4926 1 DigitalLDOLogic_VIA2 $T=107980 53860 0 0 $X=107510 $Y=53630
X4927 1 DigitalLDOLogic_VIA2 $T=107980 57940 0 0 $X=107510 $Y=57710
X4928 3 DigitalLDOLogic_VIA2 $T=111660 11700 0 0 $X=111190 $Y=11470
X4929 3 DigitalLDOLogic_VIA2 $T=111660 15780 0 0 $X=111190 $Y=15550
X4930 3 DigitalLDOLogic_VIA2 $T=111660 19860 0 0 $X=111190 $Y=19630
X4931 3 DigitalLDOLogic_VIA2 $T=111660 23940 0 0 $X=111190 $Y=23710
X4932 3 DigitalLDOLogic_VIA2 $T=111660 28020 0 0 $X=111190 $Y=27790
X4933 3 DigitalLDOLogic_VIA2 $T=111660 32100 0 0 $X=111190 $Y=31870
X4934 3 DigitalLDOLogic_VIA2 $T=111660 36180 0 0 $X=111190 $Y=35950
X4935 3 DigitalLDOLogic_VIA2 $T=111660 40260 0 0 $X=111190 $Y=40030
X4936 3 DigitalLDOLogic_VIA2 $T=111660 44340 0 0 $X=111190 $Y=44110
X4937 3 DigitalLDOLogic_VIA2 $T=111660 48420 0 0 $X=111190 $Y=48190
X4938 3 DigitalLDOLogic_VIA2 $T=111660 52500 0 0 $X=111190 $Y=52270
X4939 3 DigitalLDOLogic_VIA2 $T=111660 56580 0 0 $X=111190 $Y=56350
X4940 1 DigitalLDOLogic_VIA2 $T=113500 13060 0 0 $X=113030 $Y=12830
X4941 1 DigitalLDOLogic_VIA2 $T=113500 17140 0 0 $X=113030 $Y=16910
X4942 1 DigitalLDOLogic_VIA2 $T=113500 21220 0 0 $X=113030 $Y=20990
X4943 1 DigitalLDOLogic_VIA2 $T=113500 25300 0 0 $X=113030 $Y=25070
X4944 1 DigitalLDOLogic_VIA2 $T=113500 29380 0 0 $X=113030 $Y=29150
X4945 1 DigitalLDOLogic_VIA2 $T=113500 33460 0 0 $X=113030 $Y=33230
X4946 1 DigitalLDOLogic_VIA2 $T=113500 37540 0 0 $X=113030 $Y=37310
X4947 1 DigitalLDOLogic_VIA2 $T=113500 41620 0 0 $X=113030 $Y=41390
X4948 1 DigitalLDOLogic_VIA2 $T=113500 45700 0 0 $X=113030 $Y=45470
X4949 1 DigitalLDOLogic_VIA2 $T=113500 49780 0 0 $X=113030 $Y=49550
X4950 1 DigitalLDOLogic_VIA2 $T=113500 53860 0 0 $X=113030 $Y=53630
X4951 1 DigitalLDOLogic_VIA2 $T=113500 57940 0 0 $X=113030 $Y=57710
X4952 3 DigitalLDOLogic_VIA2 $T=117180 11700 0 0 $X=116710 $Y=11470
X4953 3 DigitalLDOLogic_VIA2 $T=117180 15780 0 0 $X=116710 $Y=15550
X4954 3 DigitalLDOLogic_VIA2 $T=117180 19860 0 0 $X=116710 $Y=19630
X4955 3 DigitalLDOLogic_VIA2 $T=117180 23940 0 0 $X=116710 $Y=23710
X4956 3 DigitalLDOLogic_VIA2 $T=117180 28020 0 0 $X=116710 $Y=27790
X4957 3 DigitalLDOLogic_VIA2 $T=117180 32100 0 0 $X=116710 $Y=31870
X4958 3 DigitalLDOLogic_VIA2 $T=117180 36180 0 0 $X=116710 $Y=35950
X4959 3 DigitalLDOLogic_VIA2 $T=117180 40260 0 0 $X=116710 $Y=40030
X4960 3 DigitalLDOLogic_VIA2 $T=117180 44340 0 0 $X=116710 $Y=44110
X4961 3 DigitalLDOLogic_VIA2 $T=117180 48420 0 0 $X=116710 $Y=48190
X4962 3 DigitalLDOLogic_VIA2 $T=117180 52500 0 0 $X=116710 $Y=52270
X4963 3 DigitalLDOLogic_VIA2 $T=117180 56580 0 0 $X=116710 $Y=56350
X4964 1 DigitalLDOLogic_VIA2 $T=119020 13060 0 0 $X=118550 $Y=12830
X4965 1 DigitalLDOLogic_VIA2 $T=119020 17140 0 0 $X=118550 $Y=16910
X4966 1 DigitalLDOLogic_VIA2 $T=119020 21220 0 0 $X=118550 $Y=20990
X4967 1 DigitalLDOLogic_VIA2 $T=119020 25300 0 0 $X=118550 $Y=25070
X4968 1 DigitalLDOLogic_VIA2 $T=119020 29380 0 0 $X=118550 $Y=29150
X4969 1 DigitalLDOLogic_VIA2 $T=119020 33460 0 0 $X=118550 $Y=33230
X4970 1 DigitalLDOLogic_VIA2 $T=119020 37540 0 0 $X=118550 $Y=37310
X4971 1 DigitalLDOLogic_VIA2 $T=119020 41620 0 0 $X=118550 $Y=41390
X4972 1 DigitalLDOLogic_VIA2 $T=119020 45700 0 0 $X=118550 $Y=45470
X4973 1 DigitalLDOLogic_VIA2 $T=119020 49780 0 0 $X=118550 $Y=49550
X4974 1 DigitalLDOLogic_VIA2 $T=119020 53860 0 0 $X=118550 $Y=53630
X4975 1 DigitalLDOLogic_VIA2 $T=119020 57940 0 0 $X=118550 $Y=57710
X4976 3 DigitalLDOLogic_VIA2 $T=122700 11700 0 0 $X=122230 $Y=11470
X4977 3 DigitalLDOLogic_VIA2 $T=122700 15780 0 0 $X=122230 $Y=15550
X4978 3 DigitalLDOLogic_VIA2 $T=122700 19860 0 0 $X=122230 $Y=19630
X4979 3 DigitalLDOLogic_VIA2 $T=122700 23940 0 0 $X=122230 $Y=23710
X4980 3 DigitalLDOLogic_VIA2 $T=122700 28020 0 0 $X=122230 $Y=27790
X4981 3 DigitalLDOLogic_VIA2 $T=122700 32100 0 0 $X=122230 $Y=31870
X4982 3 DigitalLDOLogic_VIA2 $T=122700 36180 0 0 $X=122230 $Y=35950
X4983 3 DigitalLDOLogic_VIA2 $T=122700 40260 0 0 $X=122230 $Y=40030
X4984 3 DigitalLDOLogic_VIA2 $T=122700 44340 0 0 $X=122230 $Y=44110
X4985 3 DigitalLDOLogic_VIA2 $T=122700 48420 0 0 $X=122230 $Y=48190
X4986 3 DigitalLDOLogic_VIA2 $T=122700 52500 0 0 $X=122230 $Y=52270
X4987 3 DigitalLDOLogic_VIA2 $T=122700 56580 0 0 $X=122230 $Y=56350
X4988 1 DigitalLDOLogic_VIA2 $T=124540 13060 0 0 $X=124070 $Y=12830
X4989 1 DigitalLDOLogic_VIA2 $T=124540 17140 0 0 $X=124070 $Y=16910
X4990 1 DigitalLDOLogic_VIA2 $T=124540 21220 0 0 $X=124070 $Y=20990
X4991 1 DigitalLDOLogic_VIA2 $T=124540 25300 0 0 $X=124070 $Y=25070
X4992 1 DigitalLDOLogic_VIA2 $T=124540 29380 0 0 $X=124070 $Y=29150
X4993 1 DigitalLDOLogic_VIA2 $T=124540 33460 0 0 $X=124070 $Y=33230
X4994 1 DigitalLDOLogic_VIA2 $T=124540 37540 0 0 $X=124070 $Y=37310
X4995 1 DigitalLDOLogic_VIA2 $T=124540 41620 0 0 $X=124070 $Y=41390
X4996 1 DigitalLDOLogic_VIA2 $T=124540 45700 0 0 $X=124070 $Y=45470
X4997 1 DigitalLDOLogic_VIA2 $T=124540 49780 0 0 $X=124070 $Y=49550
X4998 1 DigitalLDOLogic_VIA2 $T=124540 53860 0 0 $X=124070 $Y=53630
X4999 1 DigitalLDOLogic_VIA2 $T=124540 57940 0 0 $X=124070 $Y=57710
X5000 3 DigitalLDOLogic_VIA2 $T=128220 11700 0 0 $X=127750 $Y=11470
X5001 3 DigitalLDOLogic_VIA2 $T=128220 15780 0 0 $X=127750 $Y=15550
X5002 3 DigitalLDOLogic_VIA2 $T=128220 19860 0 0 $X=127750 $Y=19630
X5003 3 DigitalLDOLogic_VIA2 $T=128220 23940 0 0 $X=127750 $Y=23710
X5004 3 DigitalLDOLogic_VIA2 $T=128220 28020 0 0 $X=127750 $Y=27790
X5005 3 DigitalLDOLogic_VIA2 $T=128220 32100 0 0 $X=127750 $Y=31870
X5006 3 DigitalLDOLogic_VIA2 $T=128220 36180 0 0 $X=127750 $Y=35950
X5007 3 DigitalLDOLogic_VIA2 $T=128220 40260 0 0 $X=127750 $Y=40030
X5008 3 DigitalLDOLogic_VIA2 $T=128220 44340 0 0 $X=127750 $Y=44110
X5009 3 DigitalLDOLogic_VIA2 $T=128220 48420 0 0 $X=127750 $Y=48190
X5010 3 DigitalLDOLogic_VIA2 $T=128220 52500 0 0 $X=127750 $Y=52270
X5011 3 DigitalLDOLogic_VIA2 $T=128220 56580 0 0 $X=127750 $Y=56350
X5012 1 DigitalLDOLogic_VIA2 $T=130060 13060 0 0 $X=129590 $Y=12830
X5013 1 DigitalLDOLogic_VIA2 $T=130060 17140 0 0 $X=129590 $Y=16910
X5014 1 DigitalLDOLogic_VIA2 $T=130060 21220 0 0 $X=129590 $Y=20990
X5015 1 DigitalLDOLogic_VIA2 $T=130060 25300 0 0 $X=129590 $Y=25070
X5016 1 DigitalLDOLogic_VIA2 $T=130060 29380 0 0 $X=129590 $Y=29150
X5017 1 DigitalLDOLogic_VIA2 $T=130060 33460 0 0 $X=129590 $Y=33230
X5018 1 DigitalLDOLogic_VIA2 $T=130060 37540 0 0 $X=129590 $Y=37310
X5019 1 DigitalLDOLogic_VIA2 $T=130060 41620 0 0 $X=129590 $Y=41390
X5020 1 DigitalLDOLogic_VIA2 $T=130060 45700 0 0 $X=129590 $Y=45470
X5021 1 DigitalLDOLogic_VIA2 $T=130060 49780 0 0 $X=129590 $Y=49550
X5022 1 DigitalLDOLogic_VIA2 $T=130060 53860 0 0 $X=129590 $Y=53630
X5023 1 DigitalLDOLogic_VIA2 $T=130060 57940 0 0 $X=129590 $Y=57710
X5024 3 DigitalLDOLogic_VIA2 $T=133740 11700 0 0 $X=133270 $Y=11470
X5025 3 DigitalLDOLogic_VIA2 $T=133740 15780 0 0 $X=133270 $Y=15550
X5026 3 DigitalLDOLogic_VIA2 $T=133740 19860 0 0 $X=133270 $Y=19630
X5027 3 DigitalLDOLogic_VIA2 $T=133740 23940 0 0 $X=133270 $Y=23710
X5028 3 DigitalLDOLogic_VIA2 $T=133740 28020 0 0 $X=133270 $Y=27790
X5029 3 DigitalLDOLogic_VIA2 $T=133740 32100 0 0 $X=133270 $Y=31870
X5030 3 DigitalLDOLogic_VIA2 $T=133740 36180 0 0 $X=133270 $Y=35950
X5031 3 DigitalLDOLogic_VIA2 $T=133740 40260 0 0 $X=133270 $Y=40030
X5032 3 DigitalLDOLogic_VIA2 $T=133740 44340 0 0 $X=133270 $Y=44110
X5033 3 DigitalLDOLogic_VIA2 $T=133740 48420 0 0 $X=133270 $Y=48190
X5034 3 DigitalLDOLogic_VIA2 $T=133740 52500 0 0 $X=133270 $Y=52270
X5035 3 DigitalLDOLogic_VIA2 $T=133740 56580 0 0 $X=133270 $Y=56350
X5036 1 DigitalLDOLogic_VIA2 $T=135580 13060 0 0 $X=135110 $Y=12830
X5037 1 DigitalLDOLogic_VIA2 $T=135580 17140 0 0 $X=135110 $Y=16910
X5038 1 DigitalLDOLogic_VIA2 $T=135580 21220 0 0 $X=135110 $Y=20990
X5039 1 DigitalLDOLogic_VIA2 $T=135580 25300 0 0 $X=135110 $Y=25070
X5040 1 DigitalLDOLogic_VIA2 $T=135580 29380 0 0 $X=135110 $Y=29150
X5041 1 DigitalLDOLogic_VIA2 $T=135580 33460 0 0 $X=135110 $Y=33230
X5042 1 DigitalLDOLogic_VIA2 $T=135580 37540 0 0 $X=135110 $Y=37310
X5043 1 DigitalLDOLogic_VIA2 $T=135580 41620 0 0 $X=135110 $Y=41390
X5044 1 DigitalLDOLogic_VIA2 $T=135580 45700 0 0 $X=135110 $Y=45470
X5045 1 DigitalLDOLogic_VIA2 $T=135580 49780 0 0 $X=135110 $Y=49550
X5046 1 DigitalLDOLogic_VIA2 $T=135580 53860 0 0 $X=135110 $Y=53630
X5047 1 DigitalLDOLogic_VIA2 $T=135580 57940 0 0 $X=135110 $Y=57710
X5048 3 DigitalLDOLogic_VIA2 $T=139260 11700 0 0 $X=138790 $Y=11470
X5049 3 DigitalLDOLogic_VIA2 $T=139260 15780 0 0 $X=138790 $Y=15550
X5050 3 DigitalLDOLogic_VIA2 $T=139260 19860 0 0 $X=138790 $Y=19630
X5051 3 DigitalLDOLogic_VIA2 $T=139260 23940 0 0 $X=138790 $Y=23710
X5052 3 DigitalLDOLogic_VIA2 $T=139260 28020 0 0 $X=138790 $Y=27790
X5053 3 DigitalLDOLogic_VIA2 $T=139260 32100 0 0 $X=138790 $Y=31870
X5054 3 DigitalLDOLogic_VIA2 $T=139260 36180 0 0 $X=138790 $Y=35950
X5055 3 DigitalLDOLogic_VIA2 $T=139260 40260 0 0 $X=138790 $Y=40030
X5056 3 DigitalLDOLogic_VIA2 $T=139260 44340 0 0 $X=138790 $Y=44110
X5057 3 DigitalLDOLogic_VIA2 $T=139260 48420 0 0 $X=138790 $Y=48190
X5058 3 DigitalLDOLogic_VIA2 $T=139260 52500 0 0 $X=138790 $Y=52270
X5059 3 DigitalLDOLogic_VIA2 $T=139260 56580 0 0 $X=138790 $Y=56350
X5060 1 DigitalLDOLogic_VIA2 $T=141100 13060 0 0 $X=140630 $Y=12830
X5061 1 DigitalLDOLogic_VIA2 $T=141100 17140 0 0 $X=140630 $Y=16910
X5062 1 DigitalLDOLogic_VIA2 $T=141100 21220 0 0 $X=140630 $Y=20990
X5063 1 DigitalLDOLogic_VIA2 $T=141100 25300 0 0 $X=140630 $Y=25070
X5064 1 DigitalLDOLogic_VIA2 $T=141100 29380 0 0 $X=140630 $Y=29150
X5065 1 DigitalLDOLogic_VIA2 $T=141100 33460 0 0 $X=140630 $Y=33230
X5066 1 DigitalLDOLogic_VIA2 $T=141100 37540 0 0 $X=140630 $Y=37310
X5067 1 DigitalLDOLogic_VIA2 $T=141100 41620 0 0 $X=140630 $Y=41390
X5068 1 DigitalLDOLogic_VIA2 $T=141100 45700 0 0 $X=140630 $Y=45470
X5069 1 DigitalLDOLogic_VIA2 $T=141100 49780 0 0 $X=140630 $Y=49550
X5070 1 DigitalLDOLogic_VIA2 $T=141100 53860 0 0 $X=140630 $Y=53630
X5071 1 DigitalLDOLogic_VIA2 $T=141100 57940 0 0 $X=140630 $Y=57710
X5072 3 DigitalLDOLogic_VIA2 $T=144780 11700 0 0 $X=144310 $Y=11470
X5073 3 DigitalLDOLogic_VIA2 $T=144780 15780 0 0 $X=144310 $Y=15550
X5074 3 DigitalLDOLogic_VIA2 $T=144780 19860 0 0 $X=144310 $Y=19630
X5075 3 DigitalLDOLogic_VIA2 $T=144780 23940 0 0 $X=144310 $Y=23710
X5076 3 DigitalLDOLogic_VIA2 $T=144780 28020 0 0 $X=144310 $Y=27790
X5077 3 DigitalLDOLogic_VIA2 $T=144780 32100 0 0 $X=144310 $Y=31870
X5078 3 DigitalLDOLogic_VIA2 $T=144780 36180 0 0 $X=144310 $Y=35950
X5079 3 DigitalLDOLogic_VIA2 $T=144780 40260 0 0 $X=144310 $Y=40030
X5080 3 DigitalLDOLogic_VIA2 $T=144780 44340 0 0 $X=144310 $Y=44110
X5081 3 DigitalLDOLogic_VIA2 $T=144780 48420 0 0 $X=144310 $Y=48190
X5082 3 DigitalLDOLogic_VIA2 $T=144780 52500 0 0 $X=144310 $Y=52270
X5083 3 DigitalLDOLogic_VIA2 $T=144780 56580 0 0 $X=144310 $Y=56350
X5084 1 DigitalLDOLogic_VIA2 $T=146620 13060 0 0 $X=146150 $Y=12830
X5085 1 DigitalLDOLogic_VIA2 $T=146620 17140 0 0 $X=146150 $Y=16910
X5086 1 DigitalLDOLogic_VIA2 $T=146620 21220 0 0 $X=146150 $Y=20990
X5087 1 DigitalLDOLogic_VIA2 $T=146620 25300 0 0 $X=146150 $Y=25070
X5088 1 DigitalLDOLogic_VIA2 $T=146620 29380 0 0 $X=146150 $Y=29150
X5089 1 DigitalLDOLogic_VIA2 $T=146620 33460 0 0 $X=146150 $Y=33230
X5090 1 DigitalLDOLogic_VIA2 $T=146620 37540 0 0 $X=146150 $Y=37310
X5091 1 DigitalLDOLogic_VIA2 $T=146620 41620 0 0 $X=146150 $Y=41390
X5092 1 DigitalLDOLogic_VIA2 $T=146620 45700 0 0 $X=146150 $Y=45470
X5093 1 DigitalLDOLogic_VIA2 $T=146620 49780 0 0 $X=146150 $Y=49550
X5094 1 DigitalLDOLogic_VIA2 $T=146620 53860 0 0 $X=146150 $Y=53630
X5095 1 DigitalLDOLogic_VIA2 $T=146620 57940 0 0 $X=146150 $Y=57710
X5096 3 DigitalLDOLogic_VIA2 $T=150300 11700 0 0 $X=149830 $Y=11470
X5097 3 DigitalLDOLogic_VIA2 $T=150300 15780 0 0 $X=149830 $Y=15550
X5098 3 DigitalLDOLogic_VIA2 $T=150300 19860 0 0 $X=149830 $Y=19630
X5099 3 DigitalLDOLogic_VIA2 $T=150300 23940 0 0 $X=149830 $Y=23710
X5100 3 DigitalLDOLogic_VIA2 $T=150300 28020 0 0 $X=149830 $Y=27790
X5101 3 DigitalLDOLogic_VIA2 $T=150300 32100 0 0 $X=149830 $Y=31870
X5102 3 DigitalLDOLogic_VIA2 $T=150300 36180 0 0 $X=149830 $Y=35950
X5103 3 DigitalLDOLogic_VIA2 $T=150300 40260 0 0 $X=149830 $Y=40030
X5104 3 DigitalLDOLogic_VIA2 $T=150300 44340 0 0 $X=149830 $Y=44110
X5105 3 DigitalLDOLogic_VIA2 $T=150300 48420 0 0 $X=149830 $Y=48190
X5106 3 DigitalLDOLogic_VIA2 $T=150300 52500 0 0 $X=149830 $Y=52270
X5107 3 DigitalLDOLogic_VIA2 $T=150300 56580 0 0 $X=149830 $Y=56350
X5108 1 DigitalLDOLogic_VIA2 $T=152140 13060 0 0 $X=151670 $Y=12830
X5109 1 DigitalLDOLogic_VIA2 $T=152140 17140 0 0 $X=151670 $Y=16910
X5110 1 DigitalLDOLogic_VIA2 $T=152140 21220 0 0 $X=151670 $Y=20990
X5111 1 DigitalLDOLogic_VIA2 $T=152140 25300 0 0 $X=151670 $Y=25070
X5112 1 DigitalLDOLogic_VIA2 $T=152140 29380 0 0 $X=151670 $Y=29150
X5113 1 DigitalLDOLogic_VIA2 $T=152140 33460 0 0 $X=151670 $Y=33230
X5114 1 DigitalLDOLogic_VIA2 $T=152140 37540 0 0 $X=151670 $Y=37310
X5115 1 DigitalLDOLogic_VIA2 $T=152140 41620 0 0 $X=151670 $Y=41390
X5116 1 DigitalLDOLogic_VIA2 $T=152140 45700 0 0 $X=151670 $Y=45470
X5117 1 DigitalLDOLogic_VIA2 $T=152140 49780 0 0 $X=151670 $Y=49550
X5118 1 DigitalLDOLogic_VIA2 $T=152140 53860 0 0 $X=151670 $Y=53630
X5119 1 DigitalLDOLogic_VIA2 $T=152140 57940 0 0 $X=151670 $Y=57710
X5120 3 DigitalLDOLogic_VIA2 $T=155820 11700 0 0 $X=155350 $Y=11470
X5121 3 DigitalLDOLogic_VIA2 $T=155820 15780 0 0 $X=155350 $Y=15550
X5122 3 DigitalLDOLogic_VIA2 $T=155820 19860 0 0 $X=155350 $Y=19630
X5123 3 DigitalLDOLogic_VIA2 $T=155820 23940 0 0 $X=155350 $Y=23710
X5124 3 DigitalLDOLogic_VIA2 $T=155820 28020 0 0 $X=155350 $Y=27790
X5125 3 DigitalLDOLogic_VIA2 $T=155820 32100 0 0 $X=155350 $Y=31870
X5126 3 DigitalLDOLogic_VIA2 $T=155820 36180 0 0 $X=155350 $Y=35950
X5127 3 DigitalLDOLogic_VIA2 $T=155820 40260 0 0 $X=155350 $Y=40030
X5128 3 DigitalLDOLogic_VIA2 $T=155820 44340 0 0 $X=155350 $Y=44110
X5129 3 DigitalLDOLogic_VIA2 $T=155820 48420 0 0 $X=155350 $Y=48190
X5130 3 DigitalLDOLogic_VIA2 $T=155820 52500 0 0 $X=155350 $Y=52270
X5131 3 DigitalLDOLogic_VIA2 $T=155820 56580 0 0 $X=155350 $Y=56350
X5132 1 DigitalLDOLogic_VIA2 $T=157660 13060 0 0 $X=157190 $Y=12830
X5133 1 DigitalLDOLogic_VIA2 $T=157660 17140 0 0 $X=157190 $Y=16910
X5134 1 DigitalLDOLogic_VIA2 $T=157660 21220 0 0 $X=157190 $Y=20990
X5135 1 DigitalLDOLogic_VIA2 $T=157660 25300 0 0 $X=157190 $Y=25070
X5136 1 DigitalLDOLogic_VIA2 $T=157660 29380 0 0 $X=157190 $Y=29150
X5137 1 DigitalLDOLogic_VIA2 $T=157660 33460 0 0 $X=157190 $Y=33230
X5138 1 DigitalLDOLogic_VIA2 $T=157660 37540 0 0 $X=157190 $Y=37310
X5139 1 DigitalLDOLogic_VIA2 $T=157660 41620 0 0 $X=157190 $Y=41390
X5140 1 DigitalLDOLogic_VIA2 $T=157660 45700 0 0 $X=157190 $Y=45470
X5141 1 DigitalLDOLogic_VIA2 $T=157660 49780 0 0 $X=157190 $Y=49550
X5142 1 DigitalLDOLogic_VIA2 $T=157660 53860 0 0 $X=157190 $Y=53630
X5143 1 DigitalLDOLogic_VIA2 $T=157660 57940 0 0 $X=157190 $Y=57710
X5144 3 DigitalLDOLogic_VIA2 $T=161340 11700 0 0 $X=160870 $Y=11470
X5145 3 DigitalLDOLogic_VIA2 $T=161340 15780 0 0 $X=160870 $Y=15550
X5146 3 DigitalLDOLogic_VIA2 $T=161340 19860 0 0 $X=160870 $Y=19630
X5147 3 DigitalLDOLogic_VIA2 $T=161340 23940 0 0 $X=160870 $Y=23710
X5148 3 DigitalLDOLogic_VIA2 $T=161340 28020 0 0 $X=160870 $Y=27790
X5149 3 DigitalLDOLogic_VIA2 $T=161340 32100 0 0 $X=160870 $Y=31870
X5150 3 DigitalLDOLogic_VIA2 $T=161340 36180 0 0 $X=160870 $Y=35950
X5151 3 DigitalLDOLogic_VIA2 $T=161340 40260 0 0 $X=160870 $Y=40030
X5152 3 DigitalLDOLogic_VIA2 $T=161340 44340 0 0 $X=160870 $Y=44110
X5153 3 DigitalLDOLogic_VIA2 $T=161340 48420 0 0 $X=160870 $Y=48190
X5154 3 DigitalLDOLogic_VIA2 $T=161340 52500 0 0 $X=160870 $Y=52270
X5155 3 DigitalLDOLogic_VIA2 $T=161340 56580 0 0 $X=160870 $Y=56350
X5156 1 DigitalLDOLogic_VIA2 $T=163180 13060 0 0 $X=162710 $Y=12830
X5157 1 DigitalLDOLogic_VIA2 $T=163180 17140 0 0 $X=162710 $Y=16910
X5158 1 DigitalLDOLogic_VIA2 $T=163180 21220 0 0 $X=162710 $Y=20990
X5159 1 DigitalLDOLogic_VIA2 $T=163180 25300 0 0 $X=162710 $Y=25070
X5160 1 DigitalLDOLogic_VIA2 $T=163180 29380 0 0 $X=162710 $Y=29150
X5161 1 DigitalLDOLogic_VIA2 $T=163180 33460 0 0 $X=162710 $Y=33230
X5162 1 DigitalLDOLogic_VIA2 $T=163180 37540 0 0 $X=162710 $Y=37310
X5163 1 DigitalLDOLogic_VIA2 $T=163180 41620 0 0 $X=162710 $Y=41390
X5164 1 DigitalLDOLogic_VIA2 $T=163180 45700 0 0 $X=162710 $Y=45470
X5165 1 DigitalLDOLogic_VIA2 $T=163180 49780 0 0 $X=162710 $Y=49550
X5166 1 DigitalLDOLogic_VIA2 $T=163180 53860 0 0 $X=162710 $Y=53630
X5167 1 DigitalLDOLogic_VIA2 $T=163180 57940 0 0 $X=162710 $Y=57710
X5168 3 DigitalLDOLogic_VIA2 $T=166860 11700 0 0 $X=166390 $Y=11470
X5169 3 DigitalLDOLogic_VIA2 $T=166860 15780 0 0 $X=166390 $Y=15550
X5170 3 DigitalLDOLogic_VIA2 $T=166860 19860 0 0 $X=166390 $Y=19630
X5171 3 DigitalLDOLogic_VIA2 $T=166860 23940 0 0 $X=166390 $Y=23710
X5172 3 DigitalLDOLogic_VIA2 $T=166860 28020 0 0 $X=166390 $Y=27790
X5173 3 DigitalLDOLogic_VIA2 $T=166860 32100 0 0 $X=166390 $Y=31870
X5174 3 DigitalLDOLogic_VIA2 $T=166860 36180 0 0 $X=166390 $Y=35950
X5175 3 DigitalLDOLogic_VIA2 $T=166860 40260 0 0 $X=166390 $Y=40030
X5176 3 DigitalLDOLogic_VIA2 $T=166860 44340 0 0 $X=166390 $Y=44110
X5177 3 DigitalLDOLogic_VIA2 $T=166860 48420 0 0 $X=166390 $Y=48190
X5178 3 DigitalLDOLogic_VIA2 $T=166860 52500 0 0 $X=166390 $Y=52270
X5179 3 DigitalLDOLogic_VIA2 $T=166860 56580 0 0 $X=166390 $Y=56350
X5180 1 DigitalLDOLogic_VIA2 $T=168700 13060 0 0 $X=168230 $Y=12830
X5181 1 DigitalLDOLogic_VIA2 $T=168700 17140 0 0 $X=168230 $Y=16910
X5182 1 DigitalLDOLogic_VIA2 $T=168700 21220 0 0 $X=168230 $Y=20990
X5183 1 DigitalLDOLogic_VIA2 $T=168700 25300 0 0 $X=168230 $Y=25070
X5184 1 DigitalLDOLogic_VIA2 $T=168700 29380 0 0 $X=168230 $Y=29150
X5185 1 DigitalLDOLogic_VIA2 $T=168700 33460 0 0 $X=168230 $Y=33230
X5186 1 DigitalLDOLogic_VIA2 $T=168700 37540 0 0 $X=168230 $Y=37310
X5187 1 DigitalLDOLogic_VIA2 $T=168700 41620 0 0 $X=168230 $Y=41390
X5188 1 DigitalLDOLogic_VIA2 $T=168700 45700 0 0 $X=168230 $Y=45470
X5189 1 DigitalLDOLogic_VIA2 $T=168700 49780 0 0 $X=168230 $Y=49550
X5190 1 DigitalLDOLogic_VIA2 $T=168700 53860 0 0 $X=168230 $Y=53630
X5191 1 DigitalLDOLogic_VIA2 $T=168700 57940 0 0 $X=168230 $Y=57710
X5192 3 DigitalLDOLogic_VIA2 $T=172380 11700 0 0 $X=171910 $Y=11470
X5193 3 DigitalLDOLogic_VIA2 $T=172380 15780 0 0 $X=171910 $Y=15550
X5194 3 DigitalLDOLogic_VIA2 $T=172380 19860 0 0 $X=171910 $Y=19630
X5195 3 DigitalLDOLogic_VIA2 $T=172380 23940 0 0 $X=171910 $Y=23710
X5196 3 DigitalLDOLogic_VIA2 $T=172380 28020 0 0 $X=171910 $Y=27790
X5197 3 DigitalLDOLogic_VIA2 $T=172380 32100 0 0 $X=171910 $Y=31870
X5198 3 DigitalLDOLogic_VIA2 $T=172380 36180 0 0 $X=171910 $Y=35950
X5199 3 DigitalLDOLogic_VIA2 $T=172380 40260 0 0 $X=171910 $Y=40030
X5200 3 DigitalLDOLogic_VIA2 $T=172380 44340 0 0 $X=171910 $Y=44110
X5201 3 DigitalLDOLogic_VIA2 $T=172380 48420 0 0 $X=171910 $Y=48190
X5202 3 DigitalLDOLogic_VIA2 $T=172380 52500 0 0 $X=171910 $Y=52270
X5203 3 DigitalLDOLogic_VIA2 $T=172380 56580 0 0 $X=171910 $Y=56350
X5204 1 DigitalLDOLogic_VIA2 $T=174220 13060 0 0 $X=173750 $Y=12830
X5205 1 DigitalLDOLogic_VIA2 $T=174220 17140 0 0 $X=173750 $Y=16910
X5206 1 DigitalLDOLogic_VIA2 $T=174220 21220 0 0 $X=173750 $Y=20990
X5207 1 DigitalLDOLogic_VIA2 $T=174220 25300 0 0 $X=173750 $Y=25070
X5208 1 DigitalLDOLogic_VIA2 $T=174220 29380 0 0 $X=173750 $Y=29150
X5209 1 DigitalLDOLogic_VIA2 $T=174220 33460 0 0 $X=173750 $Y=33230
X5210 1 DigitalLDOLogic_VIA2 $T=174220 37540 0 0 $X=173750 $Y=37310
X5211 1 DigitalLDOLogic_VIA2 $T=174220 41620 0 0 $X=173750 $Y=41390
X5212 1 DigitalLDOLogic_VIA2 $T=174220 45700 0 0 $X=173750 $Y=45470
X5213 1 DigitalLDOLogic_VIA2 $T=174220 49780 0 0 $X=173750 $Y=49550
X5214 1 DigitalLDOLogic_VIA2 $T=174220 53860 0 0 $X=173750 $Y=53630
X5215 1 DigitalLDOLogic_VIA2 $T=174220 57940 0 0 $X=173750 $Y=57710
X5216 3 DigitalLDOLogic_VIA2 $T=177900 11700 0 0 $X=177430 $Y=11470
X5217 3 DigitalLDOLogic_VIA2 $T=177900 15780 0 0 $X=177430 $Y=15550
X5218 3 DigitalLDOLogic_VIA2 $T=177900 19860 0 0 $X=177430 $Y=19630
X5219 3 DigitalLDOLogic_VIA2 $T=177900 23940 0 0 $X=177430 $Y=23710
X5220 3 DigitalLDOLogic_VIA2 $T=177900 28020 0 0 $X=177430 $Y=27790
X5221 3 DigitalLDOLogic_VIA2 $T=177900 32100 0 0 $X=177430 $Y=31870
X5222 3 DigitalLDOLogic_VIA2 $T=177900 36180 0 0 $X=177430 $Y=35950
X5223 3 DigitalLDOLogic_VIA2 $T=177900 40260 0 0 $X=177430 $Y=40030
X5224 3 DigitalLDOLogic_VIA2 $T=177900 44340 0 0 $X=177430 $Y=44110
X5225 3 DigitalLDOLogic_VIA2 $T=177900 48420 0 0 $X=177430 $Y=48190
X5226 3 DigitalLDOLogic_VIA2 $T=177900 52500 0 0 $X=177430 $Y=52270
X5227 3 DigitalLDOLogic_VIA2 $T=177900 56580 0 0 $X=177430 $Y=56350
X5228 1 DigitalLDOLogic_VIA2 $T=179740 13060 0 0 $X=179270 $Y=12830
X5229 1 DigitalLDOLogic_VIA2 $T=179740 17140 0 0 $X=179270 $Y=16910
X5230 1 DigitalLDOLogic_VIA2 $T=179740 21220 0 0 $X=179270 $Y=20990
X5231 1 DigitalLDOLogic_VIA2 $T=179740 25300 0 0 $X=179270 $Y=25070
X5232 1 DigitalLDOLogic_VIA2 $T=179740 29380 0 0 $X=179270 $Y=29150
X5233 1 DigitalLDOLogic_VIA2 $T=179740 33460 0 0 $X=179270 $Y=33230
X5234 1 DigitalLDOLogic_VIA2 $T=179740 37540 0 0 $X=179270 $Y=37310
X5235 1 DigitalLDOLogic_VIA2 $T=179740 41620 0 0 $X=179270 $Y=41390
X5236 1 DigitalLDOLogic_VIA2 $T=179740 45700 0 0 $X=179270 $Y=45470
X5237 1 DigitalLDOLogic_VIA2 $T=179740 49780 0 0 $X=179270 $Y=49550
X5238 1 DigitalLDOLogic_VIA2 $T=179740 53860 0 0 $X=179270 $Y=53630
X5239 1 DigitalLDOLogic_VIA2 $T=179740 57940 0 0 $X=179270 $Y=57710
X5240 3 DigitalLDOLogic_VIA2 $T=183420 11700 0 0 $X=182950 $Y=11470
X5241 3 DigitalLDOLogic_VIA2 $T=183420 15780 0 0 $X=182950 $Y=15550
X5242 3 DigitalLDOLogic_VIA2 $T=183420 19860 0 0 $X=182950 $Y=19630
X5243 3 DigitalLDOLogic_VIA2 $T=183420 23940 0 0 $X=182950 $Y=23710
X5244 3 DigitalLDOLogic_VIA2 $T=183420 28020 0 0 $X=182950 $Y=27790
X5245 3 DigitalLDOLogic_VIA2 $T=183420 32100 0 0 $X=182950 $Y=31870
X5246 3 DigitalLDOLogic_VIA2 $T=183420 36180 0 0 $X=182950 $Y=35950
X5247 3 DigitalLDOLogic_VIA2 $T=183420 40260 0 0 $X=182950 $Y=40030
X5248 3 DigitalLDOLogic_VIA2 $T=183420 44340 0 0 $X=182950 $Y=44110
X5249 3 DigitalLDOLogic_VIA2 $T=183420 48420 0 0 $X=182950 $Y=48190
X5250 3 DigitalLDOLogic_VIA2 $T=183420 52500 0 0 $X=182950 $Y=52270
X5251 3 DigitalLDOLogic_VIA2 $T=183420 56580 0 0 $X=182950 $Y=56350
X5252 1 DigitalLDOLogic_VIA2 $T=185260 13060 0 0 $X=184790 $Y=12830
X5253 1 DigitalLDOLogic_VIA2 $T=185260 17140 0 0 $X=184790 $Y=16910
X5254 1 DigitalLDOLogic_VIA2 $T=185260 21220 0 0 $X=184790 $Y=20990
X5255 1 DigitalLDOLogic_VIA2 $T=185260 25300 0 0 $X=184790 $Y=25070
X5256 1 DigitalLDOLogic_VIA2 $T=185260 29380 0 0 $X=184790 $Y=29150
X5257 1 DigitalLDOLogic_VIA2 $T=185260 33460 0 0 $X=184790 $Y=33230
X5258 1 DigitalLDOLogic_VIA2 $T=185260 37540 0 0 $X=184790 $Y=37310
X5259 1 DigitalLDOLogic_VIA2 $T=185260 41620 0 0 $X=184790 $Y=41390
X5260 1 DigitalLDOLogic_VIA2 $T=185260 45700 0 0 $X=184790 $Y=45470
X5261 1 DigitalLDOLogic_VIA2 $T=185260 49780 0 0 $X=184790 $Y=49550
X5262 1 DigitalLDOLogic_VIA2 $T=185260 53860 0 0 $X=184790 $Y=53630
X5263 1 DigitalLDOLogic_VIA2 $T=185260 57940 0 0 $X=184790 $Y=57710
X5264 3 DigitalLDOLogic_VIA2 $T=188940 11700 0 0 $X=188470 $Y=11470
X5265 3 DigitalLDOLogic_VIA2 $T=188940 15780 0 0 $X=188470 $Y=15550
X5266 3 DigitalLDOLogic_VIA2 $T=188940 19860 0 0 $X=188470 $Y=19630
X5267 3 DigitalLDOLogic_VIA2 $T=188940 23940 0 0 $X=188470 $Y=23710
X5268 3 DigitalLDOLogic_VIA2 $T=188940 28020 0 0 $X=188470 $Y=27790
X5269 3 DigitalLDOLogic_VIA2 $T=188940 32100 0 0 $X=188470 $Y=31870
X5270 3 DigitalLDOLogic_VIA2 $T=188940 36180 0 0 $X=188470 $Y=35950
X5271 3 DigitalLDOLogic_VIA2 $T=188940 40260 0 0 $X=188470 $Y=40030
X5272 3 DigitalLDOLogic_VIA2 $T=188940 44340 0 0 $X=188470 $Y=44110
X5273 3 DigitalLDOLogic_VIA2 $T=188940 48420 0 0 $X=188470 $Y=48190
X5274 3 DigitalLDOLogic_VIA2 $T=188940 52500 0 0 $X=188470 $Y=52270
X5275 3 DigitalLDOLogic_VIA2 $T=188940 56580 0 0 $X=188470 $Y=56350
X5276 3 DigitalLDOLogic_VIA3 $T=12300 18500 0 0 $X=11590 $Y=17500
X5277 3 DigitalLDOLogic_VIA3 $T=12300 38900 0 0 $X=11590 $Y=37900
X5278 3 DigitalLDOLogic_VIA3 $T=17820 18500 0 0 $X=17110 $Y=17500
X5279 3 DigitalLDOLogic_VIA3 $T=17820 38900 0 0 $X=17110 $Y=37900
X5280 3 DigitalLDOLogic_VIA3 $T=23340 18500 0 0 $X=22630 $Y=17500
X5281 3 DigitalLDOLogic_VIA3 $T=23340 38900 0 0 $X=22630 $Y=37900
X5282 3 DigitalLDOLogic_VIA3 $T=28860 18500 0 0 $X=28150 $Y=17500
X5283 3 DigitalLDOLogic_VIA3 $T=28860 38900 0 0 $X=28150 $Y=37900
X5284 3 DigitalLDOLogic_VIA3 $T=34380 18500 0 0 $X=33670 $Y=17500
X5285 3 DigitalLDOLogic_VIA3 $T=34380 38900 0 0 $X=33670 $Y=37900
X5286 3 DigitalLDOLogic_VIA3 $T=39900 18500 0 0 $X=39190 $Y=17500
X5287 3 DigitalLDOLogic_VIA3 $T=39900 38900 0 0 $X=39190 $Y=37900
X5288 3 DigitalLDOLogic_VIA3 $T=45420 18500 0 0 $X=44710 $Y=17500
X5289 3 DigitalLDOLogic_VIA3 $T=45420 38900 0 0 $X=44710 $Y=37900
X5290 3 DigitalLDOLogic_VIA3 $T=50940 18500 0 0 $X=50230 $Y=17500
X5291 3 DigitalLDOLogic_VIA3 $T=50940 38900 0 0 $X=50230 $Y=37900
X5292 3 DigitalLDOLogic_VIA3 $T=56460 18500 0 0 $X=55750 $Y=17500
X5293 3 DigitalLDOLogic_VIA3 $T=56460 38900 0 0 $X=55750 $Y=37900
X5294 3 DigitalLDOLogic_VIA3 $T=61980 18500 0 0 $X=61270 $Y=17500
X5295 3 DigitalLDOLogic_VIA3 $T=61980 38900 0 0 $X=61270 $Y=37900
X5296 3 DigitalLDOLogic_VIA3 $T=67500 18500 0 0 $X=66790 $Y=17500
X5297 3 DigitalLDOLogic_VIA3 $T=67500 38900 0 0 $X=66790 $Y=37900
X5298 3 DigitalLDOLogic_VIA3 $T=73020 18500 0 0 $X=72310 $Y=17500
X5299 3 DigitalLDOLogic_VIA3 $T=73020 38900 0 0 $X=72310 $Y=37900
X5300 3 DigitalLDOLogic_VIA3 $T=78540 18500 0 0 $X=77830 $Y=17500
X5301 3 DigitalLDOLogic_VIA3 $T=78540 38900 0 0 $X=77830 $Y=37900
X5302 3 DigitalLDOLogic_VIA3 $T=84060 18500 0 0 $X=83350 $Y=17500
X5303 3 DigitalLDOLogic_VIA3 $T=84060 38900 0 0 $X=83350 $Y=37900
X5304 3 DigitalLDOLogic_VIA3 $T=89580 18500 0 0 $X=88870 $Y=17500
X5305 3 DigitalLDOLogic_VIA3 $T=89580 38900 0 0 $X=88870 $Y=37900
X5306 3 DigitalLDOLogic_VIA3 $T=95100 18500 0 0 $X=94390 $Y=17500
X5307 3 DigitalLDOLogic_VIA3 $T=95100 38900 0 0 $X=94390 $Y=37900
X5308 3 DigitalLDOLogic_VIA3 $T=100620 18500 0 0 $X=99910 $Y=17500
X5309 3 DigitalLDOLogic_VIA3 $T=100620 38900 0 0 $X=99910 $Y=37900
X5310 3 DigitalLDOLogic_VIA3 $T=106140 18500 0 0 $X=105430 $Y=17500
X5311 3 DigitalLDOLogic_VIA3 $T=106140 38900 0 0 $X=105430 $Y=37900
X5312 3 DigitalLDOLogic_VIA3 $T=111660 18500 0 0 $X=110950 $Y=17500
X5313 3 DigitalLDOLogic_VIA3 $T=111660 38900 0 0 $X=110950 $Y=37900
X5314 3 DigitalLDOLogic_VIA3 $T=117180 18500 0 0 $X=116470 $Y=17500
X5315 3 DigitalLDOLogic_VIA3 $T=117180 38900 0 0 $X=116470 $Y=37900
X5316 3 DigitalLDOLogic_VIA3 $T=122700 18500 0 0 $X=121990 $Y=17500
X5317 3 DigitalLDOLogic_VIA3 $T=122700 38900 0 0 $X=121990 $Y=37900
X5318 3 DigitalLDOLogic_VIA3 $T=128220 18500 0 0 $X=127510 $Y=17500
X5319 3 DigitalLDOLogic_VIA3 $T=128220 38900 0 0 $X=127510 $Y=37900
X5320 3 DigitalLDOLogic_VIA3 $T=133740 18500 0 0 $X=133030 $Y=17500
X5321 3 DigitalLDOLogic_VIA3 $T=133740 38900 0 0 $X=133030 $Y=37900
X5322 3 DigitalLDOLogic_VIA3 $T=139260 18500 0 0 $X=138550 $Y=17500
X5323 3 DigitalLDOLogic_VIA3 $T=139260 38900 0 0 $X=138550 $Y=37900
X5324 3 DigitalLDOLogic_VIA3 $T=144780 18500 0 0 $X=144070 $Y=17500
X5325 3 DigitalLDOLogic_VIA3 $T=144780 38900 0 0 $X=144070 $Y=37900
X5326 3 DigitalLDOLogic_VIA3 $T=150300 18500 0 0 $X=149590 $Y=17500
X5327 3 DigitalLDOLogic_VIA3 $T=150300 38900 0 0 $X=149590 $Y=37900
X5328 3 DigitalLDOLogic_VIA3 $T=155820 18500 0 0 $X=155110 $Y=17500
X5329 3 DigitalLDOLogic_VIA3 $T=155820 38900 0 0 $X=155110 $Y=37900
X5330 3 DigitalLDOLogic_VIA3 $T=161340 18500 0 0 $X=160630 $Y=17500
X5331 3 DigitalLDOLogic_VIA3 $T=161340 38900 0 0 $X=160630 $Y=37900
X5332 3 DigitalLDOLogic_VIA3 $T=166860 18500 0 0 $X=166150 $Y=17500
X5333 3 DigitalLDOLogic_VIA3 $T=166860 38900 0 0 $X=166150 $Y=37900
X5334 3 DigitalLDOLogic_VIA3 $T=172380 18500 0 0 $X=171670 $Y=17500
X5335 3 DigitalLDOLogic_VIA3 $T=172380 38900 0 0 $X=171670 $Y=37900
X5336 3 DigitalLDOLogic_VIA3 $T=177900 18500 0 0 $X=177190 $Y=17500
X5337 3 DigitalLDOLogic_VIA3 $T=177900 38900 0 0 $X=177190 $Y=37900
X5338 3 DigitalLDOLogic_VIA3 $T=183420 18500 0 0 $X=182710 $Y=17500
X5339 3 DigitalLDOLogic_VIA3 $T=183420 38900 0 0 $X=182710 $Y=37900
X5340 3 DigitalLDOLogic_VIA3 $T=188940 18500 0 0 $X=188230 $Y=17500
X5341 3 DigitalLDOLogic_VIA3 $T=188940 38900 0 0 $X=188230 $Y=37900
X5342 1 DigitalLDOLogic_VIA4 $T=12070 10110 0 0 $X=11820 $Y=9980
X5343 1 DigitalLDOLogic_VIA4 $T=14830 10110 0 0 $X=14580 $Y=9980
X5344 1 DigitalLDOLogic_VIA4 $T=17590 10110 0 0 $X=17340 $Y=9980
X5345 1 DigitalLDOLogic_VIA4 $T=20350 10110 0 0 $X=20100 $Y=9980
X5346 1 DigitalLDOLogic_VIA4 $T=23110 10110 0 0 $X=22860 $Y=9980
X5347 1 DigitalLDOLogic_VIA4 $T=25870 10110 0 0 $X=25620 $Y=9980
X5348 1 DigitalLDOLogic_VIA4 $T=28630 10110 0 0 $X=28380 $Y=9980
X5349 1 DigitalLDOLogic_VIA4 $T=31390 10110 0 0 $X=31140 $Y=9980
X5350 1 DigitalLDOLogic_VIA4 $T=34150 10110 0 0 $X=33900 $Y=9980
X5351 1 DigitalLDOLogic_VIA4 $T=36910 10110 0 0 $X=36660 $Y=9980
X5352 1 DigitalLDOLogic_VIA4 $T=39670 10110 0 0 $X=39420 $Y=9980
X5353 1 DigitalLDOLogic_VIA4 $T=42430 10110 0 0 $X=42180 $Y=9980
X5354 1 DigitalLDOLogic_VIA4 $T=45190 10110 0 0 $X=44940 $Y=9980
X5355 1 DigitalLDOLogic_VIA4 $T=47950 10110 0 0 $X=47700 $Y=9980
X5356 1 DigitalLDOLogic_VIA4 $T=50710 10110 0 0 $X=50460 $Y=9980
X5357 1 DigitalLDOLogic_VIA4 $T=53470 10110 0 0 $X=53220 $Y=9980
X5358 1 DigitalLDOLogic_VIA4 $T=56230 10110 0 0 $X=55980 $Y=9980
X5359 1 DigitalLDOLogic_VIA4 $T=58990 10110 0 0 $X=58740 $Y=9980
X5360 1 DigitalLDOLogic_VIA4 $T=61750 10110 0 0 $X=61500 $Y=9980
X5361 1 DigitalLDOLogic_VIA4 $T=64510 10110 0 0 $X=64260 $Y=9980
X5362 1 DigitalLDOLogic_VIA4 $T=67270 10110 0 0 $X=67020 $Y=9980
X5363 1 DigitalLDOLogic_VIA4 $T=70030 10110 0 0 $X=69780 $Y=9980
X5364 1 DigitalLDOLogic_VIA4 $T=72790 10110 0 0 $X=72540 $Y=9980
X5365 1 DigitalLDOLogic_VIA4 $T=75550 10110 0 0 $X=75300 $Y=9980
X5366 1 DigitalLDOLogic_VIA4 $T=78310 10110 0 0 $X=78060 $Y=9980
X5367 1 DigitalLDOLogic_VIA4 $T=81070 10110 0 0 $X=80820 $Y=9980
X5368 1 DigitalLDOLogic_VIA4 $T=83830 10110 0 0 $X=83580 $Y=9980
X5369 1 DigitalLDOLogic_VIA4 $T=86590 10110 0 0 $X=86340 $Y=9980
X5370 1 DigitalLDOLogic_VIA4 $T=89350 10110 0 0 $X=89100 $Y=9980
X5371 1 DigitalLDOLogic_VIA4 $T=92110 10110 0 0 $X=91860 $Y=9980
X5372 1 DigitalLDOLogic_VIA4 $T=94870 10110 0 0 $X=94620 $Y=9980
X5373 1 DigitalLDOLogic_VIA4 $T=97630 10110 0 0 $X=97380 $Y=9980
X5374 1 DigitalLDOLogic_VIA4 $T=100390 10110 0 0 $X=100140 $Y=9980
X5375 1 DigitalLDOLogic_VIA4 $T=103150 10110 0 0 $X=102900 $Y=9980
X5376 1 DigitalLDOLogic_VIA4 $T=105910 10110 0 0 $X=105660 $Y=9980
X5377 1 DigitalLDOLogic_VIA4 $T=108670 10110 0 0 $X=108420 $Y=9980
X5378 1 DigitalLDOLogic_VIA4 $T=111430 10110 0 0 $X=111180 $Y=9980
X5379 1 DigitalLDOLogic_VIA4 $T=114190 10110 0 0 $X=113940 $Y=9980
X5380 1 DigitalLDOLogic_VIA4 $T=116950 10110 0 0 $X=116700 $Y=9980
X5381 1 DigitalLDOLogic_VIA4 $T=119710 10110 0 0 $X=119460 $Y=9980
X5382 1 DigitalLDOLogic_VIA4 $T=122470 10110 0 0 $X=122220 $Y=9980
X5383 1 DigitalLDOLogic_VIA4 $T=125230 10110 0 0 $X=124980 $Y=9980
X5384 1 DigitalLDOLogic_VIA4 $T=127990 10110 0 0 $X=127740 $Y=9980
X5385 1 DigitalLDOLogic_VIA4 $T=130750 10110 0 0 $X=130500 $Y=9980
X5386 1 DigitalLDOLogic_VIA4 $T=133510 10110 0 0 $X=133260 $Y=9980
X5387 1 DigitalLDOLogic_VIA4 $T=136270 10110 0 0 $X=136020 $Y=9980
X5388 1 DigitalLDOLogic_VIA4 $T=139030 10110 0 0 $X=138780 $Y=9980
X5389 1 DigitalLDOLogic_VIA4 $T=141790 10110 0 0 $X=141540 $Y=9980
X5390 1 DigitalLDOLogic_VIA4 $T=144550 10110 0 0 $X=144300 $Y=9980
X5391 1 DigitalLDOLogic_VIA4 $T=147310 10110 0 0 $X=147060 $Y=9980
X5392 1 DigitalLDOLogic_VIA4 $T=150070 10110 0 0 $X=149820 $Y=9980
X5393 1 DigitalLDOLogic_VIA4 $T=152830 10110 0 0 $X=152580 $Y=9980
X5394 1 DigitalLDOLogic_VIA4 $T=155590 10110 0 0 $X=155340 $Y=9980
X5395 1 DigitalLDOLogic_VIA4 $T=158350 10110 0 0 $X=158100 $Y=9980
X5396 1 DigitalLDOLogic_VIA4 $T=161110 10110 0 0 $X=160860 $Y=9980
X5397 1 DigitalLDOLogic_VIA4 $T=163870 10110 0 0 $X=163620 $Y=9980
X5398 1 DigitalLDOLogic_VIA4 $T=166630 10110 0 0 $X=166380 $Y=9980
X5399 1 DigitalLDOLogic_VIA4 $T=169390 10110 0 0 $X=169140 $Y=9980
X5400 1 DigitalLDOLogic_VIA4 $T=172150 10110 0 0 $X=171900 $Y=9980
X5401 1 DigitalLDOLogic_VIA4 $T=174910 10110 0 0 $X=174660 $Y=9980
X5402 1 DigitalLDOLogic_VIA4 $T=177670 10110 0 0 $X=177420 $Y=9980
X5403 1 DigitalLDOLogic_VIA4 $T=180430 10110 0 0 $X=180180 $Y=9980
X5404 1 DigitalLDOLogic_VIA4 $T=183190 10110 0 0 $X=182940 $Y=9980
X5405 1 DigitalLDOLogic_VIA4 $T=185950 10110 0 0 $X=185700 $Y=9980
X5406 1 DigitalLDOLogic_VIA4 $T=188710 10110 0 0 $X=188460 $Y=9980
X5407 1 3 MASCO__Y1 $T=13430 24300 0 0 $X=13430 $Y=24300
X5408 1 3 MASCO__Y1 $T=13430 44700 0 0 $X=13430 $Y=44700
X5409 1 3 MASCO__Y1 $T=57590 24300 0 0 $X=57590 $Y=24300
X5410 1 3 MASCO__Y1 $T=57590 44700 0 0 $X=57590 $Y=44700
X5411 1 3 MASCO__Y1 $T=101750 24300 0 0 $X=101750 $Y=24300
X5412 1 3 MASCO__Y1 $T=101750 44700 0 0 $X=101750 $Y=44700
X5413 1 3 MASCO__Y1 $T=145910 24300 0 0 $X=145910 $Y=24300
X5414 1 3 MASCO__Y1 $T=145910 44700 0 0 $X=145910 $Y=44700
X5415 1 3 MASCO__B19 $T=29130 26080 0 0 $X=29130 $Y=26080
X5416 1 3 MASCO__B19 $T=29130 31520 0 0 $X=29130 $Y=31520
X5417 1 3 MASCO__B19 $T=29130 36960 0 0 $X=29130 $Y=36960
X5418 1 3 MASCO__B19 $T=29130 42400 0 0 $X=29130 $Y=42400
X5419 1 3 MASCO__B19 $T=29130 47840 0 0 $X=29130 $Y=47840
X5420 1 3 MASCO__B19 $T=29130 53280 0 0 $X=29130 $Y=53280
X5421 1 3 MASCO__B19 $T=58570 31520 0 0 $X=58570 $Y=31520
X5422 1 3 MASCO__B19 $T=58570 36960 0 0 $X=58570 $Y=36960
X5423 1 3 MASCO__B19 $T=58570 42400 0 0 $X=58570 $Y=42400
X5424 1 3 MASCO__B19 $T=58570 47840 0 0 $X=58570 $Y=47840
X5425 1 3 MASCO__B19 $T=58570 53280 0 0 $X=58570 $Y=53280
X5426 1 3 MASCO__B19 $T=88010 31520 0 0 $X=88010 $Y=31520
X5427 1 3 MASCO__B19 $T=88010 36960 0 0 $X=88010 $Y=36960
X5428 1 3 MASCO__B19 $T=88010 42400 0 0 $X=88010 $Y=42400
X5429 1 3 MASCO__B19 $T=88010 47840 0 0 $X=88010 $Y=47840
X5430 1 3 MASCO__B19 $T=88010 53280 0 0 $X=88010 $Y=53280
X5431 1 3 MASCO__B19 $T=102730 20640 0 0 $X=102730 $Y=20640
X5432 1 3 MASCO__B19 $T=146890 26080 0 0 $X=146890 $Y=26080
X5433 1 3 MASCO__B19 $T=176330 9760 0 0 $X=176330 $Y=9760
X5434 1 3 MASCO__B19 $T=176330 26080 0 0 $X=176330 $Y=26080
X5435 1 3 MASCO__B22 $T=25910 26080 0 0 $X=25910 $Y=26080
X5436 1 3 MASCO__B22 $T=25910 31520 0 0 $X=25910 $Y=31520
X5437 1 3 MASCO__B22 $T=25910 36960 0 0 $X=25910 $Y=36960
X5438 1 3 MASCO__B22 $T=25910 42400 0 0 $X=25910 $Y=42400
X5439 1 3 MASCO__B22 $T=25910 47840 0 0 $X=25910 $Y=47840
X5440 1 3 MASCO__B22 $T=25910 53280 0 0 $X=25910 $Y=53280
X5441 1 3 MASCO__B22 $T=84790 31520 0 0 $X=84790 $Y=31520
X5442 1 3 MASCO__B22 $T=84790 36960 0 0 $X=84790 $Y=36960
X5443 1 3 MASCO__B22 $T=84790 42400 0 0 $X=84790 $Y=42400
X5444 1 3 MASCO__B22 $T=84790 47840 0 0 $X=84790 $Y=47840
X5445 1 3 MASCO__B22 $T=84790 53280 0 0 $X=84790 $Y=53280
X5446 1 3 MASCO__B22 $T=114230 26080 0 0 $X=114230 $Y=26080
X5447 1 3 MASCO__B22 $T=114230 31520 0 0 $X=114230 $Y=31520
X5448 1 3 MASCO__B22 $T=114230 36960 0 0 $X=114230 $Y=36960
X5449 1 3 MASCO__B22 $T=114230 42400 0 0 $X=114230 $Y=42400
X5450 1 3 MASCO__B22 $T=114230 47840 0 0 $X=114230 $Y=47840
X5451 1 3 MASCO__B22 $T=114230 53280 0 0 $X=114230 $Y=53280
X5452 1 3 MASCO__B22 $T=173110 26080 0 0 $X=173110 $Y=26080
X5453 1 3 MASCO__B26 $T=13030 9760 0 0 $X=13030 $Y=9760
X5454 1 3 MASCO__B26 $T=13030 15200 0 0 $X=13030 $Y=15200
X5455 1 3 MASCO__B26 $T=13030 20640 0 0 $X=13030 $Y=20640
X5456 1 3 MASCO__B26 $T=13030 26080 0 0 $X=13030 $Y=26080
X5457 1 3 MASCO__B26 $T=13030 31520 0 0 $X=13030 $Y=31520
X5458 1 3 MASCO__B26 $T=13030 36960 0 0 $X=13030 $Y=36960
X5459 1 3 MASCO__B26 $T=13030 42400 0 0 $X=13030 $Y=42400
X5460 1 3 MASCO__B26 $T=13030 47840 0 0 $X=13030 $Y=47840
X5461 1 3 MASCO__B26 $T=13030 53280 0 0 $X=13030 $Y=53280
X5462 1 3 MASCO__B26 $T=42470 9760 0 0 $X=42470 $Y=9760
X5463 1 3 MASCO__B26 $T=42470 26080 0 0 $X=42470 $Y=26080
X5464 1 3 MASCO__B26 $T=42470 31520 0 0 $X=42470 $Y=31520
X5465 1 3 MASCO__B26 $T=42470 36960 0 0 $X=42470 $Y=36960
X5466 1 3 MASCO__B26 $T=42470 42400 0 0 $X=42470 $Y=42400
X5467 1 3 MASCO__B26 $T=42470 47840 0 0 $X=42470 $Y=47840
X5468 1 3 MASCO__B26 $T=42470 53280 0 0 $X=42470 $Y=53280
X5469 1 3 MASCO__B26 $T=71910 31520 0 0 $X=71910 $Y=31520
X5470 1 3 MASCO__B26 $T=71910 36960 0 0 $X=71910 $Y=36960
X5471 1 3 MASCO__B26 $T=71910 42400 0 0 $X=71910 $Y=42400
X5472 1 3 MASCO__B26 $T=71910 47840 0 0 $X=71910 $Y=47840
X5473 1 3 MASCO__B26 $T=71910 53280 0 0 $X=71910 $Y=53280
X5474 1 3 MASCO__B26 $T=101350 31520 0 0 $X=101350 $Y=31520
X5475 1 3 MASCO__B26 $T=101350 36960 0 0 $X=101350 $Y=36960
X5476 1 3 MASCO__B26 $T=101350 42400 0 0 $X=101350 $Y=42400
X5477 1 3 MASCO__B26 $T=101350 47840 0 0 $X=101350 $Y=47840
X5478 1 3 MASCO__B26 $T=101350 53280 0 0 $X=101350 $Y=53280
X5479 1 3 MASCO__B26 $T=130790 15200 0 0 $X=130790 $Y=15200
X5480 1 3 MASCO__B26 $T=160230 26080 0 0 $X=160230 $Y=26080
.ends DigitalLDOLogic
