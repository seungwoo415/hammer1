* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : digital_ldo_top                              *
* Netlisted  : Wed Jan 29 00:53:36 2025                     *
* Pegasus Version: 22.14-s007 Tue Jan 31 16:35:56 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 1 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)
*.DEVTMPLT 2 MP(pfet_01v8_hvt) hvtpfet_01v8_rec pSourceDrain(D) hvtpfet(G) pSourceDrain(s) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__diode_2                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__diode_2 1 2 3 4 5
** N=5 EP=5 FDC=0
.ends sky130_fd_sc_hd__diode_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__clkbuf_1                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__clkbuf_1 1 2 3 4 5 6
** N=7 EP=6 FDC=4
M0 3 7 2 5 nfet_01v8 L=1.5e-07 W=5.2e-07 $X=395 $Y=235 $dt=0
M1 7 4 3 5 nfet_01v8 L=1.5e-07 W=5.2e-07 $X=835 $Y=235 $dt=0
M2 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=7.9e-07 $X=395 $Y=1695 $dt=2
M3 7 4 1 6 pfet_01v8_hvt L=1.5e-07 W=7.9e-07 $X=835 $Y=1695 $dt=2
.ends sky130_fd_sc_hd__clkbuf_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__buf_8                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__buf_8 1 2 3 4 5 6 7
** N=8 EP=7 FDC=22
M0 3 4 8 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=395 $Y=235 $dt=0
M1 8 4 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=815 $Y=235 $dt=0
M2 3 4 8 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1235 $Y=235 $dt=0
M3 2 8 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1655 $Y=235 $dt=0
M4 3 8 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2075 $Y=235 $dt=0
M5 2 8 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2495 $Y=235 $dt=0
M6 3 8 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2915 $Y=235 $dt=0
M7 2 8 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=3335 $Y=235 $dt=0
M8 3 8 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=3755 $Y=235 $dt=0
M9 2 8 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=4175 $Y=235 $dt=0
M10 3 8 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=4595 $Y=235 $dt=0
M11 1 4 8 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=395 $Y=1485 $dt=2
M12 8 4 1 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=815 $Y=1485 $dt=2
M13 1 4 8 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1235 $Y=1485 $dt=2
M14 2 8 1 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1655 $Y=1485 $dt=2
M15 1 8 2 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2075 $Y=1485 $dt=2
M16 2 8 1 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2495 $Y=1485 $dt=2
M17 1 8 2 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2915 $Y=1485 $dt=2
M18 2 8 1 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=3335 $Y=1485 $dt=2
M19 1 8 2 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=3755 $Y=1485 $dt=2
M20 2 8 1 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=4175 $Y=1485 $dt=2
M21 1 8 2 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=4595 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__buf_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__dlygate4sd2_1                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__dlygate4sd2_1 1 2 3 4 5 6
** N=9 EP=6 FDC=8
M0 3 4 7 5 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=505 $Y=235 $dt=0
M1 8 7 3 5 nfet_01v8 L=1.8e-07 W=4.2e-07 $X=925 $Y=235 $dt=0
M2 3 8 9 5 nfet_01v8 L=1.8e-07 W=4.2e-07 $X=1895 $Y=235 $dt=0
M3 2 9 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2400 $Y=235 $dt=0
M4 1 4 7 6 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=505 $Y=2065 $dt=2
M5 8 7 1 6 pfet_01v8_hvt L=1.8e-07 W=4.2e-07 $X=925 $Y=2065 $dt=2
M6 1 8 9 6 pfet_01v8_hvt L=1.8e-07 W=4.2e-07 $X=1895 $Y=2065 $dt=2
M7 2 9 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2400 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__dlygate4sd2_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__clkbuf_2                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__clkbuf_2 1 2 3 4 5 6
** N=7 EP=6 FDC=6
M0 3 4 7 5 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=400 $Y=235 $dt=0
M1 2 7 3 5 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=875 $Y=235 $dt=0
M2 3 7 2 5 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1295 $Y=235 $dt=0
M3 1 4 7 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=400 $Y=1485 $dt=2
M4 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=875 $Y=1485 $dt=2
M5 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1295 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__clkbuf_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__clkbuf_1_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__clkbuf_1_DigitalLDOLogic_gds 1 2 3 4 5 6
** N=7 EP=6 FDC=4
M0 3 7 1 5 nfet_01v8 L=1.5e-07 W=5.2e-07 $X=395 $Y=235 $dt=0
M1 7 4 3 5 nfet_01v8 L=1.5e-07 W=5.2e-07 $X=835 $Y=235 $dt=0
M2 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=7.9e-07 $X=395 $Y=1695 $dt=2
M3 7 4 2 6 pfet_01v8_hvt L=1.5e-07 W=7.9e-07 $X=835 $Y=1695 $dt=2
.ends sky130_fd_sc_hd__clkbuf_1_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds 1 2 3 4 5 6
** N=7 EP=6 FDC=22
M0 3 4 7 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=395 $Y=235 $dt=0
M1 7 4 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=815 $Y=235 $dt=0
M2 3 4 7 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1235 $Y=235 $dt=0
M3 2 7 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1655 $Y=235 $dt=0
M4 3 7 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2075 $Y=235 $dt=0
M5 2 7 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2495 $Y=235 $dt=0
M6 3 7 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2915 $Y=235 $dt=0
M7 2 7 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=3335 $Y=235 $dt=0
M8 3 7 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=3755 $Y=235 $dt=0
M9 2 7 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=4175 $Y=235 $dt=0
M10 3 7 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=4595 $Y=235 $dt=0
M11 1 4 7 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=395 $Y=1485 $dt=2
M12 7 4 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=815 $Y=1485 $dt=2
M13 1 4 7 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1235 $Y=1485 $dt=2
M14 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1655 $Y=1485 $dt=2
M15 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2075 $Y=1485 $dt=2
M16 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2495 $Y=1485 $dt=2
M17 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2915 $Y=1485 $dt=2
M18 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=3335 $Y=1485 $dt=2
M19 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=3755 $Y=1485 $dt=2
M20 2 7 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=4175 $Y=1485 $dt=2
M21 1 7 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=4595 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__dfxtp_1                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__dfxtp_1 1 2 3 4 5 6 7
** N=22 EP=7 FDC=24
M0 3 4 9 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=395 $Y=235 $dt=0
M1 8 9 3 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=815 $Y=235 $dt=0
M2 10 5 3 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1755 $Y=235 $dt=0
M3 11 9 10 6 nfet_01v8 L=1.5e-07 W=3.6e-07 $X=2315 $Y=235 $dt=0
M4 17 8 11 6 nfet_01v8 L=1.5e-07 W=3.6e-07 $X=2810 $Y=235 $dt=0
M5 3 12 17 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=3305 $Y=235 $dt=0
M6 12 11 3 6 nfet_01v8 L=1.5e-07 W=6.4e-07 $X=3900 $Y=235 $dt=0
M7 13 8 12 6 nfet_01v8 L=1.5e-07 W=3.6e-07 $X=4405 $Y=235 $dt=0
M8 18 9 13 6 nfet_01v8 L=1.5e-07 W=3.6e-07 $X=4935 $Y=235 $dt=0
M9 3 14 18 6 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=5410 $Y=235 $dt=0
M10 3 13 14 6 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=6355 $Y=235 $dt=0
M11 2 14 3 6 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=6775 $Y=235 $dt=0
M12 1 4 9 7 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=395 $Y=1815 $dt=2
M13 8 9 1 7 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=815 $Y=1815 $dt=2
M14 10 5 1 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=1755 $Y=2065 $dt=2
M15 11 8 10 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=2180 $Y=2065 $dt=2
M16 15 9 11 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=2655 $Y=2065 $dt=2
M17 1 12 15 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=3170 $Y=2065 $dt=2
M18 12 11 1 7 pfet_01v8_hvt L=1.5e-07 W=7.5e-07 $X=3830 $Y=1735 $dt=2
M19 13 9 12 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=4305 $Y=2065 $dt=2
M20 16 8 13 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=4725 $Y=2065 $dt=2
M21 1 14 16 7 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=5295 $Y=2065 $dt=2
M22 1 13 14 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=6345 $Y=1485 $dt=2
M23 2 14 1 7 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=6765 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__dfxtp_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__a221o_1                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__a221o_1 1 2 3 4 5 6 7 8 9 10
** N=17 EP=10 FDC=12
M0 3 4 13 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=395 $Y=235 $dt=0
M1 14 5 3 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=875 $Y=235 $dt=0
M2 13 6 14 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1235 $Y=235 $dt=0
M3 15 7 13 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2175 $Y=235 $dt=0
M4 3 8 15 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2655 $Y=235 $dt=0
M5 1 13 3 9 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=3120 $Y=235 $dt=0
M6 11 4 13 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=395 $Y=1485 $dt=2
M7 12 5 11 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=815 $Y=1485 $dt=2
M8 11 6 12 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1235 $Y=1485 $dt=2
M9 12 7 2 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2175 $Y=1485 $dt=2
M10 2 8 12 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2655 $Y=1485 $dt=2
M11 1 13 2 10 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=3120 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__a221o_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__a21o_1                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__a21o_1 1 2 3 4 5 6 7 8
** N=12 EP=8 FDC=8
M0 3 9 1 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=405 $Y=235 $dt=0
M1 9 4 3 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1345 $Y=235 $dt=0
M2 11 5 9 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1770 $Y=235 $dt=0
M3 3 6 11 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=2200 $Y=235 $dt=0
M4 2 9 1 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=405 $Y=1485 $dt=2
M5 10 4 9 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1345 $Y=1485 $dt=2
M6 2 5 10 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1770 $Y=1485 $dt=2
M7 10 6 2 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=2200 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__a21o_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__or3_1                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__or3_1 1 2 3 4 5 6 7 8
** N=13 EP=8 FDC=8
M0 3 4 9 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=405 $Y=265 $dt=0
M1 9 5 3 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=825 $Y=265 $dt=0
M2 3 6 9 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1245 $Y=265 $dt=0
M3 2 9 3 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=1735 $Y=235 $dt=0
M4 10 4 9 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=405 $Y=1485 $dt=2
M5 11 5 10 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=765 $Y=1485 $dt=2
M6 1 6 11 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=1245 $Y=1485 $dt=2
M7 2 9 1 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=1735 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__or3_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__inv_2                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__inv_2 1 2 3 4 5 6
** N=6 EP=6 FDC=4
M0 2 4 3 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=405 $Y=235 $dt=0
M1 3 4 2 5 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=825 $Y=235 $dt=0
M2 2 4 1 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=405 $Y=1485 $dt=2
M3 1 4 2 6 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=825 $Y=1485 $dt=2
.ends sky130_fd_sc_hd__inv_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds 1 2
** N=2 EP=2 FDC=0
.ends sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=1.97e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=1.97e-06 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=5.9e-07 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=5.9e-07 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=4.73e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=4.73e-06 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=1.05e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=1.05e-06 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=2.89e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=2.89e-06 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_PR_DigitalLDOLogic_gds                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_PR_DigitalLDOLogic_gds 1
** N=1 EP=1 FDC=0
.ends L1M1_PR_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_PR_M                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_PR_M 1
** N=1 EP=1 FDC=0
.ends M1M2_PR_M

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_PR_DigitalLDOLogic_gds                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_PR_DigitalLDOLogic_gds 1
** N=1 EP=1 FDC=0
.ends M1M2_PR_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2M3_PR_DigitalLDOLogic_gds                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2M3_PR_DigitalLDOLogic_gds 1
** N=1 EP=1 FDC=0
.ends M2M3_PR_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3M4_PR_DigitalLDOLogic_gds                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3M4_PR_DigitalLDOLogic_gds 1
** N=1 EP=1 FDC=0
.ends M3M4_PR_DigitalLDOLogic_gds

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA0                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA0 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA1                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA1 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA2                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA2 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA3                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA3 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic_VIA4                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic_VIA4 1
** N=1 EP=1 FDC=0
.ends DigitalLDOLogic_VIA4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y3 1 2
** N=2 EP=2 FDC=0
X0 1 DigitalLDOLogic_VIA3 $T=710 1000 0 0 $X=0 $Y=0
X1 1 DigitalLDOLogic_VIA3 $T=6230 1000 0 0 $X=5520 $Y=0
X2 1 DigitalLDOLogic_VIA3 $T=11750 1000 0 0 $X=11040 $Y=0
X3 1 DigitalLDOLogic_VIA3 $T=17270 1000 0 0 $X=16560 $Y=0
X4 1 DigitalLDOLogic_VIA3 $T=22790 1000 0 0 $X=22080 $Y=0
X5 1 DigitalLDOLogic_VIA3 $T=28310 1000 0 0 $X=27600 $Y=0
X6 1 DigitalLDOLogic_VIA3 $T=33830 1000 0 0 $X=33120 $Y=0
X7 1 DigitalLDOLogic_VIA3 $T=39350 1000 0 0 $X=38640 $Y=0
.ends MASCO__Y3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B94                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B94 1 2
** N=2 EP=2 FDC=4
X0 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=190 2960 1 0 $X=0 $Y=0
X1 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=190 2960 0 0 $X=0 $Y=2720
X2 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=650 2960 1 0 $X=460 $Y=0
X3 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=650 2960 0 0 $X=460 $Y=2720
.ends MASCO__B94

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B97                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B97 1 2
** N=2 EP=2 FDC=8
X0 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=2030 2960 1 0 $X=1840 $Y=0
X1 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=2030 2960 0 0 $X=1840 $Y=2720
X2 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=190 2960 1 0 $X=0 $Y=0
X3 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=190 2960 0 0 $X=0 $Y=2720
.ends MASCO__B97

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B101                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B101 1 2
** N=2 EP=2 FDC=4
X0 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=1570 2960 1 0 $X=1380 $Y=0
X1 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=1570 2960 0 0 $X=1380 $Y=2720
X2 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=190 2960 1 0 $X=0 $Y=0
X3 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=190 2960 0 0 $X=0 $Y=2720
.ends MASCO__B101

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DigitalLDOLogic                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DigitalLDOLogic 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75
** N=181 EP=75 FDC=3456
X0 1 76 2 77 2 1 sky130_fd_sc_hd__dlygate4sd2_1 $T=162260 18160 0 0 $X=162070 $Y=17920
X1 1 78 2 29 2 1 sky130_fd_sc_hd__clkbuf_2 $T=171460 23600 1 0 $X=171270 $Y=20640
X2 1 79 2 37 2 1 sky130_fd_sc_hd__clkbuf_2 $T=172840 18160 0 0 $X=172650 $Y=17920
X3 80 1 2 14 2 1 sky130_fd_sc_hd__clkbuf_1_DigitalLDOLogic_gds $T=60140 23600 1 0 $X=59950 $Y=20640
X4 81 1 2 14 2 1 sky130_fd_sc_hd__clkbuf_1_DigitalLDOLogic_gds $T=80840 23600 0 180 $X=79270 $Y=20640
X5 82 1 2 14 2 1 sky130_fd_sc_hd__clkbuf_1_DigitalLDOLogic_gds $T=134660 23600 0 180 $X=133090 $Y=20640
X6 83 1 2 14 2 1 sky130_fd_sc_hd__clkbuf_1_DigitalLDOLogic_gds $T=171460 23600 0 180 $X=169890 $Y=20640
X7 1 3 2 84 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=19200 12720 0 0 $X=19010 $Y=12480
X8 1 4 2 85 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=19200 18160 1 0 $X=19010 $Y=15200
X9 1 5 2 86 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=21040 23600 0 0 $X=20850 $Y=23360
X10 1 6 2 87 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=29780 12720 1 0 $X=29590 $Y=9760
X11 1 7 2 88 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=29780 18160 1 0 $X=29590 $Y=15200
X12 1 8 2 10 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=38060 12720 1 180 $X=32350 $Y=12480
X13 1 9 2 89 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=40820 29040 0 180 $X=35110 $Y=26080
X14 1 11 2 90 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=41280 18160 0 180 $X=35570 $Y=15200
X15 1 12 2 91 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=47720 12720 1 0 $X=47530 $Y=9760
X16 1 15 2 92 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=62440 12720 1 0 $X=62250 $Y=9760
X17 1 16 2 93 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=65660 12720 0 0 $X=65470 $Y=12480
X18 1 13 2 94 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=65660 23600 0 0 $X=65470 $Y=23360
X19 1 19 2 18 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=73940 12720 1 0 $X=73750 $Y=9760
X20 1 17 2 95 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=73940 18160 1 0 $X=73750 $Y=15200
X21 1 21 2 96 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=82680 12720 1 0 $X=82490 $Y=9760
X22 1 20 2 97 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=91420 12720 1 0 $X=91230 $Y=9760
X23 1 22 2 98 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=97400 12720 1 0 $X=97210 $Y=9760
X24 1 24 2 99 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=103380 12720 0 0 $X=103190 $Y=12480
X25 1 23 2 100 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=103380 18160 1 0 $X=103190 $Y=15200
X26 1 25 2 101 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=114880 18160 1 180 $X=109170 $Y=17920
X27 1 26 2 102 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=115800 12720 1 180 $X=110090 $Y=12480
X28 1 27 2 103 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=123620 12720 0 180 $X=117910 $Y=9760
X29 1 28 2 104 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=123620 18160 0 180 $X=117910 $Y=15200
X30 1 30 2 105 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=132820 12720 0 0 $X=132630 $Y=12480
X31 1 31 2 106 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=138340 12720 1 0 $X=138150 $Y=9760
X32 1 32 2 107 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=144780 12720 1 180 $X=139070 $Y=12480
X33 1 33 2 108 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=153060 23600 1 180 $X=147350 $Y=23360
X34 1 34 2 109 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=148460 12720 1 0 $X=148270 $Y=9760
X35 1 36 2 110 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=162260 18160 1 0 $X=162070 $Y=15200
X36 1 35 2 111 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=163180 12720 1 0 $X=162990 $Y=9760
X37 1 38 2 112 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=176980 18160 1 0 $X=176790 $Y=15200
X38 1 39 2 113 2 1 sky130_fd_sc_hd__buf_8_DigitalLDOLogic_gds $T=180200 23600 0 0 $X=180010 $Y=23360
X39 1 88 2 80 114 2 1 sky130_fd_sc_hd__dfxtp_1 $T=48180 34480 0 0 $X=47990 $Y=34240
X40 1 89 2 80 115 2 1 sky130_fd_sc_hd__dfxtp_1 $T=48640 34480 1 0 $X=48450 $Y=31520
X41 1 87 2 80 116 2 1 sky130_fd_sc_hd__dfxtp_1 $T=49560 18160 0 0 $X=49370 $Y=17920
X42 1 86 2 80 117 2 1 sky130_fd_sc_hd__dfxtp_1 $T=49560 23600 0 0 $X=49370 $Y=23360
X43 1 84 2 80 118 2 1 sky130_fd_sc_hd__dfxtp_1 $T=50020 18160 1 0 $X=49830 $Y=15200
X44 1 92 2 81 119 2 1 sky130_fd_sc_hd__dfxtp_1 $T=51400 23600 1 0 $X=51210 $Y=20640
X45 1 91 2 80 120 2 1 sky130_fd_sc_hd__dfxtp_1 $T=59220 18160 1 0 $X=59030 $Y=15200
X46 1 10 2 80 121 2 1 sky130_fd_sc_hd__dfxtp_1 $T=59220 18160 0 0 $X=59030 $Y=17920
X47 1 94 2 80 122 2 1 sky130_fd_sc_hd__dfxtp_1 $T=59220 29040 1 0 $X=59030 $Y=26080
X48 1 90 2 80 123 2 1 sky130_fd_sc_hd__dfxtp_1 $T=59220 29040 0 0 $X=59030 $Y=28800
X49 1 18 2 81 124 2 1 sky130_fd_sc_hd__dfxtp_1 $T=66120 23600 1 0 $X=65930 $Y=20640
X50 1 95 2 81 125 2 1 sky130_fd_sc_hd__dfxtp_1 $T=75320 18160 0 0 $X=75130 $Y=17920
X51 1 93 2 81 126 2 1 sky130_fd_sc_hd__dfxtp_1 $T=77160 23600 0 0 $X=76970 $Y=23360
X52 1 97 2 81 127 2 1 sky130_fd_sc_hd__dfxtp_1 $T=80840 23600 1 0 $X=80650 $Y=20640
X53 1 98 2 81 128 2 1 sky130_fd_sc_hd__dfxtp_1 $T=90960 23600 0 0 $X=90770 $Y=23360
X54 1 96 2 81 129 2 1 sky130_fd_sc_hd__dfxtp_1 $T=93720 18160 0 0 $X=93530 $Y=17920
X55 1 100 2 81 130 2 1 sky130_fd_sc_hd__dfxtp_1 $T=95560 23600 1 0 $X=95370 $Y=20640
X56 1 101 2 82 131 2 1 sky130_fd_sc_hd__dfxtp_1 $T=110280 23600 1 0 $X=110090 $Y=20640
X57 1 99 2 82 132 2 1 sky130_fd_sc_hd__dfxtp_1 $T=118100 18160 0 0 $X=117910 $Y=17920
X58 1 85 2 82 133 2 1 sky130_fd_sc_hd__dfxtp_1 $T=118100 23600 0 0 $X=117910 $Y=23360
X59 1 104 2 82 134 2 1 sky130_fd_sc_hd__dfxtp_1 $T=124540 23600 1 0 $X=124350 $Y=20640
X60 1 113 2 82 135 2 1 sky130_fd_sc_hd__dfxtp_1 $T=124540 29040 1 0 $X=124350 $Y=26080
X61 1 102 2 82 136 2 1 sky130_fd_sc_hd__dfxtp_1 $T=132820 18160 0 0 $X=132630 $Y=17920
X62 1 106 2 82 137 2 1 sky130_fd_sc_hd__dfxtp_1 $T=134660 23600 1 0 $X=134470 $Y=20640
X63 1 108 2 82 138 2 1 sky130_fd_sc_hd__dfxtp_1 $T=135120 29040 1 0 $X=134930 $Y=26080
X64 1 105 2 83 139 2 1 sky130_fd_sc_hd__dfxtp_1 $T=153060 18160 0 0 $X=152870 $Y=17920
X65 1 103 2 83 140 2 1 sky130_fd_sc_hd__dfxtp_1 $T=153520 18160 1 0 $X=153330 $Y=15200
X66 1 110 2 83 141 2 1 sky130_fd_sc_hd__dfxtp_1 $T=153520 23600 1 0 $X=153330 $Y=20640
X67 1 112 2 83 142 2 1 sky130_fd_sc_hd__dfxtp_1 $T=162260 23600 1 0 $X=162070 $Y=20640
X68 1 109 2 83 76 2 1 sky130_fd_sc_hd__dfxtp_1 $T=165480 18160 0 0 $X=165290 $Y=17920
X69 1 107 2 83 143 2 1 sky130_fd_sc_hd__dfxtp_1 $T=169160 18160 1 0 $X=168970 $Y=15200
X70 1 111 2 83 144 2 1 sky130_fd_sc_hd__dfxtp_1 $T=176980 23600 1 0 $X=176790 $Y=20640
X71 116 1 2 79 78 84 10 145 2 1 sky130_fd_sc_hd__a221o_1 $T=44500 18160 1 0 $X=44310 $Y=15200
X72 117 1 2 79 78 85 88 145 2 1 sky130_fd_sc_hd__a221o_1 $T=45880 23600 1 0 $X=45690 $Y=20640
X73 114 1 2 79 78 86 89 145 2 1 sky130_fd_sc_hd__a221o_1 $T=45880 29040 1 0 $X=45690 $Y=26080
X74 115 1 2 79 78 88 90 145 2 1 sky130_fd_sc_hd__a221o_1 $T=45880 29040 0 0 $X=45690 $Y=28800
X75 121 1 2 79 78 87 91 145 2 1 sky130_fd_sc_hd__a221o_1 $T=50480 12720 0 0 $X=50290 $Y=12480
X76 120 1 2 79 78 10 92 145 2 1 sky130_fd_sc_hd__a221o_1 $T=64280 12720 1 180 $X=60410 $Y=12480
X77 122 1 2 79 78 90 93 145 2 1 sky130_fd_sc_hd__a221o_1 $T=72100 18160 0 180 $X=68230 $Y=15200
X78 119 1 2 79 78 91 95 145 2 1 sky130_fd_sc_hd__a221o_1 $T=72100 18160 1 180 $X=68230 $Y=17920
X79 123 1 2 79 78 89 94 145 2 1 sky130_fd_sc_hd__a221o_1 $T=72100 29040 0 180 $X=68230 $Y=26080
X80 126 1 2 79 78 94 18 145 2 1 sky130_fd_sc_hd__a221o_1 $T=73940 29040 0 0 $X=73750 $Y=28800
X81 127 1 2 79 78 18 98 145 2 1 sky130_fd_sc_hd__a221o_1 $T=80380 29040 0 0 $X=80190 $Y=28800
X82 125 1 2 79 78 92 96 145 2 1 sky130_fd_sc_hd__a221o_1 $T=84980 18160 0 180 $X=81110 $Y=15200
X83 124 1 2 79 78 93 97 145 2 1 sky130_fd_sc_hd__a221o_1 $T=82680 18160 0 0 $X=82490 $Y=17920
X84 128 1 2 79 78 97 99 145 2 1 sky130_fd_sc_hd__a221o_1 $T=92800 12720 0 0 $X=92610 $Y=12480
X85 130 1 2 79 78 96 101 145 2 1 sky130_fd_sc_hd__a221o_1 $T=93720 29040 0 0 $X=93530 $Y=28800
X86 129 1 2 79 78 95 100 145 2 1 sky130_fd_sc_hd__a221o_1 $T=98320 18160 0 180 $X=94450 $Y=15200
X87 131 1 2 79 78 100 104 145 2 1 sky130_fd_sc_hd__a221o_1 $T=111200 18160 1 0 $X=111010 $Y=15200
X88 133 1 2 79 78 113 86 145 2 1 sky130_fd_sc_hd__a221o_1 $T=112580 23600 0 0 $X=112390 $Y=23360
X89 132 1 2 79 78 98 102 145 2 1 sky130_fd_sc_hd__a221o_1 $T=118100 12720 0 0 $X=117910 $Y=12480
X90 135 1 2 79 78 112 85 145 2 1 sky130_fd_sc_hd__a221o_1 $T=119480 29040 1 0 $X=119290 $Y=26080
X91 134 1 2 79 78 101 106 145 2 1 sky130_fd_sc_hd__a221o_1 $T=119480 29040 0 0 $X=119290 $Y=28800
X92 136 1 2 79 78 99 103 145 2 1 sky130_fd_sc_hd__a221o_1 $T=125460 18160 1 0 $X=125270 $Y=15200
X93 140 1 2 79 78 102 105 145 2 1 sky130_fd_sc_hd__a221o_1 $T=134660 18160 1 0 $X=134470 $Y=15200
X94 137 1 2 79 78 104 108 145 2 1 sky130_fd_sc_hd__a221o_1 $T=141560 23600 1 180 $X=137690 $Y=23360
X95 138 1 2 79 78 106 110 145 2 1 sky130_fd_sc_hd__a221o_1 $T=141560 29040 1 180 $X=137690 $Y=28800
X96 139 1 2 79 78 103 107 145 2 1 sky130_fd_sc_hd__a221o_1 $T=142480 18160 1 0 $X=142290 $Y=15200
X97 143 1 2 79 78 105 109 145 2 1 sky130_fd_sc_hd__a221o_1 $T=142480 18160 0 0 $X=142290 $Y=17920
X98 141 1 2 79 78 108 112 145 2 1 sky130_fd_sc_hd__a221o_1 $T=158580 23600 1 180 $X=154710 $Y=23360
X99 142 1 2 79 78 110 113 145 2 1 sky130_fd_sc_hd__a221o_1 $T=156740 29040 1 0 $X=156550 $Y=26080
X100 77 1 2 37 29 107 111 145 2 1 sky130_fd_sc_hd__a221o_1 $T=171460 12720 1 180 $X=167590 $Y=12480
X101 144 1 2 79 109 78 2 1 sky130_fd_sc_hd__a21o_1 $T=169160 23600 0 0 $X=168970 $Y=23360
X102 1 118 2 87 79 78 2 1 sky130_fd_sc_hd__or3_1 $T=45420 12720 0 0 $X=45230 $Y=12480
X103 1 145 2 29 2 1 sky130_fd_sc_hd__inv_2 $T=120400 34480 0 180 $X=118830 $Y=31520
X104 146 40 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 12720 1 0 $X=9810 $Y=9760
X105 147 41 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 12720 0 0 $X=9810 $Y=12480
X106 148 42 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 18160 1 0 $X=9810 $Y=15200
X107 149 43 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 18160 0 0 $X=9810 $Y=17920
X108 150 44 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 23600 1 0 $X=9810 $Y=20640
X109 151 45 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 23600 0 0 $X=9810 $Y=23360
X110 152 46 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 29040 1 0 $X=9810 $Y=26080
X111 153 47 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 29040 0 0 $X=9810 $Y=28800
X112 154 48 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 34480 1 0 $X=9810 $Y=31520
X113 155 49 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 34480 0 0 $X=9810 $Y=34240
X114 156 50 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 39920 1 0 $X=9810 $Y=36960
X115 157 51 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 39920 0 0 $X=9810 $Y=39680
X116 158 52 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 45360 1 0 $X=9810 $Y=42400
X117 159 53 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 45360 0 0 $X=9810 $Y=45120
X118 160 54 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 50800 1 0 $X=9810 $Y=47840
X119 161 55 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 50800 0 0 $X=9810 $Y=50560
X120 162 56 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 56240 1 0 $X=9810 $Y=53280
X121 163 57 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=10000 56240 0 0 $X=9810 $Y=56000
X122 164 58 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 12720 0 180 $X=189210 $Y=9760
X123 165 59 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 12720 1 180 $X=189210 $Y=12480
X124 166 60 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 18160 0 180 $X=189210 $Y=15200
X125 167 61 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 18160 1 180 $X=189210 $Y=17920
X126 168 62 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 23600 0 180 $X=189210 $Y=20640
X127 169 63 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 23600 1 180 $X=189210 $Y=23360
X128 170 64 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 29040 0 180 $X=189210 $Y=26080
X129 171 65 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 29040 1 180 $X=189210 $Y=28800
X130 172 66 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 34480 0 180 $X=189210 $Y=31520
X131 173 67 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 34480 1 180 $X=189210 $Y=34240
X132 174 68 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 39920 0 180 $X=189210 $Y=36960
X133 175 69 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 39920 1 180 $X=189210 $Y=39680
X134 176 70 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 45360 0 180 $X=189210 $Y=42400
X135 177 71 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 45360 1 180 $X=189210 $Y=45120
X136 178 72 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 50800 0 180 $X=189210 $Y=47840
X137 179 73 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 50800 1 180 $X=189210 $Y=50560
X138 180 74 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 56240 0 180 $X=189210 $Y=53280
X139 181 75 2 1 sky130_fd_sc_hd__tap_1_DigitalLDOLogic_gds $T=189860 56240 1 180 $X=189210 $Y=56000
X140 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=29320 12720 1 0 $X=29130 $Y=9760
X141 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=29320 12720 0 0 $X=29130 $Y=12480
X142 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=29320 18160 1 0 $X=29130 $Y=15200
X143 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=29320 18160 0 0 $X=29130 $Y=17920
X144 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=29320 23600 1 0 $X=29130 $Y=20640
X145 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=29320 23600 0 0 $X=29130 $Y=23360
X146 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=44040 18160 1 0 $X=43850 $Y=15200
X147 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=44040 18160 0 0 $X=43850 $Y=17920
X148 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=44040 23600 1 0 $X=43850 $Y=20640
X149 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=44040 23600 0 0 $X=43850 $Y=23360
X150 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=58760 12720 1 0 $X=58570 $Y=9760
X151 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=58760 12720 0 0 $X=58570 $Y=12480
X152 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=58760 18160 1 0 $X=58570 $Y=15200
X153 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=58760 18160 0 0 $X=58570 $Y=17920
X154 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=58760 23600 1 0 $X=58570 $Y=20640
X155 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=58760 23600 0 0 $X=58570 $Y=23360
X156 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=58760 29040 1 0 $X=58570 $Y=26080
X157 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=58760 29040 0 0 $X=58570 $Y=28800
X158 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=73480 12720 1 0 $X=73290 $Y=9760
X159 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=73480 12720 0 0 $X=73290 $Y=12480
X160 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=73480 18160 1 0 $X=73290 $Y=15200
X161 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=73480 18160 0 0 $X=73290 $Y=17920
X162 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=73480 23600 1 0 $X=73290 $Y=20640
X163 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=73480 23600 0 0 $X=73290 $Y=23360
X164 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=73480 29040 1 0 $X=73290 $Y=26080
X165 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=73480 29040 0 0 $X=73290 $Y=28800
X166 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=88200 12720 1 0 $X=88010 $Y=9760
X167 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=88200 12720 0 0 $X=88010 $Y=12480
X168 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=88200 18160 1 0 $X=88010 $Y=15200
X169 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=88200 18160 0 0 $X=88010 $Y=17920
X170 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=88200 23600 1 0 $X=88010 $Y=20640
X171 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=88200 23600 0 0 $X=88010 $Y=23360
X172 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=88200 29040 1 0 $X=88010 $Y=26080
X173 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=88200 29040 0 0 $X=88010 $Y=28800
X174 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=102920 12720 1 0 $X=102730 $Y=9760
X175 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=102920 12720 0 0 $X=102730 $Y=12480
X176 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=102920 18160 1 0 $X=102730 $Y=15200
X177 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=102920 18160 0 0 $X=102730 $Y=17920
X178 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=102920 29040 1 0 $X=102730 $Y=26080
X179 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=102920 29040 0 0 $X=102730 $Y=28800
X180 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 12720 1 0 $X=117450 $Y=9760
X181 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 12720 0 0 $X=117450 $Y=12480
X182 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 18160 1 0 $X=117450 $Y=15200
X183 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 18160 0 0 $X=117450 $Y=17920
X184 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 23600 1 0 $X=117450 $Y=20640
X185 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 23600 0 0 $X=117450 $Y=23360
X186 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 29040 1 0 $X=117450 $Y=26080
X187 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 29040 0 0 $X=117450 $Y=28800
X188 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 34480 1 0 $X=117450 $Y=31520
X189 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 34480 0 0 $X=117450 $Y=34240
X190 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 39920 1 0 $X=117450 $Y=36960
X191 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 39920 0 0 $X=117450 $Y=39680
X192 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 45360 1 0 $X=117450 $Y=42400
X193 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 45360 0 0 $X=117450 $Y=45120
X194 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 50800 1 0 $X=117450 $Y=47840
X195 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 50800 0 0 $X=117450 $Y=50560
X196 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 56240 1 0 $X=117450 $Y=53280
X197 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=117640 56240 0 0 $X=117450 $Y=56000
X198 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 12720 1 0 $X=132170 $Y=9760
X199 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 12720 0 0 $X=132170 $Y=12480
X200 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 23600 1 0 $X=132170 $Y=20640
X201 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 23600 0 0 $X=132170 $Y=23360
X202 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 29040 1 0 $X=132170 $Y=26080
X203 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 29040 0 0 $X=132170 $Y=28800
X204 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 34480 1 0 $X=132170 $Y=31520
X205 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 34480 0 0 $X=132170 $Y=34240
X206 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 39920 1 0 $X=132170 $Y=36960
X207 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 39920 0 0 $X=132170 $Y=39680
X208 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 45360 1 0 $X=132170 $Y=42400
X209 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 45360 0 0 $X=132170 $Y=45120
X210 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 50800 1 0 $X=132170 $Y=47840
X211 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 50800 0 0 $X=132170 $Y=50560
X212 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 56240 1 0 $X=132170 $Y=53280
X213 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=132360 56240 0 0 $X=132170 $Y=56000
X214 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 12720 1 0 $X=146890 $Y=9760
X215 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 12720 0 0 $X=146890 $Y=12480
X216 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 18160 1 0 $X=146890 $Y=15200
X217 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 18160 0 0 $X=146890 $Y=17920
X218 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 23600 1 0 $X=146890 $Y=20640
X219 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 23600 0 0 $X=146890 $Y=23360
X220 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 34480 1 0 $X=146890 $Y=31520
X221 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 34480 0 0 $X=146890 $Y=34240
X222 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 39920 1 0 $X=146890 $Y=36960
X223 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 39920 0 0 $X=146890 $Y=39680
X224 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 45360 1 0 $X=146890 $Y=42400
X225 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 45360 0 0 $X=146890 $Y=45120
X226 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 50800 1 0 $X=146890 $Y=47840
X227 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 50800 0 0 $X=146890 $Y=50560
X228 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 56240 1 0 $X=146890 $Y=53280
X229 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=147080 56240 0 0 $X=146890 $Y=56000
X230 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 12720 1 0 $X=161610 $Y=9760
X231 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 12720 0 0 $X=161610 $Y=12480
X232 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 18160 1 0 $X=161610 $Y=15200
X233 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 18160 0 0 $X=161610 $Y=17920
X234 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 23600 1 0 $X=161610 $Y=20640
X235 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 23600 0 0 $X=161610 $Y=23360
X236 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 34480 1 0 $X=161610 $Y=31520
X237 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 34480 0 0 $X=161610 $Y=34240
X238 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 39920 1 0 $X=161610 $Y=36960
X239 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 39920 0 0 $X=161610 $Y=39680
X240 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 45360 1 0 $X=161610 $Y=42400
X241 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 45360 0 0 $X=161610 $Y=45120
X242 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 50800 1 0 $X=161610 $Y=47840
X243 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 50800 0 0 $X=161610 $Y=50560
X244 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 56240 1 0 $X=161610 $Y=53280
X245 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=161800 56240 0 0 $X=161610 $Y=56000
X246 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 18160 1 0 $X=176330 $Y=15200
X247 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 18160 0 0 $X=176330 $Y=17920
X248 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 23600 1 0 $X=176330 $Y=20640
X249 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 23600 0 0 $X=176330 $Y=23360
X250 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 34480 1 0 $X=176330 $Y=31520
X251 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 34480 0 0 $X=176330 $Y=34240
X252 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 39920 1 0 $X=176330 $Y=36960
X253 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 39920 0 0 $X=176330 $Y=39680
X254 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 45360 1 0 $X=176330 $Y=42400
X255 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 45360 0 0 $X=176330 $Y=45120
X256 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 50800 1 0 $X=176330 $Y=47840
X257 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 50800 0 0 $X=176330 $Y=50560
X258 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 56240 1 0 $X=176330 $Y=53280
X259 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=176520 56240 0 0 $X=176330 $Y=56000
X260 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 12720 1 0 $X=188750 $Y=9760
X261 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 12720 0 0 $X=188750 $Y=12480
X262 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 18160 1 0 $X=188750 $Y=15200
X263 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 18160 0 0 $X=188750 $Y=17920
X264 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 23600 1 0 $X=188750 $Y=20640
X265 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 23600 0 0 $X=188750 $Y=23360
X266 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 29040 1 0 $X=188750 $Y=26080
X267 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 29040 0 0 $X=188750 $Y=28800
X268 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 34480 1 0 $X=188750 $Y=31520
X269 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 34480 0 0 $X=188750 $Y=34240
X270 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 39920 1 0 $X=188750 $Y=36960
X271 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 39920 0 0 $X=188750 $Y=39680
X272 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 45360 1 0 $X=188750 $Y=42400
X273 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 45360 0 0 $X=188750 $Y=45120
X274 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 50800 1 0 $X=188750 $Y=47840
X275 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 50800 0 0 $X=188750 $Y=50560
X276 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 56240 1 0 $X=188750 $Y=53280
X277 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1_DigitalLDOLogic_gds $T=188940 56240 0 0 $X=188750 $Y=56000
X278 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 12720 1 0 $X=10270 $Y=9760
X279 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 12720 0 0 $X=10270 $Y=12480
X280 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 18160 1 0 $X=10270 $Y=15200
X281 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 18160 0 0 $X=10270 $Y=17920
X282 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 23600 1 0 $X=10270 $Y=20640
X283 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 23600 0 0 $X=10270 $Y=23360
X284 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 29040 1 0 $X=10270 $Y=26080
X285 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 29040 0 0 $X=10270 $Y=28800
X286 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 34480 1 0 $X=10270 $Y=31520
X287 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 34480 0 0 $X=10270 $Y=34240
X288 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 39920 1 0 $X=10270 $Y=36960
X289 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 39920 0 0 $X=10270 $Y=39680
X290 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 45360 1 0 $X=10270 $Y=42400
X291 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 45360 0 0 $X=10270 $Y=45120
X292 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 50800 1 0 $X=10270 $Y=47840
X293 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 50800 0 0 $X=10270 $Y=50560
X294 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 56240 1 0 $X=10270 $Y=53280
X295 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=10460 56240 0 0 $X=10270 $Y=56000
X296 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=15060 12720 0 0 $X=14870 $Y=12480
X297 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=15060 18160 1 0 $X=14870 $Y=15200
X298 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=15060 23600 0 0 $X=14870 $Y=23360
X299 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=24720 12720 0 0 $X=24530 $Y=12480
X300 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=24720 18160 1 0 $X=24530 $Y=15200
X301 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=26560 23600 0 0 $X=26370 $Y=23360
X302 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=29780 12720 0 0 $X=29590 $Y=12480
X303 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=38060 12720 0 0 $X=37870 $Y=12480
X304 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=41280 18160 1 0 $X=41090 $Y=15200
X305 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=44500 34480 1 0 $X=44310 $Y=31520
X306 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=47720 12720 0 0 $X=47530 $Y=12480
X307 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=54160 12720 0 0 $X=53970 $Y=12480
X308 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=56000 34480 1 0 $X=55810 $Y=31520
X309 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=61520 23600 1 0 $X=61330 $Y=20640
X310 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=62900 23600 0 0 $X=62710 $Y=23360
X311 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=77620 29040 0 0 $X=77430 $Y=28800
X312 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=84060 29040 0 0 $X=83870 $Y=28800
X313 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=88660 12720 1 0 $X=88470 $Y=9760
X314 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=88660 12720 0 0 $X=88470 $Y=12480
X315 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=88660 18160 1 0 $X=88470 $Y=15200
X316 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=98320 18160 1 0 $X=98130 $Y=15200
X317 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=98320 23600 0 0 $X=98130 $Y=23360
X318 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=100160 12720 0 0 $X=99970 $Y=12480
X319 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=103380 18160 0 0 $X=103190 $Y=17920
X320 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=114880 18160 1 0 $X=114690 $Y=15200
X321 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=114880 18160 0 0 $X=114690 $Y=17920
X322 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=121780 23600 1 0 $X=121590 $Y=20640
X323 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=129600 34480 1 0 $X=129410 $Y=31520
X324 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=138340 18160 1 0 $X=138150 $Y=15200
X325 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=142480 29040 1 0 $X=142290 $Y=26080
X326 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=147540 18160 1 0 $X=147350 $Y=15200
X327 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=147540 23600 1 0 $X=147350 $Y=20640
X328 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=157660 12720 1 0 $X=157470 $Y=9760
X329 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=171920 23600 0 0 $X=171730 $Y=23360
X330 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=172380 12720 1 0 $X=172190 $Y=9760
X331 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=184340 23600 1 0 $X=184150 $Y=20640
X332 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 12720 1 0 $X=185990 $Y=9760
X333 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 12720 0 0 $X=185990 $Y=12480
X334 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 18160 1 0 $X=185990 $Y=15200
X335 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 18160 0 0 $X=185990 $Y=17920
X336 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 29040 1 0 $X=185990 $Y=26080
X337 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 29040 0 0 $X=185990 $Y=28800
X338 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 34480 1 0 $X=185990 $Y=31520
X339 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 34480 0 0 $X=185990 $Y=34240
X340 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 39920 1 0 $X=185990 $Y=36960
X341 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 39920 0 0 $X=185990 $Y=39680
X342 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 45360 1 0 $X=185990 $Y=42400
X343 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 45360 0 0 $X=185990 $Y=45120
X344 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 50800 1 0 $X=185990 $Y=47840
X345 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 50800 0 0 $X=185990 $Y=50560
X346 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 56240 1 0 $X=185990 $Y=53280
X347 1 2 2 1 sky130_fd_sc_hd__decap_6_DigitalLDOLogic_gds $T=186180 56240 0 0 $X=185990 $Y=56000
X348 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=17820 12720 0 0 $X=17630 $Y=12480
X349 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=17820 18160 1 0 $X=17630 $Y=15200
X350 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=19660 23600 0 0 $X=19470 $Y=23360
X351 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=27940 12720 1 0 $X=27750 $Y=9760
X352 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=27940 18160 0 0 $X=27750 $Y=17920
X353 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=27940 23600 1 0 $X=27750 $Y=20640
X354 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=42660 18160 0 0 $X=42470 $Y=17920
X355 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=42660 23600 1 0 $X=42470 $Y=20640
X356 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=42660 23600 0 0 $X=42470 $Y=23360
X357 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=44500 23600 1 0 $X=44310 $Y=20640
X358 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=44500 29040 1 0 $X=44310 $Y=26080
X359 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=44500 29040 0 0 $X=44310 $Y=28800
X360 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=46340 12720 1 0 $X=46150 $Y=9760
X361 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=47260 34480 1 0 $X=47070 $Y=31520
X362 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=48180 18160 0 0 $X=47990 $Y=17920
X363 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=48180 23600 0 0 $X=47990 $Y=23360
X364 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 18160 1 0 $X=57190 $Y=15200
X365 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 34480 0 0 $X=57190 $Y=34240
X366 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 39920 1 0 $X=57190 $Y=36960
X367 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 39920 0 0 $X=57190 $Y=39680
X368 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 45360 1 0 $X=57190 $Y=42400
X369 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 45360 0 0 $X=57190 $Y=45120
X370 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 50800 1 0 $X=57190 $Y=47840
X371 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 50800 0 0 $X=57190 $Y=50560
X372 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 56240 1 0 $X=57190 $Y=53280
X373 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=57380 56240 0 0 $X=57190 $Y=56000
X374 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=59220 12720 0 0 $X=59030 $Y=12480
X375 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=61060 12720 1 0 $X=60870 $Y=9760
X376 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=64280 12720 0 0 $X=64090 $Y=12480
X377 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=71180 12720 0 0 $X=70990 $Y=12480
X378 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=71180 23600 0 0 $X=70990 $Y=23360
X379 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=72100 18160 1 0 $X=71910 $Y=15200
X380 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=72100 18160 0 0 $X=71910 $Y=17920
X381 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=72100 29040 1 0 $X=71910 $Y=26080
X382 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=72100 29040 0 0 $X=71910 $Y=28800
X383 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=73940 18160 0 0 $X=73750 $Y=17920
X384 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=75780 23600 0 0 $X=75590 $Y=23360
X385 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=81300 12720 1 0 $X=81110 $Y=9760
X386 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=86820 12720 0 0 $X=86630 $Y=12480
X387 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=86820 18160 1 0 $X=86630 $Y=15200
X388 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=86820 29040 1 0 $X=86630 $Y=26080
X389 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=86820 29040 0 0 $X=86630 $Y=28800
X390 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=88660 23600 0 0 $X=88470 $Y=23360
X391 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=91420 12720 0 0 $X=91230 $Y=12480
X392 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=92340 18160 0 0 $X=92150 $Y=17920
X393 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=92340 29040 0 0 $X=92150 $Y=28800
X394 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=93260 18160 1 0 $X=93070 $Y=15200
X395 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=94180 23600 1 0 $X=93990 $Y=20640
X396 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=101540 29040 1 0 $X=101350 $Y=26080
X397 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=107980 18160 0 0 $X=107790 $Y=17920
X398 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=108900 12720 0 0 $X=108710 $Y=12480
X399 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=108900 18160 1 0 $X=108710 $Y=15200
X400 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=108900 23600 1 0 $X=108710 $Y=20640
X401 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=116260 12720 1 0 $X=116070 $Y=9760
X402 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=116260 23600 0 0 $X=116070 $Y=23360
X403 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=118100 29040 1 0 $X=117910 $Y=26080
X404 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=118100 29040 0 0 $X=117910 $Y=28800
X405 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=123160 29040 1 0 $X=122970 $Y=26080
X406 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 12720 1 0 $X=130790 $Y=9760
X407 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 12720 0 0 $X=130790 $Y=12480
X408 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 23600 0 0 $X=130790 $Y=23360
X409 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 34480 0 0 $X=130790 $Y=34240
X410 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 39920 1 0 $X=130790 $Y=36960
X411 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 39920 0 0 $X=130790 $Y=39680
X412 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 45360 1 0 $X=130790 $Y=42400
X413 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 45360 0 0 $X=130790 $Y=45120
X414 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 50800 1 0 $X=130790 $Y=47840
X415 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 50800 0 0 $X=130790 $Y=50560
X416 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 56240 1 0 $X=130790 $Y=53280
X417 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=130980 56240 0 0 $X=130790 $Y=56000
X418 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=132820 29040 1 0 $X=132630 $Y=26080
X419 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=136500 23600 0 0 $X=136310 $Y=23360
X420 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=136500 29040 0 0 $X=136310 $Y=28800
X421 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=140180 18160 0 0 $X=139990 $Y=17920
X422 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=141100 18160 1 0 $X=140910 $Y=15200
X423 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=144780 12720 0 0 $X=144590 $Y=12480
X424 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 12720 1 0 $X=145510 $Y=9760
X425 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 23600 1 0 $X=145510 $Y=20640
X426 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 34480 1 0 $X=145510 $Y=31520
X427 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 34480 0 0 $X=145510 $Y=34240
X428 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 39920 1 0 $X=145510 $Y=36960
X429 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 39920 0 0 $X=145510 $Y=39680
X430 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 45360 1 0 $X=145510 $Y=42400
X431 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 45360 0 0 $X=145510 $Y=45120
X432 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 50800 1 0 $X=145510 $Y=47840
X433 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 50800 0 0 $X=145510 $Y=50560
X434 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 56240 1 0 $X=145510 $Y=53280
X435 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=145700 56240 0 0 $X=145510 $Y=56000
X436 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=152140 18160 1 0 $X=151950 $Y=15200
X437 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=152140 23600 1 0 $X=151950 $Y=20640
X438 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 12720 1 0 $X=160230 $Y=9760
X439 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 12720 0 0 $X=160230 $Y=12480
X440 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 18160 0 0 $X=160230 $Y=17920
X441 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 23600 0 0 $X=160230 $Y=23360
X442 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 34480 1 0 $X=160230 $Y=31520
X443 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 34480 0 0 $X=160230 $Y=34240
X444 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 39920 1 0 $X=160230 $Y=36960
X445 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 39920 0 0 $X=160230 $Y=39680
X446 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 45360 1 0 $X=160230 $Y=42400
X447 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 45360 0 0 $X=160230 $Y=45120
X448 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 50800 1 0 $X=160230 $Y=47840
X449 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 50800 0 0 $X=160230 $Y=50560
X450 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 56240 1 0 $X=160230 $Y=53280
X451 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=160420 56240 0 0 $X=160230 $Y=56000
X452 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=167780 18160 1 0 $X=167590 $Y=15200
X453 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=167780 23600 0 0 $X=167590 $Y=23360
X454 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 12720 1 0 $X=174950 $Y=9760
X455 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 12720 0 0 $X=174950 $Y=12480
X456 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 23600 1 0 $X=174950 $Y=20640
X457 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 34480 1 0 $X=174950 $Y=31520
X458 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 34480 0 0 $X=174950 $Y=34240
X459 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 39920 1 0 $X=174950 $Y=36960
X460 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 39920 0 0 $X=174950 $Y=39680
X461 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 45360 1 0 $X=174950 $Y=42400
X462 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 45360 0 0 $X=174950 $Y=45120
X463 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 50800 1 0 $X=174950 $Y=47840
X464 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 50800 0 0 $X=174950 $Y=50560
X465 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 56240 1 0 $X=174950 $Y=53280
X466 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=175140 56240 0 0 $X=174950 $Y=56000
X467 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=178820 23600 0 0 $X=178630 $Y=23360
X468 1 2 2 1 sky130_fd_sc_hd__decap_3_DigitalLDOLogic_gds $T=187560 23600 0 0 $X=187370 $Y=23360
X469 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 12720 1 0 $X=14870 $Y=9760
X470 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 18160 0 0 $X=14870 $Y=17920
X471 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 23600 1 0 $X=14870 $Y=20640
X472 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 29040 1 0 $X=14870 $Y=26080
X473 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 29040 0 0 $X=14870 $Y=28800
X474 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 34480 1 0 $X=14870 $Y=31520
X475 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 34480 0 0 $X=14870 $Y=34240
X476 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 39920 1 0 $X=14870 $Y=36960
X477 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 39920 0 0 $X=14870 $Y=39680
X478 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 45360 1 0 $X=14870 $Y=42400
X479 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 45360 0 0 $X=14870 $Y=45120
X480 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 50800 1 0 $X=14870 $Y=47840
X481 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 50800 0 0 $X=14870 $Y=50560
X482 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 56240 1 0 $X=14870 $Y=53280
X483 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=15060 56240 0 0 $X=14870 $Y=56000
X484 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 12720 1 0 $X=20390 $Y=9760
X485 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 18160 0 0 $X=20390 $Y=17920
X486 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 23600 1 0 $X=20390 $Y=20640
X487 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 29040 1 0 $X=20390 $Y=26080
X488 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 29040 0 0 $X=20390 $Y=28800
X489 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 34480 1 0 $X=20390 $Y=31520
X490 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 34480 0 0 $X=20390 $Y=34240
X491 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 39920 1 0 $X=20390 $Y=36960
X492 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 39920 0 0 $X=20390 $Y=39680
X493 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 45360 1 0 $X=20390 $Y=42400
X494 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 45360 0 0 $X=20390 $Y=45120
X495 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 50800 1 0 $X=20390 $Y=47840
X496 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 50800 0 0 $X=20390 $Y=50560
X497 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 56240 1 0 $X=20390 $Y=53280
X498 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=20580 56240 0 0 $X=20390 $Y=56000
X499 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=29780 18160 0 0 $X=29590 $Y=17920
X500 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=29780 23600 1 0 $X=29590 $Y=20640
X501 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=29780 23600 0 0 $X=29590 $Y=23360
X502 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 12720 1 0 $X=35110 $Y=9760
X503 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 18160 0 0 $X=35110 $Y=17920
X504 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 23600 1 0 $X=35110 $Y=20640
X505 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 23600 0 0 $X=35110 $Y=23360
X506 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 29040 0 0 $X=35110 $Y=28800
X507 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 34480 1 0 $X=35110 $Y=31520
X508 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 34480 0 0 $X=35110 $Y=34240
X509 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 39920 1 0 $X=35110 $Y=36960
X510 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 39920 0 0 $X=35110 $Y=39680
X511 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 45360 1 0 $X=35110 $Y=42400
X512 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 45360 0 0 $X=35110 $Y=45120
X513 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 50800 1 0 $X=35110 $Y=47840
X514 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 50800 0 0 $X=35110 $Y=50560
X515 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 56240 1 0 $X=35110 $Y=53280
X516 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=35300 56240 0 0 $X=35110 $Y=56000
X517 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=44500 39920 1 0 $X=44310 $Y=36960
X518 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=44500 39920 0 0 $X=44310 $Y=39680
X519 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=44500 45360 1 0 $X=44310 $Y=42400
X520 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=44500 45360 0 0 $X=44310 $Y=45120
X521 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=44500 50800 1 0 $X=44310 $Y=47840
X522 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=44500 50800 0 0 $X=44310 $Y=50560
X523 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=44500 56240 1 0 $X=44310 $Y=53280
X524 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=44500 56240 0 0 $X=44310 $Y=56000
X525 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=49560 29040 1 0 $X=49370 $Y=26080
X526 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=49560 29040 0 0 $X=49370 $Y=28800
X527 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=50020 39920 1 0 $X=49830 $Y=36960
X528 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=50020 39920 0 0 $X=49830 $Y=39680
X529 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=50020 45360 1 0 $X=49830 $Y=42400
X530 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=50020 45360 0 0 $X=49830 $Y=45120
X531 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=50020 50800 1 0 $X=49830 $Y=47840
X532 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=50020 50800 0 0 $X=49830 $Y=50560
X533 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=50020 56240 1 0 $X=49830 $Y=53280
X534 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=50020 56240 0 0 $X=49830 $Y=56000
X535 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=53240 12720 1 0 $X=53050 $Y=9760
X536 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 34480 1 0 $X=64550 $Y=31520
X537 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 34480 0 0 $X=64550 $Y=34240
X538 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 39920 1 0 $X=64550 $Y=36960
X539 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 39920 0 0 $X=64550 $Y=39680
X540 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 45360 1 0 $X=64550 $Y=42400
X541 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 45360 0 0 $X=64550 $Y=45120
X542 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 50800 1 0 $X=64550 $Y=47840
X543 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 50800 0 0 $X=64550 $Y=50560
X544 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 56240 1 0 $X=64550 $Y=53280
X545 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=64740 56240 0 0 $X=64550 $Y=56000
X546 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=66580 29040 0 0 $X=66390 $Y=28800
X547 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=67960 12720 1 0 $X=67770 $Y=9760
X548 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 12720 0 0 $X=73750 $Y=12480
X549 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 23600 1 0 $X=73750 $Y=20640
X550 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 29040 1 0 $X=73750 $Y=26080
X551 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 34480 1 0 $X=73750 $Y=31520
X552 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 34480 0 0 $X=73750 $Y=34240
X553 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 39920 1 0 $X=73750 $Y=36960
X554 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 39920 0 0 $X=73750 $Y=39680
X555 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 45360 1 0 $X=73750 $Y=42400
X556 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 45360 0 0 $X=73750 $Y=45120
X557 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 50800 1 0 $X=73750 $Y=47840
X558 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 50800 0 0 $X=73750 $Y=50560
X559 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 56240 1 0 $X=73750 $Y=53280
X560 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=73940 56240 0 0 $X=73750 $Y=56000
X561 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 12720 0 0 $X=79270 $Y=12480
X562 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 29040 1 0 $X=79270 $Y=26080
X563 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 34480 1 0 $X=79270 $Y=31520
X564 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 34480 0 0 $X=79270 $Y=34240
X565 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 39920 1 0 $X=79270 $Y=36960
X566 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 39920 0 0 $X=79270 $Y=39680
X567 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 45360 1 0 $X=79270 $Y=42400
X568 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 45360 0 0 $X=79270 $Y=45120
X569 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 50800 1 0 $X=79270 $Y=47840
X570 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 50800 0 0 $X=79270 $Y=50560
X571 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 56240 1 0 $X=79270 $Y=53280
X572 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=79460 56240 0 0 $X=79270 $Y=56000
X573 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=88660 23600 1 0 $X=88470 $Y=20640
X574 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=88660 29040 1 0 $X=88470 $Y=26080
X575 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 29040 1 0 $X=93990 $Y=26080
X576 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 34480 1 0 $X=93990 $Y=31520
X577 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 34480 0 0 $X=93990 $Y=34240
X578 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 39920 1 0 $X=93990 $Y=36960
X579 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 39920 0 0 $X=93990 $Y=39680
X580 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 45360 1 0 $X=93990 $Y=42400
X581 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 45360 0 0 $X=93990 $Y=45120
X582 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 50800 1 0 $X=93990 $Y=47840
X583 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 50800 0 0 $X=93990 $Y=50560
X584 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 56240 1 0 $X=93990 $Y=53280
X585 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=94180 56240 0 0 $X=93990 $Y=56000
X586 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=97400 29040 0 0 $X=97210 $Y=28800
X587 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 12720 1 0 $X=103190 $Y=9760
X588 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 29040 1 0 $X=103190 $Y=26080
X589 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 29040 0 0 $X=103190 $Y=28800
X590 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 34480 1 0 $X=103190 $Y=31520
X591 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 34480 0 0 $X=103190 $Y=34240
X592 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 39920 1 0 $X=103190 $Y=36960
X593 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 39920 0 0 $X=103190 $Y=39680
X594 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 45360 1 0 $X=103190 $Y=42400
X595 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 45360 0 0 $X=103190 $Y=45120
X596 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 50800 1 0 $X=103190 $Y=47840
X597 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 50800 0 0 $X=103190 $Y=50560
X598 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 56240 1 0 $X=103190 $Y=53280
X599 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=103380 56240 0 0 $X=103190 $Y=56000
X600 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 12720 1 0 $X=108710 $Y=9760
X601 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 29040 1 0 $X=108710 $Y=26080
X602 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 29040 0 0 $X=108710 $Y=28800
X603 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 34480 1 0 $X=108710 $Y=31520
X604 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 34480 0 0 $X=108710 $Y=34240
X605 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 39920 1 0 $X=108710 $Y=36960
X606 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 39920 0 0 $X=108710 $Y=39680
X607 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 45360 1 0 $X=108710 $Y=42400
X608 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 45360 0 0 $X=108710 $Y=45120
X609 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 50800 1 0 $X=108710 $Y=47840
X610 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 50800 0 0 $X=108710 $Y=50560
X611 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 56240 1 0 $X=108710 $Y=53280
X612 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=108900 56240 0 0 $X=108710 $Y=56000
X613 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 34480 0 0 $X=117910 $Y=34240
X614 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 39920 1 0 $X=117910 $Y=36960
X615 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 39920 0 0 $X=117910 $Y=39680
X616 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 45360 1 0 $X=117910 $Y=42400
X617 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 45360 0 0 $X=117910 $Y=45120
X618 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 50800 1 0 $X=117910 $Y=47840
X619 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 50800 0 0 $X=117910 $Y=50560
X620 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 56240 1 0 $X=117910 $Y=53280
X621 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=118100 56240 0 0 $X=117910 $Y=56000
X622 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=120400 34480 1 0 $X=120210 $Y=31520
X623 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=121780 12720 0 0 $X=121590 $Y=12480
X624 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123160 29040 0 0 $X=122970 $Y=28800
X625 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 12720 1 0 $X=123430 $Y=9760
X626 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 34480 0 0 $X=123430 $Y=34240
X627 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 39920 1 0 $X=123430 $Y=36960
X628 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 39920 0 0 $X=123430 $Y=39680
X629 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 45360 1 0 $X=123430 $Y=42400
X630 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 45360 0 0 $X=123430 $Y=45120
X631 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 50800 1 0 $X=123430 $Y=47840
X632 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 50800 0 0 $X=123430 $Y=50560
X633 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 56240 1 0 $X=123430 $Y=53280
X634 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=123620 56240 0 0 $X=123430 $Y=56000
X635 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=125460 18160 0 0 $X=125270 $Y=17920
X636 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=125460 23600 0 0 $X=125270 $Y=23360
X637 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 12720 1 0 $X=132630 $Y=9760
X638 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 34480 1 0 $X=132630 $Y=31520
X639 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 34480 0 0 $X=132630 $Y=34240
X640 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 39920 1 0 $X=132630 $Y=36960
X641 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 39920 0 0 $X=132630 $Y=39680
X642 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 45360 1 0 $X=132630 $Y=42400
X643 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 45360 0 0 $X=132630 $Y=45120
X644 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 50800 1 0 $X=132630 $Y=47840
X645 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 50800 0 0 $X=132630 $Y=50560
X646 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 56240 1 0 $X=132630 $Y=53280
X647 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=132820 56240 0 0 $X=132630 $Y=56000
X648 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 34480 1 0 $X=138150 $Y=31520
X649 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 34480 0 0 $X=138150 $Y=34240
X650 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 39920 1 0 $X=138150 $Y=36960
X651 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 39920 0 0 $X=138150 $Y=39680
X652 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 45360 1 0 $X=138150 $Y=42400
X653 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 45360 0 0 $X=138150 $Y=45120
X654 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 50800 1 0 $X=138150 $Y=47840
X655 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 50800 0 0 $X=138150 $Y=50560
X656 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 56240 1 0 $X=138150 $Y=53280
X657 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=138340 56240 0 0 $X=138150 $Y=56000
X658 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=141560 23600 0 0 $X=141370 $Y=23360
X659 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=141560 29040 0 0 $X=141370 $Y=28800
X660 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 12720 0 0 $X=147350 $Y=12480
X661 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 18160 0 0 $X=147350 $Y=17920
X662 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 34480 1 0 $X=147350 $Y=31520
X663 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 34480 0 0 $X=147350 $Y=34240
X664 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 39920 1 0 $X=147350 $Y=36960
X665 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 39920 0 0 $X=147350 $Y=39680
X666 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 45360 1 0 $X=147350 $Y=42400
X667 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 45360 0 0 $X=147350 $Y=45120
X668 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 50800 1 0 $X=147350 $Y=47840
X669 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 50800 0 0 $X=147350 $Y=50560
X670 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 56240 1 0 $X=147350 $Y=53280
X671 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=147540 56240 0 0 $X=147350 $Y=56000
X672 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 12720 0 0 $X=152870 $Y=12480
X673 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 29040 0 0 $X=152870 $Y=28800
X674 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 34480 1 0 $X=152870 $Y=31520
X675 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 34480 0 0 $X=152870 $Y=34240
X676 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 39920 1 0 $X=152870 $Y=36960
X677 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 39920 0 0 $X=152870 $Y=39680
X678 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 45360 1 0 $X=152870 $Y=42400
X679 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 45360 0 0 $X=152870 $Y=45120
X680 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 50800 1 0 $X=152870 $Y=47840
X681 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 50800 0 0 $X=152870 $Y=50560
X682 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 56240 1 0 $X=152870 $Y=53280
X683 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=153060 56240 0 0 $X=152870 $Y=56000
X684 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 12720 0 0 $X=162070 $Y=12480
X685 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 23600 0 0 $X=162070 $Y=23360
X686 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 29040 1 0 $X=162070 $Y=26080
X687 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 29040 0 0 $X=162070 $Y=28800
X688 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 34480 1 0 $X=162070 $Y=31520
X689 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 34480 0 0 $X=162070 $Y=34240
X690 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 39920 1 0 $X=162070 $Y=36960
X691 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 39920 0 0 $X=162070 $Y=39680
X692 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 45360 1 0 $X=162070 $Y=42400
X693 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 45360 0 0 $X=162070 $Y=45120
X694 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 50800 1 0 $X=162070 $Y=47840
X695 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 50800 0 0 $X=162070 $Y=50560
X696 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 56240 1 0 $X=162070 $Y=53280
X697 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=162260 56240 0 0 $X=162070 $Y=56000
X698 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 29040 1 0 $X=167590 $Y=26080
X699 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 29040 0 0 $X=167590 $Y=28800
X700 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 34480 1 0 $X=167590 $Y=31520
X701 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 34480 0 0 $X=167590 $Y=34240
X702 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 39920 1 0 $X=167590 $Y=36960
X703 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 39920 0 0 $X=167590 $Y=39680
X704 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 45360 1 0 $X=167590 $Y=42400
X705 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 45360 0 0 $X=167590 $Y=45120
X706 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 50800 1 0 $X=167590 $Y=47840
X707 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 50800 0 0 $X=167590 $Y=50560
X708 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 56240 1 0 $X=167590 $Y=53280
X709 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=167780 56240 0 0 $X=167590 $Y=56000
X710 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 18160 0 0 $X=176790 $Y=17920
X711 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 34480 1 0 $X=176790 $Y=31520
X712 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 34480 0 0 $X=176790 $Y=34240
X713 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 39920 1 0 $X=176790 $Y=36960
X714 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 39920 0 0 $X=176790 $Y=39680
X715 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 45360 1 0 $X=176790 $Y=42400
X716 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 45360 0 0 $X=176790 $Y=45120
X717 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 50800 1 0 $X=176790 $Y=47840
X718 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 50800 0 0 $X=176790 $Y=50560
X719 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 56240 1 0 $X=176790 $Y=53280
X720 1 2 2 1 sky130_fd_sc_hd__decap_12_DigitalLDOLogic_gds $T=176980 56240 0 0 $X=176790 $Y=56000
X721 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=17820 23600 0 0 $X=17630 $Y=23360
X722 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=26100 12720 1 0 $X=25910 $Y=9760
X723 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=26100 18160 0 0 $X=25910 $Y=17920
X724 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=26100 23600 1 0 $X=25910 $Y=20640
X725 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=27480 12720 0 0 $X=27290 $Y=12480
X726 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=27480 18160 1 0 $X=27290 $Y=15200
X727 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 12720 1 0 $X=40630 $Y=9760
X728 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 12720 0 0 $X=40630 $Y=12480
X729 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 18160 0 0 $X=40630 $Y=17920
X730 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 23600 1 0 $X=40630 $Y=20640
X731 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 23600 0 0 $X=40630 $Y=23360
X732 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 29040 1 0 $X=40630 $Y=26080
X733 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 29040 0 0 $X=40630 $Y=28800
X734 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 34480 1 0 $X=40630 $Y=31520
X735 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 34480 0 0 $X=40630 $Y=34240
X736 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 39920 1 0 $X=40630 $Y=36960
X737 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 39920 0 0 $X=40630 $Y=39680
X738 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 45360 1 0 $X=40630 $Y=42400
X739 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 45360 0 0 $X=40630 $Y=45120
X740 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 50800 1 0 $X=40630 $Y=47840
X741 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 50800 0 0 $X=40630 $Y=50560
X742 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 56240 1 0 $X=40630 $Y=53280
X743 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=40820 56240 0 0 $X=40630 $Y=56000
X744 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=44500 12720 1 0 $X=44310 $Y=9760
X745 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=48180 18160 1 0 $X=47990 $Y=15200
X746 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=49560 23600 1 0 $X=49370 $Y=20640
X747 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 34480 0 0 $X=55350 $Y=34240
X748 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 39920 1 0 $X=55350 $Y=36960
X749 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 39920 0 0 $X=55350 $Y=39680
X750 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 45360 1 0 $X=55350 $Y=42400
X751 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 45360 0 0 $X=55350 $Y=45120
X752 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 50800 1 0 $X=55350 $Y=47840
X753 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 50800 0 0 $X=55350 $Y=50560
X754 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 56240 1 0 $X=55350 $Y=53280
X755 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=55540 56240 0 0 $X=55350 $Y=56000
X756 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=56920 12720 0 0 $X=56730 $Y=12480
X757 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=56920 18160 0 0 $X=56730 $Y=17920
X758 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=56920 23600 0 0 $X=56730 $Y=23360
X759 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=59220 12720 1 0 $X=59030 $Y=9760
X760 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=64280 23600 1 0 $X=64090 $Y=20640
X761 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=66580 18160 1 0 $X=66390 $Y=15200
X762 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=66580 18160 0 0 $X=66390 $Y=17920
X763 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=66580 29040 1 0 $X=66390 $Y=26080
X764 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 34480 1 0 $X=70070 $Y=31520
X765 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 34480 0 0 $X=70070 $Y=34240
X766 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 39920 1 0 $X=70070 $Y=36960
X767 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 39920 0 0 $X=70070 $Y=39680
X768 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 45360 1 0 $X=70070 $Y=42400
X769 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 45360 0 0 $X=70070 $Y=45120
X770 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 50800 1 0 $X=70070 $Y=47840
X771 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 50800 0 0 $X=70070 $Y=50560
X772 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 56240 1 0 $X=70070 $Y=53280
X773 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=70260 56240 0 0 $X=70070 $Y=56000
X774 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=73940 23600 0 0 $X=73750 $Y=23360
X775 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=79460 12720 1 0 $X=79270 $Y=9760
X776 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=79460 18160 1 0 $X=79270 $Y=15200
X777 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=84980 12720 0 0 $X=84790 $Y=12480
X778 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=84980 18160 1 0 $X=84790 $Y=15200
X779 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=84980 29040 1 0 $X=84790 $Y=26080
X780 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=86360 18160 0 0 $X=86170 $Y=17920
X781 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=91420 18160 1 0 $X=91230 $Y=15200
X782 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 29040 1 0 $X=99510 $Y=26080
X783 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 34480 1 0 $X=99510 $Y=31520
X784 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 34480 0 0 $X=99510 $Y=34240
X785 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 39920 1 0 $X=99510 $Y=36960
X786 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 39920 0 0 $X=99510 $Y=39680
X787 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 45360 1 0 $X=99510 $Y=42400
X788 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 45360 0 0 $X=99510 $Y=45120
X789 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 50800 1 0 $X=99510 $Y=47840
X790 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 50800 0 0 $X=99510 $Y=50560
X791 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 56240 1 0 $X=99510 $Y=53280
X792 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=99700 56240 0 0 $X=99510 $Y=56000
X793 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=101080 18160 1 0 $X=100890 $Y=15200
X794 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=101080 18160 0 0 $X=100890 $Y=17920
X795 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=101080 23600 0 0 $X=100890 $Y=23360
X796 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=106140 18160 0 0 $X=105950 $Y=17920
X797 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=114420 12720 1 0 $X=114230 $Y=9760
X798 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=115800 12720 0 0 $X=115610 $Y=12480
X799 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=123620 18160 1 0 $X=123430 $Y=15200
X800 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 12720 1 0 $X=128950 $Y=9760
X801 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 18160 1 0 $X=128950 $Y=15200
X802 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 34480 0 0 $X=128950 $Y=34240
X803 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 39920 1 0 $X=128950 $Y=36960
X804 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 39920 0 0 $X=128950 $Y=39680
X805 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 45360 1 0 $X=128950 $Y=42400
X806 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 45360 0 0 $X=128950 $Y=45120
X807 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 50800 1 0 $X=128950 $Y=47840
X808 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 50800 0 0 $X=128950 $Y=50560
X809 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 56240 1 0 $X=128950 $Y=53280
X810 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=129140 56240 0 0 $X=128950 $Y=56000
X811 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=132820 18160 1 0 $X=132630 $Y=15200
X812 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 12720 1 0 $X=143670 $Y=9760
X813 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 34480 1 0 $X=143670 $Y=31520
X814 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 34480 0 0 $X=143670 $Y=34240
X815 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 39920 1 0 $X=143670 $Y=36960
X816 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 39920 0 0 $X=143670 $Y=39680
X817 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 45360 1 0 $X=143670 $Y=42400
X818 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 45360 0 0 $X=143670 $Y=45120
X819 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 50800 1 0 $X=143670 $Y=47840
X820 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 50800 0 0 $X=143670 $Y=50560
X821 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 56240 1 0 $X=143670 $Y=53280
X822 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=143860 56240 0 0 $X=143670 $Y=56000
X823 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=145240 29040 1 0 $X=145050 $Y=26080
X824 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=150300 18160 1 0 $X=150110 $Y=15200
X825 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=150300 23600 1 0 $X=150110 $Y=20640
X826 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=153060 23600 0 0 $X=152870 $Y=23360
X827 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 12720 0 0 $X=158390 $Y=12480
X828 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 23600 0 0 $X=158390 $Y=23360
X829 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 29040 0 0 $X=158390 $Y=28800
X830 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 34480 1 0 $X=158390 $Y=31520
X831 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 34480 0 0 $X=158390 $Y=34240
X832 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 39920 1 0 $X=158390 $Y=36960
X833 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 39920 0 0 $X=158390 $Y=39680
X834 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 45360 1 0 $X=158390 $Y=42400
X835 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 45360 0 0 $X=158390 $Y=45120
X836 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 50800 1 0 $X=158390 $Y=47840
X837 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 50800 0 0 $X=158390 $Y=50560
X838 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 56240 1 0 $X=158390 $Y=53280
X839 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=158580 56240 0 0 $X=158390 $Y=56000
X840 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 23600 1 0 $X=173110 $Y=20640
X841 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 34480 1 0 $X=173110 $Y=31520
X842 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 34480 0 0 $X=173110 $Y=34240
X843 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 39920 1 0 $X=173110 $Y=36960
X844 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 39920 0 0 $X=173110 $Y=39680
X845 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 45360 1 0 $X=173110 $Y=42400
X846 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 45360 0 0 $X=173110 $Y=45120
X847 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 50800 1 0 $X=173110 $Y=47840
X848 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 50800 0 0 $X=173110 $Y=50560
X849 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 56240 1 0 $X=173110 $Y=53280
X850 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=173300 56240 0 0 $X=173110 $Y=56000
X851 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=174680 18160 0 0 $X=174490 $Y=17920
X852 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=174680 23600 0 0 $X=174490 $Y=23360
X853 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=176980 23600 0 0 $X=176790 $Y=23360
X854 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=185720 23600 0 0 $X=185530 $Y=23360
X855 1 2 2 1 sky130_fd_sc_hd__decap_4_DigitalLDOLogic_gds $T=187100 23600 1 0 $X=186910 $Y=20640
X856 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=44500 18160 0 0 $X=44310 $Y=17920
X857 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=44500 23600 0 0 $X=44310 $Y=23360
X858 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=44500 34480 0 0 $X=44310 $Y=34240
X859 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=55080 29040 1 0 $X=54890 $Y=26080
X860 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=55080 29040 0 0 $X=54890 $Y=28800
X861 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=59220 23600 0 0 $X=59030 $Y=23360
X862 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=84520 23600 0 0 $X=84330 $Y=23360
X863 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=88660 18160 0 0 $X=88470 $Y=17920
X864 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=88660 29040 0 0 $X=88470 $Y=28800
X865 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=96480 12720 0 0 $X=96290 $Y=12480
X866 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=108900 23600 0 0 $X=108710 $Y=23360
X867 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=118100 23600 1 0 $X=117910 $Y=20640
X868 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=125920 34480 1 0 $X=125730 $Y=31520
X869 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=127300 12720 0 0 $X=127110 $Y=12480
X870 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=128680 29040 0 0 $X=128490 $Y=28800
X871 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=132820 23600 0 0 $X=132630 $Y=23360
X872 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=132820 29040 0 0 $X=132630 $Y=28800
X873 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=142020 23600 1 0 $X=141830 $Y=20640
X874 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=153060 29040 1 0 $X=152870 $Y=26080
X875 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=153980 12720 1 0 $X=153790 $Y=9760
X876 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=168700 12720 1 0 $X=168510 $Y=9760
X877 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=171460 12720 0 0 $X=171270 $Y=12480
X878 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 12720 1 0 $X=182310 $Y=9760
X879 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 12720 0 0 $X=182310 $Y=12480
X880 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 18160 1 0 $X=182310 $Y=15200
X881 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 18160 0 0 $X=182310 $Y=17920
X882 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 29040 1 0 $X=182310 $Y=26080
X883 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 29040 0 0 $X=182310 $Y=28800
X884 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 34480 1 0 $X=182310 $Y=31520
X885 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 34480 0 0 $X=182310 $Y=34240
X886 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 39920 1 0 $X=182310 $Y=36960
X887 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 39920 0 0 $X=182310 $Y=39680
X888 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 45360 1 0 $X=182310 $Y=42400
X889 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 45360 0 0 $X=182310 $Y=45120
X890 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 50800 1 0 $X=182310 $Y=47840
X891 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 50800 0 0 $X=182310 $Y=50560
X892 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 56240 1 0 $X=182310 $Y=53280
X893 1 2 2 1 sky130_fd_sc_hd__decap_8_DigitalLDOLogic_gds $T=182500 56240 0 0 $X=182310 $Y=56000
X894 1 2 2 1 sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds $T=35300 18160 1 0 $X=35110 $Y=15200
X895 1 2 2 1 sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds $T=96940 12720 1 0 $X=96750 $Y=9760
X896 1 2 2 1 sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds $T=131900 23600 1 0 $X=131710 $Y=20640
X897 1 2 2 1 sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds $T=131900 29040 1 0 $X=131710 $Y=26080
X898 1 2 2 1 sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds $T=132820 23600 1 0 $X=132630 $Y=20640
X899 1 2 2 1 sky130_fd_sc_hd__fill_1_DigitalLDOLogic_gds $T=169620 23600 1 0 $X=169430 $Y=20640
X900 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=44500 12720 0 0 $X=44310 $Y=12480
X901 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=59220 23600 1 0 $X=59030 $Y=20640
X902 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=72560 12720 0 0 $X=72370 $Y=12480
X903 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=72560 23600 0 0 $X=72370 $Y=23360
X904 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=90040 23600 0 0 $X=89850 $Y=23360
X905 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=110280 18160 1 0 $X=110090 $Y=15200
X906 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=118100 34480 1 0 $X=117910 $Y=31520
X907 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=134200 29040 1 0 $X=134010 $Y=26080
X908 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=138340 12720 0 0 $X=138150 $Y=12480
X909 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=141560 18160 0 0 $X=141370 $Y=17920
X910 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=146160 12720 0 0 $X=145970 $Y=12480
X911 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=146160 18160 1 0 $X=145970 $Y=15200
X912 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=146160 18160 0 0 $X=145970 $Y=17920
X913 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=147540 12720 1 0 $X=147350 $Y=9760
X914 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=160880 18160 1 0 $X=160690 $Y=15200
X915 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=160880 23600 1 0 $X=160690 $Y=20640
X916 1 2 2 1 sky130_fd_sc_hd__fill_2_DigitalLDOLogic_gds $T=162260 12720 1 0 $X=162070 $Y=9760
X917 84 L1M1_PR_DigitalLDOLogic_gds $T=20350 13910 0 0 $X=20205 $Y=13795
X918 85 L1M1_PR_DigitalLDOLogic_gds $T=20350 16970 0 0 $X=20205 $Y=16855
X919 3 L1M1_PR_DigitalLDOLogic_gds $T=21270 14250 0 0 $X=21125 $Y=14135
X920 4 L1M1_PR_DigitalLDOLogic_gds $T=21270 16630 0 0 $X=21125 $Y=16515
X921 86 L1M1_PR_DigitalLDOLogic_gds $T=22190 24790 0 0 $X=22045 $Y=24675
X922 5 L1M1_PR_DigitalLDOLogic_gds $T=23110 25130 0 0 $X=22965 $Y=25015
X923 87 L1M1_PR_DigitalLDOLogic_gds $T=30930 11530 0 0 $X=30785 $Y=11415
X924 88 L1M1_PR_DigitalLDOLogic_gds $T=30930 16970 0 0 $X=30785 $Y=16855
X925 6 L1M1_PR_DigitalLDOLogic_gds $T=31850 11190 0 0 $X=31705 $Y=11075
X926 7 L1M1_PR_DigitalLDOLogic_gds $T=31850 16630 0 0 $X=31705 $Y=16515
X927 8 L1M1_PR_DigitalLDOLogic_gds $T=35070 14250 0 0 $X=34925 $Y=14135
X928 10 L1M1_PR_DigitalLDOLogic_gds $T=37830 13910 0 0 $X=37685 $Y=13795
X929 9 L1M1_PR_DigitalLDOLogic_gds $T=37830 27510 0 0 $X=37685 $Y=27395
X930 11 L1M1_PR_DigitalLDOLogic_gds $T=39210 16630 0 0 $X=39065 $Y=16515
X931 90 L1M1_PR_DigitalLDOLogic_gds $T=40590 16970 0 0 $X=40445 $Y=16855
X932 89 L1M1_PR_DigitalLDOLogic_gds $T=40590 27850 0 0 $X=40445 $Y=27735
X933 79 L1M1_PR_DigitalLDOLogic_gds $T=44730 16970 0 0 $X=44585 $Y=16855
X934 78 L1M1_PR_DigitalLDOLogic_gds $T=45420 16970 0 0 $X=45275 $Y=16855
X935 79 L1M1_PR_DigitalLDOLogic_gds $T=45650 14930 0 0 $X=45505 $Y=14815
X936 87 L1M1_PR_DigitalLDOLogic_gds $T=45675 13910 0 0 $X=45530 $Y=13795
X937 78 L1M1_PR_DigitalLDOLogic_gds $T=46110 13910 0 0 $X=45965 $Y=13795
X938 84 L1M1_PR_DigitalLDOLogic_gds $T=46110 17310 0 0 $X=45965 $Y=17195
X939 79 L1M1_PR_DigitalLDOLogic_gds $T=46110 22410 0 0 $X=45965 $Y=22295
X940 79 L1M1_PR_DigitalLDOLogic_gds $T=46110 27850 0 0 $X=45965 $Y=27735
X941 79 L1M1_PR_DigitalLDOLogic_gds $T=46110 30230 0 0 $X=45965 $Y=30115
X942 10 L1M1_PR_DigitalLDOLogic_gds $T=46570 16970 0 0 $X=46425 $Y=16855
X943 78 L1M1_PR_DigitalLDOLogic_gds $T=46800 22410 0 0 $X=46655 $Y=22295
X944 78 L1M1_PR_DigitalLDOLogic_gds $T=46800 27850 0 0 $X=46655 $Y=27735
X945 78 L1M1_PR_DigitalLDOLogic_gds $T=46800 30230 0 0 $X=46655 $Y=30115
X946 145 L1M1_PR_DigitalLDOLogic_gds $T=47260 16970 0 0 $X=47115 $Y=16855
X947 86 L1M1_PR_DigitalLDOLogic_gds $T=47260 27850 0 0 $X=47115 $Y=27735
X948 118 L1M1_PR_DigitalLDOLogic_gds $T=47490 14930 0 0 $X=47345 $Y=14815
X949 85 L1M1_PR_DigitalLDOLogic_gds $T=47490 22750 0 0 $X=47345 $Y=22635
X950 88 L1M1_PR_DigitalLDOLogic_gds $T=47490 30230 0 0 $X=47345 $Y=30115
X951 116 L1M1_PR_DigitalLDOLogic_gds $T=47950 17650 0 0 $X=47805 $Y=17535
X952 88 L1M1_PR_DigitalLDOLogic_gds $T=47950 22410 0 0 $X=47805 $Y=22295
X953 89 L1M1_PR_DigitalLDOLogic_gds $T=47950 28190 0 0 $X=47805 $Y=28075
X954 90 L1M1_PR_DigitalLDOLogic_gds $T=47950 29890 0 0 $X=47805 $Y=29775
X955 80 L1M1_PR_DigitalLDOLogic_gds $T=48410 36010 0 0 $X=48265 $Y=35895
X956 145 L1M1_PR_DigitalLDOLogic_gds $T=48640 22410 0 0 $X=48495 $Y=22295
X957 145 L1M1_PR_DigitalLDOLogic_gds $T=48640 27850 0 0 $X=48495 $Y=27735
X958 145 L1M1_PR_DigitalLDOLogic_gds $T=48640 30230 0 0 $X=48495 $Y=30115
X959 91 L1M1_PR_DigitalLDOLogic_gds $T=48870 11530 0 0 $X=48725 $Y=11415
X960 80 L1M1_PR_DigitalLDOLogic_gds $T=48870 32950 0 0 $X=48725 $Y=32835
X961 117 L1M1_PR_DigitalLDOLogic_gds $T=49330 23090 0 0 $X=49185 $Y=22975
X962 114 L1M1_PR_DigitalLDOLogic_gds $T=49330 28530 0 0 $X=49185 $Y=28415
X963 115 L1M1_PR_DigitalLDOLogic_gds $T=49330 31250 0 0 $X=49185 $Y=31135
X964 12 L1M1_PR_DigitalLDOLogic_gds $T=49715 11190 0 0 $X=49570 $Y=11075
X965 114 L1M1_PR_DigitalLDOLogic_gds $T=49715 35330 0 0 $X=49570 $Y=35215
X966 80 L1M1_PR_DigitalLDOLogic_gds $T=49790 19350 0 0 $X=49645 $Y=19235
X967 80 L1M1_PR_DigitalLDOLogic_gds $T=49790 24790 0 0 $X=49645 $Y=24675
X968 115 L1M1_PR_DigitalLDOLogic_gds $T=50175 33290 0 0 $X=50030 $Y=33175
X969 80 L1M1_PR_DigitalLDOLogic_gds $T=50250 16970 0 0 $X=50105 $Y=16855
X970 79 L1M1_PR_DigitalLDOLogic_gds $T=50740 13910 0 0 $X=50595 $Y=13795
X971 116 L1M1_PR_DigitalLDOLogic_gds $T=51095 19010 0 0 $X=50950 $Y=18895
X972 117 L1M1_PR_DigitalLDOLogic_gds $T=51095 24450 0 0 $X=50950 $Y=24335
X973 78 L1M1_PR_DigitalLDOLogic_gds $T=51175 13910 0 0 $X=51030 $Y=13795
X974 118 L1M1_PR_DigitalLDOLogic_gds $T=51555 16970 0 0 $X=51410 $Y=16855
X975 81 L1M1_PR_DigitalLDOLogic_gds $T=51630 22410 0 0 $X=51485 $Y=22295
X976 87 L1M1_PR_DigitalLDOLogic_gds $T=52090 13570 0 0 $X=51945 $Y=13455
X977 91 L1M1_PR_DigitalLDOLogic_gds $T=52550 13570 0 0 $X=52405 $Y=13455
X978 119 L1M1_PR_DigitalLDOLogic_gds $T=52935 22750 0 0 $X=52790 $Y=22635
X979 145 L1M1_PR_DigitalLDOLogic_gds $T=53240 13910 0 0 $X=53095 $Y=13795
X980 121 L1M1_PR_DigitalLDOLogic_gds $T=53930 14930 0 0 $X=53785 $Y=14815
X981 88 L1M1_PR_DigitalLDOLogic_gds $T=55310 34990 0 0 $X=55165 $Y=34875
X982 89 L1M1_PR_DigitalLDOLogic_gds $T=55770 32270 0 0 $X=55625 $Y=32155
X983 87 L1M1_PR_DigitalLDOLogic_gds $T=56690 18670 0 0 $X=56545 $Y=18555
X984 86 L1M1_PR_DigitalLDOLogic_gds $T=56690 24110 0 0 $X=56545 $Y=23995
X985 84 L1M1_PR_DigitalLDOLogic_gds $T=57150 15950 0 0 $X=57005 $Y=15835
X986 92 L1M1_PR_DigitalLDOLogic_gds $T=58530 21390 0 0 $X=58385 $Y=21275
X987 80 L1M1_PR_DigitalLDOLogic_gds $T=59450 16970 0 0 $X=59305 $Y=16855
X988 80 L1M1_PR_DigitalLDOLogic_gds $T=59450 19350 0 0 $X=59305 $Y=19235
X989 80 L1M1_PR_DigitalLDOLogic_gds $T=59450 27850 0 0 $X=59305 $Y=27735
X990 80 L1M1_PR_DigitalLDOLogic_gds $T=59450 30230 0 0 $X=59305 $Y=30115
X991 80 L1M1_PR_DigitalLDOLogic_gds $T=60370 23090 0 0 $X=60225 $Y=22975
X992 120 L1M1_PR_DigitalLDOLogic_gds $T=60755 16970 0 0 $X=60610 $Y=16855
X993 121 L1M1_PR_DigitalLDOLogic_gds $T=60755 19010 0 0 $X=60610 $Y=18895
X994 122 L1M1_PR_DigitalLDOLogic_gds $T=60755 27850 0 0 $X=60610 $Y=27735
X995 123 L1M1_PR_DigitalLDOLogic_gds $T=60755 29890 0 0 $X=60610 $Y=29775
X996 120 L1M1_PR_DigitalLDOLogic_gds $T=60830 14930 0 0 $X=60685 $Y=14815
X997 14 L1M1_PR_DigitalLDOLogic_gds $T=61290 22410 0 0 $X=61145 $Y=22295
X998 145 L1M1_PR_DigitalLDOLogic_gds $T=61520 13910 0 0 $X=61375 $Y=13795
X999 92 L1M1_PR_DigitalLDOLogic_gds $T=62210 13570 0 0 $X=62065 $Y=13455
X1000 92 L1M1_PR_DigitalLDOLogic_gds $T=62670 11530 0 0 $X=62525 $Y=11415
X1001 10 L1M1_PR_DigitalLDOLogic_gds $T=62670 13910 0 0 $X=62525 $Y=13795
X1002 78 L1M1_PR_DigitalLDOLogic_gds $T=63360 13910 0 0 $X=63215 $Y=13795
X1003 79 L1M1_PR_DigitalLDOLogic_gds $T=64050 13910 0 0 $X=63905 $Y=13795
X1004 15 L1M1_PR_DigitalLDOLogic_gds $T=65430 11190 0 0 $X=65285 $Y=11075
X1005 94 L1M1_PR_DigitalLDOLogic_gds $T=65890 24790 0 0 $X=65745 $Y=24675
X1006 91 L1M1_PR_DigitalLDOLogic_gds $T=66350 15950 0 0 $X=66205 $Y=15835
X1007 10 L1M1_PR_DigitalLDOLogic_gds $T=66350 18670 0 0 $X=66205 $Y=18555
X1008 81 L1M1_PR_DigitalLDOLogic_gds $T=66350 22410 0 0 $X=66205 $Y=22295
X1009 94 L1M1_PR_DigitalLDOLogic_gds $T=66350 26830 0 0 $X=66205 $Y=26715
X1010 90 L1M1_PR_DigitalLDOLogic_gds $T=66350 31250 0 0 $X=66205 $Y=31135
X1011 93 L1M1_PR_DigitalLDOLogic_gds $T=66810 13910 0 0 $X=66665 $Y=13795
X1012 124 L1M1_PR_DigitalLDOLogic_gds $T=67655 22410 0 0 $X=67510 $Y=22295
X1013 16 L1M1_PR_DigitalLDOLogic_gds $T=68190 14250 0 0 $X=68045 $Y=14135
X1014 122 L1M1_PR_DigitalLDOLogic_gds $T=68650 17650 0 0 $X=68505 $Y=17535
X1015 119 L1M1_PR_DigitalLDOLogic_gds $T=68650 20370 0 0 $X=68505 $Y=20255
X1016 123 L1M1_PR_DigitalLDOLogic_gds $T=68650 28530 0 0 $X=68505 $Y=28415
X1017 145 L1M1_PR_DigitalLDOLogic_gds $T=69340 16970 0 0 $X=69195 $Y=16855
X1018 145 L1M1_PR_DigitalLDOLogic_gds $T=69340 19350 0 0 $X=69195 $Y=19235
X1019 145 L1M1_PR_DigitalLDOLogic_gds $T=69340 27850 0 0 $X=69195 $Y=27735
X1020 93 L1M1_PR_DigitalLDOLogic_gds $T=70030 16970 0 0 $X=69885 $Y=16855
X1021 95 L1M1_PR_DigitalLDOLogic_gds $T=70030 19010 0 0 $X=69885 $Y=18895
X1022 13 L1M1_PR_DigitalLDOLogic_gds $T=70030 24450 0 0 $X=69885 $Y=24335
X1023 94 L1M1_PR_DigitalLDOLogic_gds $T=70030 27850 0 0 $X=69885 $Y=27735
X1024 90 L1M1_PR_DigitalLDOLogic_gds $T=70490 17310 0 0 $X=70345 $Y=17195
X1025 91 L1M1_PR_DigitalLDOLogic_gds $T=70490 19350 0 0 $X=70345 $Y=19235
X1026 89 L1M1_PR_DigitalLDOLogic_gds $T=70490 28190 0 0 $X=70345 $Y=28075
X1027 78 L1M1_PR_DigitalLDOLogic_gds $T=71180 27850 0 0 $X=71035 $Y=27735
X1028 78 L1M1_PR_DigitalLDOLogic_gds $T=71265 16970 0 0 $X=71120 $Y=16855
X1029 78 L1M1_PR_DigitalLDOLogic_gds $T=71265 19350 0 0 $X=71120 $Y=19235
X1030 79 L1M1_PR_DigitalLDOLogic_gds $T=71835 16970 0 0 $X=71690 $Y=16855
X1031 79 L1M1_PR_DigitalLDOLogic_gds $T=71870 19350 0 0 $X=71725 $Y=19235
X1032 79 L1M1_PR_DigitalLDOLogic_gds $T=71870 27850 0 0 $X=71725 $Y=27735
X1033 18 L1M1_PR_DigitalLDOLogic_gds $T=73250 23090 0 0 $X=73105 $Y=22975
X1034 18 L1M1_PR_DigitalLDOLogic_gds $T=74170 11530 0 0 $X=74025 $Y=11415
X1035 95 L1M1_PR_DigitalLDOLogic_gds $T=74170 16970 0 0 $X=74025 $Y=16855
X1036 79 L1M1_PR_DigitalLDOLogic_gds $T=74170 30230 0 0 $X=74025 $Y=30115
X1037 78 L1M1_PR_DigitalLDOLogic_gds $T=74860 30230 0 0 $X=74715 $Y=30115
X1038 81 L1M1_PR_DigitalLDOLogic_gds $T=75550 19350 0 0 $X=75405 $Y=19235
X1039 94 L1M1_PR_DigitalLDOLogic_gds $T=75550 29890 0 0 $X=75405 $Y=29775
X1040 18 L1M1_PR_DigitalLDOLogic_gds $T=76010 29890 0 0 $X=75865 $Y=29775
X1041 17 L1M1_PR_DigitalLDOLogic_gds $T=76470 16630 0 0 $X=76325 $Y=16515
X1042 145 L1M1_PR_DigitalLDOLogic_gds $T=76700 30230 0 0 $X=76555 $Y=30115
X1043 125 L1M1_PR_DigitalLDOLogic_gds $T=76855 19010 0 0 $X=76710 $Y=18895
X1044 81 L1M1_PR_DigitalLDOLogic_gds $T=77390 25130 0 0 $X=77245 $Y=25015
X1045 126 L1M1_PR_DigitalLDOLogic_gds $T=77390 29550 0 0 $X=77245 $Y=29435
X1046 19 L1M1_PR_DigitalLDOLogic_gds $T=78310 11190 0 0 $X=78165 $Y=11075
X1047 126 L1M1_PR_DigitalLDOLogic_gds $T=78695 24450 0 0 $X=78550 $Y=24335
X1048 14 L1M1_PR_DigitalLDOLogic_gds $T=79690 22410 0 0 $X=79545 $Y=22295
X1049 81 L1M1_PR_DigitalLDOLogic_gds $T=80610 23090 0 0 $X=80465 $Y=22975
X1050 79 L1M1_PR_DigitalLDOLogic_gds $T=80610 30230 0 0 $X=80465 $Y=30115
X1051 81 L1M1_PR_DigitalLDOLogic_gds $T=81070 22410 0 0 $X=80925 $Y=22295
X1052 78 L1M1_PR_DigitalLDOLogic_gds $T=81300 30230 0 0 $X=81155 $Y=30115
X1053 125 L1M1_PR_DigitalLDOLogic_gds $T=81530 17650 0 0 $X=81385 $Y=17535
X1054 18 L1M1_PR_DigitalLDOLogic_gds $T=81990 29830 0 0 $X=81845 $Y=29715
X1055 145 L1M1_PR_DigitalLDOLogic_gds $T=82220 16970 0 0 $X=82075 $Y=16855
X1056 127 L1M1_PR_DigitalLDOLogic_gds $T=82405 22750 0 0 $X=82260 $Y=22635
X1057 95 L1M1_PR_DigitalLDOLogic_gds $T=82450 18670 0 0 $X=82305 $Y=18555
X1058 98 L1M1_PR_DigitalLDOLogic_gds $T=82490 29890 0 0 $X=82345 $Y=29775
X1059 96 L1M1_PR_DigitalLDOLogic_gds $T=82910 11530 0 0 $X=82765 $Y=11415
X1060 96 L1M1_PR_DigitalLDOLogic_gds $T=82910 16970 0 0 $X=82765 $Y=16855
X1061 79 L1M1_PR_DigitalLDOLogic_gds $T=82910 19350 0 0 $X=82765 $Y=19235
X1062 145 L1M1_PR_DigitalLDOLogic_gds $T=83140 30230 0 0 $X=82995 $Y=30115
X1063 92 L1M1_PR_DigitalLDOLogic_gds $T=83370 16970 0 0 $X=83225 $Y=16855
X1064 78 L1M1_PR_DigitalLDOLogic_gds $T=83600 19350 0 0 $X=83455 $Y=19235
X1065 127 L1M1_PR_DigitalLDOLogic_gds $T=83830 29550 0 0 $X=83685 $Y=29435
X1066 78 L1M1_PR_DigitalLDOLogic_gds $T=84060 16970 0 0 $X=83915 $Y=16855
X1067 93 L1M1_PR_DigitalLDOLogic_gds $T=84290 19010 0 0 $X=84145 $Y=18895
X1068 93 L1M1_PR_DigitalLDOLogic_gds $T=84290 24110 0 0 $X=84145 $Y=23995
X1069 79 L1M1_PR_DigitalLDOLogic_gds $T=84750 16970 0 0 $X=84605 $Y=16855
X1070 97 L1M1_PR_DigitalLDOLogic_gds $T=84750 19350 0 0 $X=84605 $Y=19235
X1071 145 L1M1_PR_DigitalLDOLogic_gds $T=85440 19350 0 0 $X=85295 $Y=19235
X1072 124 L1M1_PR_DigitalLDOLogic_gds $T=86130 20370 0 0 $X=85985 $Y=20255
X1073 21 L1M1_PR_DigitalLDOLogic_gds $T=87050 11190 0 0 $X=86905 $Y=11075
X1074 97 L1M1_PR_DigitalLDOLogic_gds $T=87970 21390 0 0 $X=87825 $Y=21275
X1075 81 L1M1_PR_DigitalLDOLogic_gds $T=91190 24790 0 0 $X=91045 $Y=24675
X1076 97 L1M1_PR_DigitalLDOLogic_gds $T=91650 11530 0 0 $X=91505 $Y=11415
X1077 128 L1M1_PR_DigitalLDOLogic_gds $T=92495 24450 0 0 $X=92350 $Y=24335
X1078 79 L1M1_PR_DigitalLDOLogic_gds $T=93030 13910 0 0 $X=92885 $Y=13795
X1079 20 L1M1_PR_DigitalLDOLogic_gds $T=93490 11190 0 0 $X=93345 $Y=11075
X1080 78 L1M1_PR_DigitalLDOLogic_gds $T=93720 13910 0 0 $X=93575 $Y=13795
X1081 81 L1M1_PR_DigitalLDOLogic_gds $T=93950 19690 0 0 $X=93805 $Y=19575
X1082 79 L1M1_PR_DigitalLDOLogic_gds $T=93950 30230 0 0 $X=93805 $Y=30115
X1083 97 L1M1_PR_DigitalLDOLogic_gds $T=94410 13910 0 0 $X=94265 $Y=13795
X1084 78 L1M1_PR_DigitalLDOLogic_gds $T=94640 30230 0 0 $X=94495 $Y=30115
X1085 99 L1M1_PR_DigitalLDOLogic_gds $T=94870 13570 0 0 $X=94725 $Y=13455
X1086 129 L1M1_PR_DigitalLDOLogic_gds $T=94870 17650 0 0 $X=94725 $Y=17535
X1087 129 L1M1_PR_DigitalLDOLogic_gds $T=95255 19010 0 0 $X=95110 $Y=18895
X1088 96 L1M1_PR_DigitalLDOLogic_gds $T=95330 29890 0 0 $X=95185 $Y=29775
X1089 145 L1M1_PR_DigitalLDOLogic_gds $T=95560 13910 0 0 $X=95415 $Y=13795
X1090 145 L1M1_PR_DigitalLDOLogic_gds $T=95560 16970 0 0 $X=95415 $Y=16855
X1091 81 L1M1_PR_DigitalLDOLogic_gds $T=95790 22410 0 0 $X=95645 $Y=22295
X1092 101 L1M1_PR_DigitalLDOLogic_gds $T=95790 30230 0 0 $X=95645 $Y=30115
X1093 128 L1M1_PR_DigitalLDOLogic_gds $T=96245 13230 0 0 $X=96100 $Y=13115
X1094 100 L1M1_PR_DigitalLDOLogic_gds $T=96250 16970 0 0 $X=96105 $Y=16855
X1095 145 L1M1_PR_DigitalLDOLogic_gds $T=96480 30230 0 0 $X=96335 $Y=30115
X1096 95 L1M1_PR_DigitalLDOLogic_gds $T=96710 17310 0 0 $X=96565 $Y=17195
X1097 130 L1M1_PR_DigitalLDOLogic_gds $T=97095 22750 0 0 $X=96950 $Y=22635
X1098 130 L1M1_PR_DigitalLDOLogic_gds $T=97170 29550 0 0 $X=97025 $Y=29435
X1099 78 L1M1_PR_DigitalLDOLogic_gds $T=97485 16970 0 0 $X=97340 $Y=16855
X1100 79 L1M1_PR_DigitalLDOLogic_gds $T=98090 16970 0 0 $X=97945 $Y=16855
X1101 98 L1M1_PR_DigitalLDOLogic_gds $T=98090 24110 0 0 $X=97945 $Y=23995
X1102 98 L1M1_PR_DigitalLDOLogic_gds $T=98550 11530 0 0 $X=98405 $Y=11415
X1103 22 L1M1_PR_DigitalLDOLogic_gds $T=99470 11190 0 0 $X=99325 $Y=11075
X1104 96 L1M1_PR_DigitalLDOLogic_gds $T=100850 18670 0 0 $X=100705 $Y=18555
X1105 96 L1M1_PR_DigitalLDOLogic_gds $T=100850 20370 0 0 $X=100705 $Y=20255
X1106 100 L1M1_PR_DigitalLDOLogic_gds $T=102690 21390 0 0 $X=102545 $Y=21275
X1107 99 L1M1_PR_DigitalLDOLogic_gds $T=103610 13910 0 0 $X=103465 $Y=13795
X1108 100 L1M1_PR_DigitalLDOLogic_gds $T=103610 16970 0 0 $X=103465 $Y=16855
X1109 24 L1M1_PR_DigitalLDOLogic_gds $T=105450 14250 0 0 $X=105305 $Y=14135
X1110 23 L1M1_PR_DigitalLDOLogic_gds $T=105450 16630 0 0 $X=105305 $Y=16515
X1111 25 L1M1_PR_DigitalLDOLogic_gds $T=110510 19010 0 0 $X=110365 $Y=18895
X1112 82 L1M1_PR_DigitalLDOLogic_gds $T=110510 22410 0 0 $X=110365 $Y=22295
X1113 79 L1M1_PR_DigitalLDOLogic_gds $T=111430 16970 0 0 $X=111285 $Y=16855
X1114 131 L1M1_PR_DigitalLDOLogic_gds $T=111815 22750 0 0 $X=111670 $Y=22635
X1115 78 L1M1_PR_DigitalLDOLogic_gds $T=112120 16970 0 0 $X=111975 $Y=16855
X1116 100 L1M1_PR_DigitalLDOLogic_gds $T=112810 16970 0 0 $X=112665 $Y=16855
X1117 79 L1M1_PR_DigitalLDOLogic_gds $T=112810 24790 0 0 $X=112665 $Y=24675
X1118 104 L1M1_PR_DigitalLDOLogic_gds $T=113270 17310 0 0 $X=113125 $Y=17195
X1119 78 L1M1_PR_DigitalLDOLogic_gds $T=113500 24790 0 0 $X=113355 $Y=24675
X1120 26 L1M1_PR_DigitalLDOLogic_gds $T=113730 14250 0 0 $X=113585 $Y=14135
X1121 145 L1M1_PR_DigitalLDOLogic_gds $T=113960 16970 0 0 $X=113815 $Y=16855
X1122 113 L1M1_PR_DigitalLDOLogic_gds $T=114190 24450 0 0 $X=114045 $Y=24335
X1123 131 L1M1_PR_DigitalLDOLogic_gds $T=114650 17650 0 0 $X=114505 $Y=17535
X1124 101 L1M1_PR_DigitalLDOLogic_gds $T=114650 19350 0 0 $X=114505 $Y=19235
X1125 86 L1M1_PR_DigitalLDOLogic_gds $T=114650 24790 0 0 $X=114505 $Y=24675
X1126 145 L1M1_PR_DigitalLDOLogic_gds $T=115340 24790 0 0 $X=115195 $Y=24675
X1127 102 L1M1_PR_DigitalLDOLogic_gds $T=115570 13910 0 0 $X=115425 $Y=13795
X1128 133 L1M1_PR_DigitalLDOLogic_gds $T=116030 24110 0 0 $X=115885 $Y=23995
X1129 101 L1M1_PR_DigitalLDOLogic_gds $T=117410 21390 0 0 $X=117265 $Y=21275
X1130 79 L1M1_PR_DigitalLDOLogic_gds $T=118330 13910 0 0 $X=118185 $Y=13795
X1131 82 L1M1_PR_DigitalLDOLogic_gds $T=118330 19690 0 0 $X=118185 $Y=19575
X1132 82 L1M1_PR_DigitalLDOLogic_gds $T=118330 24790 0 0 $X=118185 $Y=24675
X1133 78 L1M1_PR_DigitalLDOLogic_gds $T=119070 13910 0 0 $X=118925 $Y=13795
X1134 98 L1M1_PR_DigitalLDOLogic_gds $T=119635 13570 0 0 $X=119490 $Y=13455
X1135 132 L1M1_PR_DigitalLDOLogic_gds $T=119635 19010 0 0 $X=119490 $Y=18895
X1136 133 L1M1_PR_DigitalLDOLogic_gds $T=119635 24450 0 0 $X=119490 $Y=24335
X1137 145 L1M1_PR_DigitalLDOLogic_gds $T=119635 32270 0 0 $X=119490 $Y=32155
X1138 79 L1M1_PR_DigitalLDOLogic_gds $T=119710 27850 0 0 $X=119565 $Y=27735
X1139 79 L1M1_PR_DigitalLDOLogic_gds $T=119710 30230 0 0 $X=119565 $Y=30115
X1140 102 L1M1_PR_DigitalLDOLogic_gds $T=120170 13570 0 0 $X=120025 $Y=13455
X1141 29 L1M1_PR_DigitalLDOLogic_gds $T=120170 33290 0 0 $X=120025 $Y=33175
X1142 78 L1M1_PR_DigitalLDOLogic_gds $T=120400 27850 0 0 $X=120255 $Y=27735
X1143 78 L1M1_PR_DigitalLDOLogic_gds $T=120400 30230 0 0 $X=120255 $Y=30115
X1144 28 L1M1_PR_DigitalLDOLogic_gds $T=120630 16630 0 0 $X=120485 $Y=16515
X1145 145 L1M1_PR_DigitalLDOLogic_gds $T=120910 13910 0 0 $X=120765 $Y=13795
X1146 112 L1M1_PR_DigitalLDOLogic_gds $T=121090 27850 0 0 $X=120945 $Y=27735
X1147 101 L1M1_PR_DigitalLDOLogic_gds $T=121090 29890 0 0 $X=120945 $Y=29775
X1148 27 L1M1_PR_DigitalLDOLogic_gds $T=121550 11190 0 0 $X=121405 $Y=11075
X1149 132 L1M1_PR_DigitalLDOLogic_gds $T=121550 13230 0 0 $X=121405 $Y=13115
X1150 85 L1M1_PR_DigitalLDOLogic_gds $T=121550 28190 0 0 $X=121405 $Y=28075
X1151 106 L1M1_PR_DigitalLDOLogic_gds $T=121550 29890 0 0 $X=121405 $Y=29775
X1152 145 L1M1_PR_DigitalLDOLogic_gds $T=122240 27850 0 0 $X=122095 $Y=27735
X1153 145 L1M1_PR_DigitalLDOLogic_gds $T=122240 30230 0 0 $X=122095 $Y=30115
X1154 104 L1M1_PR_DigitalLDOLogic_gds $T=122470 16970 0 0 $X=122325 $Y=16855
X1155 103 L1M1_PR_DigitalLDOLogic_gds $T=122930 11530 0 0 $X=122785 $Y=11415
X1156 135 L1M1_PR_DigitalLDOLogic_gds $T=122930 28530 0 0 $X=122785 $Y=28415
X1157 134 L1M1_PR_DigitalLDOLogic_gds $T=122930 29550 0 0 $X=122785 $Y=29435
X1158 82 L1M1_PR_DigitalLDOLogic_gds $T=124770 22410 0 0 $X=124625 $Y=22295
X1159 82 L1M1_PR_DigitalLDOLogic_gds $T=124770 27510 0 0 $X=124625 $Y=27395
X1160 99 L1M1_PR_DigitalLDOLogic_gds $T=125230 18670 0 0 $X=125085 $Y=18555
X1161 85 L1M1_PR_DigitalLDOLogic_gds $T=125230 25810 0 0 $X=125085 $Y=25695
X1162 79 L1M1_PR_DigitalLDOLogic_gds $T=125690 16970 0 0 $X=125545 $Y=16855
X1163 134 L1M1_PR_DigitalLDOLogic_gds $T=126075 22750 0 0 $X=125930 $Y=22635
X1164 135 L1M1_PR_DigitalLDOLogic_gds $T=126075 28190 0 0 $X=125930 $Y=28075
X1165 78 L1M1_PR_DigitalLDOLogic_gds $T=126290 16970 0 0 $X=126145 $Y=16855
X1166 99 L1M1_PR_DigitalLDOLogic_gds $T=127070 17310 0 0 $X=126925 $Y=17195
X1167 103 L1M1_PR_DigitalLDOLogic_gds $T=127530 16970 0 0 $X=127385 $Y=16855
X1168 145 L1M1_PR_DigitalLDOLogic_gds $T=128220 16970 0 0 $X=128075 $Y=16855
X1169 136 L1M1_PR_DigitalLDOLogic_gds $T=128910 17650 0 0 $X=128765 $Y=17535
X1170 104 L1M1_PR_DigitalLDOLogic_gds $T=131670 21390 0 0 $X=131525 $Y=21275
X1171 113 L1M1_PR_DigitalLDOLogic_gds $T=131670 26830 0 0 $X=131525 $Y=26715
X1172 113 L1M1_PR_DigitalLDOLogic_gds $T=131670 28530 0 0 $X=131525 $Y=28415
X1173 82 L1M1_PR_DigitalLDOLogic_gds $T=133050 19690 0 0 $X=132905 $Y=19575
X1174 14 L1M1_PR_DigitalLDOLogic_gds $T=133510 22410 0 0 $X=133365 $Y=22295
X1175 105 L1M1_PR_DigitalLDOLogic_gds $T=133970 13910 0 0 $X=133825 $Y=13795
X1176 136 L1M1_PR_DigitalLDOLogic_gds $T=134355 19350 0 0 $X=134210 $Y=19235
X1177 82 L1M1_PR_DigitalLDOLogic_gds $T=134430 23090 0 0 $X=134285 $Y=22975
X1178 30 L1M1_PR_DigitalLDOLogic_gds $T=134890 14250 0 0 $X=134745 $Y=14135
X1179 79 L1M1_PR_DigitalLDOLogic_gds $T=134890 16970 0 0 $X=134745 $Y=16855
X1180 82 L1M1_PR_DigitalLDOLogic_gds $T=134890 22410 0 0 $X=134745 $Y=22295
X1181 82 L1M1_PR_DigitalLDOLogic_gds $T=135350 27510 0 0 $X=135205 $Y=27395
X1182 78 L1M1_PR_DigitalLDOLogic_gds $T=135580 16970 0 0 $X=135435 $Y=16855
X1183 137 L1M1_PR_DigitalLDOLogic_gds $T=136195 22750 0 0 $X=136050 $Y=22635
X1184 102 L1M1_PR_DigitalLDOLogic_gds $T=136270 17310 0 0 $X=136125 $Y=17195
X1185 105 L1M1_PR_DigitalLDOLogic_gds $T=136655 16970 0 0 $X=136510 $Y=16855
X1186 138 L1M1_PR_DigitalLDOLogic_gds $T=136655 28190 0 0 $X=136510 $Y=28075
X1187 145 L1M1_PR_DigitalLDOLogic_gds $T=137420 16970 0 0 $X=137275 $Y=16855
X1188 140 L1M1_PR_DigitalLDOLogic_gds $T=138110 17650 0 0 $X=137965 $Y=17535
X1189 137 L1M1_PR_DigitalLDOLogic_gds $T=138110 24110 0 0 $X=137965 $Y=23995
X1190 138 L1M1_PR_DigitalLDOLogic_gds $T=138110 29550 0 0 $X=137965 $Y=29435
X1191 145 L1M1_PR_DigitalLDOLogic_gds $T=138800 24790 0 0 $X=138655 $Y=24675
X1192 145 L1M1_PR_DigitalLDOLogic_gds $T=138800 30230 0 0 $X=138655 $Y=30115
X1193 106 L1M1_PR_DigitalLDOLogic_gds $T=139490 11530 0 0 $X=139345 $Y=11415
X1194 108 L1M1_PR_DigitalLDOLogic_gds $T=139490 24450 0 0 $X=139345 $Y=24335
X1195 110 L1M1_PR_DigitalLDOLogic_gds $T=139490 30230 0 0 $X=139345 $Y=30115
X1196 102 L1M1_PR_DigitalLDOLogic_gds $T=139950 18670 0 0 $X=139805 $Y=18555
X1197 104 L1M1_PR_DigitalLDOLogic_gds $T=139950 24790 0 0 $X=139805 $Y=24675
X1198 106 L1M1_PR_DigitalLDOLogic_gds $T=139950 29890 0 0 $X=139805 $Y=29775
X1199 31 L1M1_PR_DigitalLDOLogic_gds $T=140410 11190 0 0 $X=140265 $Y=11075
X1200 78 L1M1_PR_DigitalLDOLogic_gds $T=140640 24790 0 0 $X=140495 $Y=24675
X1201 78 L1M1_PR_DigitalLDOLogic_gds $T=140640 30230 0 0 $X=140495 $Y=30115
X1202 79 L1M1_PR_DigitalLDOLogic_gds $T=141330 24790 0 0 $X=141185 $Y=24675
X1203 79 L1M1_PR_DigitalLDOLogic_gds $T=141330 30230 0 0 $X=141185 $Y=30115
X1204 106 L1M1_PR_DigitalLDOLogic_gds $T=141790 23090 0 0 $X=141645 $Y=22975
X1205 108 L1M1_PR_DigitalLDOLogic_gds $T=142250 26830 0 0 $X=142105 $Y=26715
X1206 32 L1M1_PR_DigitalLDOLogic_gds $T=142710 14250 0 0 $X=142565 $Y=14135
X1207 79 L1M1_PR_DigitalLDOLogic_gds $T=142710 16970 0 0 $X=142565 $Y=16855
X1208 79 L1M1_PR_DigitalLDOLogic_gds $T=142710 19350 0 0 $X=142565 $Y=19235
X1209 78 L1M1_PR_DigitalLDOLogic_gds $T=143175 16970 0 0 $X=143030 $Y=16855
X1210 78 L1M1_PR_DigitalLDOLogic_gds $T=143400 19350 0 0 $X=143255 $Y=19235
X1211 103 L1M1_PR_DigitalLDOLogic_gds $T=144090 16970 0 0 $X=143945 $Y=16855
X1212 105 L1M1_PR_DigitalLDOLogic_gds $T=144090 19350 0 0 $X=143945 $Y=19235
X1213 107 L1M1_PR_DigitalLDOLogic_gds $T=144550 13910 0 0 $X=144405 $Y=13795
X1214 109 L1M1_PR_DigitalLDOLogic_gds $T=144550 19350 0 0 $X=144405 $Y=19235
X1215 107 L1M1_PR_DigitalLDOLogic_gds $T=144695 16970 0 0 $X=144550 $Y=16855
X1216 145 L1M1_PR_DigitalLDOLogic_gds $T=145240 19350 0 0 $X=145095 $Y=19235
X1217 145 L1M1_PR_DigitalLDOLogic_gds $T=145290 16970 0 0 $X=145145 $Y=16855
X1218 139 L1M1_PR_DigitalLDOLogic_gds $T=145930 17650 0 0 $X=145785 $Y=17535
X1219 143 L1M1_PR_DigitalLDOLogic_gds $T=145930 18670 0 0 $X=145785 $Y=18555
X1220 109 L1M1_PR_DigitalLDOLogic_gds $T=148690 11530 0 0 $X=148545 $Y=11415
X1221 33 L1M1_PR_DigitalLDOLogic_gds $T=150990 25130 0 0 $X=150845 $Y=25015
X1222 108 L1M1_PR_DigitalLDOLogic_gds $T=151910 24790 0 0 $X=151765 $Y=24675
X1223 34 L1M1_PR_DigitalLDOLogic_gds $T=152830 11190 0 0 $X=152685 $Y=11075
X1224 83 L1M1_PR_DigitalLDOLogic_gds $T=153290 19350 0 0 $X=153145 $Y=19235
X1225 83 L1M1_PR_DigitalLDOLogic_gds $T=153750 16970 0 0 $X=153605 $Y=16855
X1226 83 L1M1_PR_DigitalLDOLogic_gds $T=153750 22070 0 0 $X=153605 $Y=21955
X1227 139 L1M1_PR_DigitalLDOLogic_gds $T=154595 19010 0 0 $X=154450 $Y=18895
X1228 140 L1M1_PR_DigitalLDOLogic_gds $T=155055 16970 0 0 $X=154910 $Y=16855
X1229 141 L1M1_PR_DigitalLDOLogic_gds $T=155055 22750 0 0 $X=154910 $Y=22635
X1230 141 L1M1_PR_DigitalLDOLogic_gds $T=155130 24110 0 0 $X=154985 $Y=23995
X1231 145 L1M1_PR_DigitalLDOLogic_gds $T=155820 24790 0 0 $X=155675 $Y=24675
X1232 112 L1M1_PR_DigitalLDOLogic_gds $T=156510 24450 0 0 $X=156365 $Y=24335
X1233 108 L1M1_PR_DigitalLDOLogic_gds $T=156970 24790 0 0 $X=156825 $Y=24675
X1234 79 L1M1_PR_DigitalLDOLogic_gds $T=156970 27850 0 0 $X=156825 $Y=27735
X1235 78 L1M1_PR_DigitalLDOLogic_gds $T=157660 24790 0 0 $X=157515 $Y=24675
X1236 78 L1M1_PR_DigitalLDOLogic_gds $T=157660 27850 0 0 $X=157515 $Y=27735
X1237 79 L1M1_PR_DigitalLDOLogic_gds $T=158350 24790 0 0 $X=158205 $Y=24675
X1238 110 L1M1_PR_DigitalLDOLogic_gds $T=158350 28190 0 0 $X=158205 $Y=28075
X1239 113 L1M1_PR_DigitalLDOLogic_gds $T=158810 28190 0 0 $X=158665 $Y=28075
X1240 145 L1M1_PR_DigitalLDOLogic_gds $T=159500 27850 0 0 $X=159355 $Y=27735
X1241 105 L1M1_PR_DigitalLDOLogic_gds $T=160190 20370 0 0 $X=160045 $Y=20255
X1242 142 L1M1_PR_DigitalLDOLogic_gds $T=160190 26830 0 0 $X=160045 $Y=26715
X1243 103 L1M1_PR_DigitalLDOLogic_gds $T=160650 15950 0 0 $X=160505 $Y=15835
X1244 110 L1M1_PR_DigitalLDOLogic_gds $T=160650 23090 0 0 $X=160505 $Y=22975
X1245 110 L1M1_PR_DigitalLDOLogic_gds $T=162490 16970 0 0 $X=162345 $Y=16855
X1246 77 L1M1_PR_DigitalLDOLogic_gds $T=162490 19350 0 0 $X=162345 $Y=19235
X1247 83 L1M1_PR_DigitalLDOLogic_gds $T=162490 22410 0 0 $X=162345 $Y=22295
X1248 142 L1M1_PR_DigitalLDOLogic_gds $T=163795 22750 0 0 $X=163650 $Y=22635
X1249 111 L1M1_PR_DigitalLDOLogic_gds $T=164330 11530 0 0 $X=164185 $Y=11415
X1250 36 L1M1_PR_DigitalLDOLogic_gds $T=164790 16630 0 0 $X=164645 $Y=16515
X1251 35 L1M1_PR_DigitalLDOLogic_gds $T=165250 11190 0 0 $X=165105 $Y=11075
X1252 76 L1M1_PR_DigitalLDOLogic_gds $T=165250 19010 0 0 $X=165105 $Y=18895
X1253 83 L1M1_PR_DigitalLDOLogic_gds $T=165710 19350 0 0 $X=165565 $Y=19235
X1254 76 L1M1_PR_DigitalLDOLogic_gds $T=167015 19010 0 0 $X=166870 $Y=18895
X1255 77 L1M1_PR_DigitalLDOLogic_gds $T=168010 14930 0 0 $X=167865 $Y=14815
X1256 145 L1M1_PR_DigitalLDOLogic_gds $T=168700 13910 0 0 $X=168555 $Y=13795
X1257 111 L1M1_PR_DigitalLDOLogic_gds $T=169390 13570 0 0 $X=169245 $Y=13455
X1258 83 L1M1_PR_DigitalLDOLogic_gds $T=169390 16970 0 0 $X=169245 $Y=16855
X1259 112 L1M1_PR_DigitalLDOLogic_gds $T=169390 21390 0 0 $X=169245 $Y=21275
X1260 112 L1M1_PR_DigitalLDOLogic_gds $T=169390 23090 0 0 $X=169245 $Y=22975
X1261 144 L1M1_PR_DigitalLDOLogic_gds $T=169390 24450 0 0 $X=169245 $Y=24335
X1262 107 L1M1_PR_DigitalLDOLogic_gds $T=169850 13910 0 0 $X=169705 $Y=13795
X1263 14 L1M1_PR_DigitalLDOLogic_gds $T=170310 22410 0 0 $X=170165 $Y=22295
X1264 79 L1M1_PR_DigitalLDOLogic_gds $T=170310 24790 0 0 $X=170165 $Y=24675
X1265 29 L1M1_PR_DigitalLDOLogic_gds $T=170540 13910 0 0 $X=170395 $Y=13795
X1266 143 L1M1_PR_DigitalLDOLogic_gds $T=170725 16970 0 0 $X=170580 $Y=16855
X1267 37 L1M1_PR_DigitalLDOLogic_gds $T=171230 13910 0 0 $X=171085 $Y=13795
X1268 83 L1M1_PR_DigitalLDOLogic_gds $T=171230 21730 0 0 $X=171085 $Y=21615
X1269 109 L1M1_PR_DigitalLDOLogic_gds $T=171230 24110 0 0 $X=171085 $Y=23995
X1270 78 L1M1_PR_DigitalLDOLogic_gds $T=171690 24790 0 0 $X=171545 $Y=24675
X1271 29 L1M1_PR_DigitalLDOLogic_gds $T=172150 22750 0 0 $X=172005 $Y=22635
X1272 109 L1M1_PR_DigitalLDOLogic_gds $T=172610 20030 0 0 $X=172465 $Y=19915
X1273 78 L1M1_PR_DigitalLDOLogic_gds $T=173070 22750 0 0 $X=172925 $Y=22635
X1274 37 L1M1_PR_DigitalLDOLogic_gds $T=173530 19350 0 0 $X=173385 $Y=19235
X1275 79 L1M1_PR_DigitalLDOLogic_gds $T=173990 20370 0 0 $X=173845 $Y=20255
X1276 107 L1M1_PR_DigitalLDOLogic_gds $T=176290 15950 0 0 $X=176145 $Y=15835
X1277 112 L1M1_PR_DigitalLDOLogic_gds $T=177210 16970 0 0 $X=177065 $Y=16855
X1278 83 L1M1_PR_DigitalLDOLogic_gds $T=177210 22070 0 0 $X=177065 $Y=21955
X1279 144 L1M1_PR_DigitalLDOLogic_gds $T=178515 22750 0 0 $X=178370 $Y=22635
X1280 38 L1M1_PR_DigitalLDOLogic_gds $T=179050 16630 0 0 $X=178905 $Y=16515
X1281 113 L1M1_PR_DigitalLDOLogic_gds $T=181350 24790 0 0 $X=181205 $Y=24675
X1282 111 L1M1_PR_DigitalLDOLogic_gds $T=184110 21390 0 0 $X=183965 $Y=21275
X1283 39 L1M1_PR_DigitalLDOLogic_gds $T=184570 24450 0 0 $X=184425 $Y=24335
X1284 78 M1M2_PR_M $T=43350 13570 0 0 $X=43190 $Y=13440
X1285 84 M1M2_PR_M $T=43350 14250 0 0 $X=43190 $Y=14120
X1286 79 M1M2_PR_M $T=43350 16290 0 0 $X=43190 $Y=16160
X1287 86 M1M2_PR_M $T=46110 24450 0 0 $X=45950 $Y=24320
X1288 87 M1M2_PR_M $T=48870 13570 0 0 $X=48710 $Y=13440
X1289 90 M1M2_PR_M $T=70950 17650 0 0 $X=70790 $Y=17520
X1290 79 M1M2_PR_M $T=109590 14590 0 0 $X=109430 $Y=14460
X1291 78 M1M2_PR_M $T=112350 27170 0 0 $X=112190 $Y=27040
X1292 79 M1M2_PR_M $T=128910 16290 0 0 $X=128750 $Y=16160
X1293 145 M1M2_PR_M $T=148230 16970 0 0 $X=148070 $Y=16840
X1294 4 M1M2_PR_DigitalLDOLogic_gds $T=10230 16630 0 0 $X=10070 $Y=16470
X1295 3 M1M2_PR_DigitalLDOLogic_gds $T=15750 14250 0 0 $X=15590 $Y=14090
X1296 5 M1M2_PR_DigitalLDOLogic_gds $T=18510 25130 0 0 $X=18350 $Y=24970
X1297 6 M1M2_PR_DigitalLDOLogic_gds $T=26790 11190 0 0 $X=26630 $Y=11030
X1298 7 M1M2_PR_DigitalLDOLogic_gds $T=29550 16630 0 0 $X=29390 $Y=16470
X1299 85 M1M2_PR_DigitalLDOLogic_gds $T=29550 17310 0 0 $X=29390 $Y=17150
X1300 85 M1M2_PR_DigitalLDOLogic_gds $T=29550 22750 0 0 $X=29390 $Y=22590
X1301 88 M1M2_PR_DigitalLDOLogic_gds $T=32310 17310 0 0 $X=32150 $Y=17150
X1302 88 M1M2_PR_DigitalLDOLogic_gds $T=32310 21390 0 0 $X=32150 $Y=21230
X1303 8 M1M2_PR_DigitalLDOLogic_gds $T=35070 14250 0 0 $X=34910 $Y=14090
X1304 84 M1M2_PR_DigitalLDOLogic_gds $T=35070 14930 0 0 $X=34910 $Y=14770
X1305 84 M1M2_PR_DigitalLDOLogic_gds $T=35070 17650 0 0 $X=34910 $Y=17490
X1306 9 M1M2_PR_DigitalLDOLogic_gds $T=37830 27510 0 0 $X=37670 $Y=27350
X1307 11 M1M2_PR_DigitalLDOLogic_gds $T=40590 650 0 0 $X=40430 $Y=490
X1308 11 M1M2_PR_DigitalLDOLogic_gds $T=40590 16290 0 0 $X=40430 $Y=16130
X1309 90 M1M2_PR_DigitalLDOLogic_gds $T=40590 16970 0 0 $X=40430 $Y=16810
X1310 85 M1M2_PR_DigitalLDOLogic_gds $T=40590 22750 0 0 $X=40430 $Y=22590
X1311 90 M1M2_PR_DigitalLDOLogic_gds $T=40590 29890 0 0 $X=40430 $Y=29730
X1312 85 M1M2_PR_DigitalLDOLogic_gds $T=40590 38390 0 0 $X=40430 $Y=38230
X1313 84 M1M2_PR_DigitalLDOLogic_gds $T=42890 9490 0 0 $X=42730 $Y=9330
X1314 79 M1M2_PR_DigitalLDOLogic_gds $T=43350 14930 0 0 $X=43190 $Y=14770
X1315 78 M1M2_PR_DigitalLDOLogic_gds $T=43350 17310 0 0 $X=43190 $Y=17150
X1316 78 M1M2_PR_DigitalLDOLogic_gds $T=43350 22070 0 0 $X=43190 $Y=21910
X1317 78 M1M2_PR_DigitalLDOLogic_gds $T=43350 27510 0 0 $X=43190 $Y=27350
X1318 78 M1M2_PR_DigitalLDOLogic_gds $T=43350 30570 0 0 $X=43190 $Y=30410
X1319 87 M1M2_PR_DigitalLDOLogic_gds $T=46110 11530 0 0 $X=45950 $Y=11370
X1320 10 M1M2_PR_DigitalLDOLogic_gds $T=46110 13230 0 0 $X=45950 $Y=13070
X1321 87 M1M2_PR_DigitalLDOLogic_gds $T=46110 14590 0 0 $X=45950 $Y=14430
X1322 10 M1M2_PR_DigitalLDOLogic_gds $T=46110 15950 0 0 $X=45950 $Y=15790
X1323 79 M1M2_PR_DigitalLDOLogic_gds $T=46110 16630 0 0 $X=45950 $Y=16470
X1324 79 M1M2_PR_DigitalLDOLogic_gds $T=46110 22410 0 0 $X=45950 $Y=22250
X1325 88 M1M2_PR_DigitalLDOLogic_gds $T=46110 23090 0 0 $X=45950 $Y=22930
X1326 86 M1M2_PR_DigitalLDOLogic_gds $T=46110 26830 0 0 $X=45950 $Y=26670
X1327 79 M1M2_PR_DigitalLDOLogic_gds $T=46110 27850 0 0 $X=45950 $Y=27690
X1328 79 M1M2_PR_DigitalLDOLogic_gds $T=46110 29550 0 0 $X=45950 $Y=29390
X1329 79 M1M2_PR_DigitalLDOLogic_gds $T=46110 30230 0 0 $X=45950 $Y=30070
X1330 88 M1M2_PR_DigitalLDOLogic_gds $T=46110 30910 0 0 $X=45950 $Y=30750
X1331 11 M1M2_PR_DigitalLDOLogic_gds $T=48410 650 0 0 $X=48250 $Y=490
X1332 84 M1M2_PR_DigitalLDOLogic_gds $T=48410 9490 0 0 $X=48250 $Y=9330
X1333 87 M1M2_PR_DigitalLDOLogic_gds $T=48525 14590 0 0 $X=48365 $Y=14430
X1334 87 M1M2_PR_DigitalLDOLogic_gds $T=48525 18670 0 0 $X=48365 $Y=18510
X1335 12 M1M2_PR_DigitalLDOLogic_gds $T=48870 10510 0 0 $X=48710 $Y=10350
X1336 84 M1M2_PR_DigitalLDOLogic_gds $T=48870 15950 0 0 $X=48710 $Y=15790
X1337 80 M1M2_PR_DigitalLDOLogic_gds $T=48870 16970 0 0 $X=48710 $Y=16810
X1338 80 M1M2_PR_DigitalLDOLogic_gds $T=48870 19350 0 0 $X=48710 $Y=19190
X1339 80 M1M2_PR_DigitalLDOLogic_gds $T=48870 24790 0 0 $X=48710 $Y=24630
X1340 80 M1M2_PR_DigitalLDOLogic_gds $T=48870 32950 0 0 $X=48710 $Y=32790
X1341 80 M1M2_PR_DigitalLDOLogic_gds $T=48870 35670 0 0 $X=48710 $Y=35510
X1342 91 M1M2_PR_DigitalLDOLogic_gds $T=51630 12210 0 0 $X=51470 $Y=12050
X1343 91 M1M2_PR_DigitalLDOLogic_gds $T=51630 13230 0 0 $X=51470 $Y=13070
X1344 79 M1M2_PR_DigitalLDOLogic_gds $T=51630 14250 0 0 $X=51470 $Y=14090
X1345 118 M1M2_PR_DigitalLDOLogic_gds $T=51630 14930 0 0 $X=51470 $Y=14770
X1346 118 M1M2_PR_DigitalLDOLogic_gds $T=51630 16970 0 0 $X=51470 $Y=16810
X1347 116 M1M2_PR_DigitalLDOLogic_gds $T=51630 17650 0 0 $X=51470 $Y=17490
X1348 116 M1M2_PR_DigitalLDOLogic_gds $T=51630 19010 0 0 $X=51470 $Y=18850
X1349 145 M1M2_PR_DigitalLDOLogic_gds $T=51630 21390 0 0 $X=51470 $Y=21230
X1350 117 M1M2_PR_DigitalLDOLogic_gds $T=51630 23090 0 0 $X=51470 $Y=22930
X1351 117 M1M2_PR_DigitalLDOLogic_gds $T=51630 24450 0 0 $X=51470 $Y=24290
X1352 145 M1M2_PR_DigitalLDOLogic_gds $T=51630 27510 0 0 $X=51470 $Y=27350
X1353 114 M1M2_PR_DigitalLDOLogic_gds $T=51630 28530 0 0 $X=51470 $Y=28370
X1354 115 M1M2_PR_DigitalLDOLogic_gds $T=51630 31250 0 0 $X=51470 $Y=31090
X1355 115 M1M2_PR_DigitalLDOLogic_gds $T=51630 33290 0 0 $X=51470 $Y=33130
X1356 114 M1M2_PR_DigitalLDOLogic_gds $T=51630 35330 0 0 $X=51470 $Y=35170
X1357 121 M1M2_PR_DigitalLDOLogic_gds $T=54390 14930 0 0 $X=54230 $Y=14770
X1358 121 M1M2_PR_DigitalLDOLogic_gds $T=54390 19010 0 0 $X=54230 $Y=18850
X1359 119 M1M2_PR_DigitalLDOLogic_gds $T=54390 20370 0 0 $X=54230 $Y=20210
X1360 119 M1M2_PR_DigitalLDOLogic_gds $T=54390 22750 0 0 $X=54230 $Y=22590
X1361 145 M1M2_PR_DigitalLDOLogic_gds $T=54390 27510 0 0 $X=54230 $Y=27350
X1362 145 M1M2_PR_DigitalLDOLogic_gds $T=54390 30230 0 0 $X=54230 $Y=30070
X1363 88 M1M2_PR_DigitalLDOLogic_gds $T=54390 30910 0 0 $X=54230 $Y=30750
X1364 88 M1M2_PR_DigitalLDOLogic_gds $T=54390 34990 0 0 $X=54230 $Y=34830
X1365 145 M1M2_PR_DigitalLDOLogic_gds $T=57150 13910 0 0 $X=56990 $Y=13750
X1366 145 M1M2_PR_DigitalLDOLogic_gds $T=57150 17310 0 0 $X=56990 $Y=17150
X1367 145 M1M2_PR_DigitalLDOLogic_gds $T=57150 18670 0 0 $X=56990 $Y=18510
X1368 145 M1M2_PR_DigitalLDOLogic_gds $T=57150 21390 0 0 $X=56990 $Y=21230
X1369 13 M1M2_PR_DigitalLDOLogic_gds $T=57150 24110 0 0 $X=56990 $Y=23950
X1370 89 M1M2_PR_DigitalLDOLogic_gds $T=57150 28190 0 0 $X=56990 $Y=28030
X1371 89 M1M2_PR_DigitalLDOLogic_gds $T=57150 32270 0 0 $X=56990 $Y=32110
X1372 78 M1M2_PR_DigitalLDOLogic_gds $T=59910 14250 0 0 $X=59750 $Y=14090
X1373 80 M1M2_PR_DigitalLDOLogic_gds $T=59910 16970 0 0 $X=59750 $Y=16810
X1374 80 M1M2_PR_DigitalLDOLogic_gds $T=59910 19350 0 0 $X=59750 $Y=19190
X1375 80 M1M2_PR_DigitalLDOLogic_gds $T=59910 23090 0 0 $X=59750 $Y=22930
X1376 80 M1M2_PR_DigitalLDOLogic_gds $T=59910 27850 0 0 $X=59750 $Y=27690
X1377 80 M1M2_PR_DigitalLDOLogic_gds $T=59910 30230 0 0 $X=59750 $Y=30070
X1378 92 M1M2_PR_DigitalLDOLogic_gds $T=62670 11530 0 0 $X=62510 $Y=11370
X1379 92 M1M2_PR_DigitalLDOLogic_gds $T=62670 13230 0 0 $X=62510 $Y=13070
X1380 10 M1M2_PR_DigitalLDOLogic_gds $T=62670 13910 0 0 $X=62510 $Y=13750
X1381 120 M1M2_PR_DigitalLDOLogic_gds $T=62670 14930 0 0 $X=62510 $Y=14770
X1382 120 M1M2_PR_DigitalLDOLogic_gds $T=62670 16970 0 0 $X=62510 $Y=16810
X1383 10 M1M2_PR_DigitalLDOLogic_gds $T=62670 18670 0 0 $X=62510 $Y=18510
X1384 92 M1M2_PR_DigitalLDOLogic_gds $T=62670 21390 0 0 $X=62510 $Y=21230
X1385 94 M1M2_PR_DigitalLDOLogic_gds $T=62670 25470 0 0 $X=62510 $Y=25310
X1386 94 M1M2_PR_DigitalLDOLogic_gds $T=62670 26830 0 0 $X=62510 $Y=26670
X1387 123 M1M2_PR_DigitalLDOLogic_gds $T=62670 28530 0 0 $X=62510 $Y=28370
X1388 123 M1M2_PR_DigitalLDOLogic_gds $T=62670 29890 0 0 $X=62510 $Y=29730
X1389 15 M1M2_PR_DigitalLDOLogic_gds $T=65430 11190 0 0 $X=65270 $Y=11030
X1390 91 M1M2_PR_DigitalLDOLogic_gds $T=65430 12210 0 0 $X=65270 $Y=12050
X1391 91 M1M2_PR_DigitalLDOLogic_gds $T=65430 15950 0 0 $X=65270 $Y=15790
X1392 91 M1M2_PR_DigitalLDOLogic_gds $T=65430 19690 0 0 $X=65270 $Y=19530
X1393 81 M1M2_PR_DigitalLDOLogic_gds $T=65430 22410 0 0 $X=65270 $Y=22250
X1394 145 M1M2_PR_DigitalLDOLogic_gds $T=65430 27510 0 0 $X=65270 $Y=27350
X1395 145 M1M2_PR_DigitalLDOLogic_gds $T=65430 32610 0 0 $X=65270 $Y=32450
X1396 16 M1M2_PR_DigitalLDOLogic_gds $T=68190 14250 0 0 $X=68030 $Y=14090
X1397 93 M1M2_PR_DigitalLDOLogic_gds $T=68190 14930 0 0 $X=68030 $Y=14770
X1398 93 M1M2_PR_DigitalLDOLogic_gds $T=68190 16630 0 0 $X=68030 $Y=16470
X1399 122 M1M2_PR_DigitalLDOLogic_gds $T=68190 17650 0 0 $X=68030 $Y=17490
X1400 93 M1M2_PR_DigitalLDOLogic_gds $T=68190 24110 0 0 $X=68030 $Y=23950
X1401 122 M1M2_PR_DigitalLDOLogic_gds $T=68190 27850 0 0 $X=68030 $Y=27690
X1402 79 M1M2_PR_DigitalLDOLogic_gds $T=70950 13910 0 0 $X=70790 $Y=13750
X1403 79 M1M2_PR_DigitalLDOLogic_gds $T=70950 16290 0 0 $X=70790 $Y=16130
X1404 90 M1M2_PR_DigitalLDOLogic_gds $T=70950 31250 0 0 $X=70790 $Y=31090
X1405 18 M1M2_PR_DigitalLDOLogic_gds $T=73710 11530 0 0 $X=73550 $Y=11370
X1406 92 M1M2_PR_DigitalLDOLogic_gds $T=73710 13230 0 0 $X=73550 $Y=13070
X1407 92 M1M2_PR_DigitalLDOLogic_gds $T=73710 15950 0 0 $X=73550 $Y=15790
X1408 78 M1M2_PR_DigitalLDOLogic_gds $T=73710 16630 0 0 $X=73550 $Y=16470
X1409 95 M1M2_PR_DigitalLDOLogic_gds $T=73710 17650 0 0 $X=73550 $Y=17490
X1410 95 M1M2_PR_DigitalLDOLogic_gds $T=73710 18670 0 0 $X=73550 $Y=18510
X1411 81 M1M2_PR_DigitalLDOLogic_gds $T=73710 19350 0 0 $X=73550 $Y=19190
X1412 81 M1M2_PR_DigitalLDOLogic_gds $T=73710 25130 0 0 $X=73550 $Y=24970
X1413 78 M1M2_PR_DigitalLDOLogic_gds $T=73710 27170 0 0 $X=73550 $Y=27010
X1414 79 M1M2_PR_DigitalLDOLogic_gds $T=73710 27850 0 0 $X=73550 $Y=27690
X1415 94 M1M2_PR_DigitalLDOLogic_gds $T=73710 28530 0 0 $X=73550 $Y=28370
X1416 94 M1M2_PR_DigitalLDOLogic_gds $T=73710 29550 0 0 $X=73550 $Y=29390
X1417 79 M1M2_PR_DigitalLDOLogic_gds $T=73710 30230 0 0 $X=73550 $Y=30070
X1418 78 M1M2_PR_DigitalLDOLogic_gds $T=73710 30910 0 0 $X=73550 $Y=30750
X1419 78 M1M2_PR_DigitalLDOLogic_gds $T=73710 32270 0 0 $X=73550 $Y=32110
X1420 17 M1M2_PR_DigitalLDOLogic_gds $T=76470 16630 0 0 $X=76310 $Y=16470
X1421 18 M1M2_PR_DigitalLDOLogic_gds $T=76470 23090 0 0 $X=76310 $Y=22930
X1422 18 M1M2_PR_DigitalLDOLogic_gds $T=76470 29550 0 0 $X=76310 $Y=29390
X1423 145 M1M2_PR_DigitalLDOLogic_gds $T=76470 30230 0 0 $X=76310 $Y=30070
X1424 145 M1M2_PR_DigitalLDOLogic_gds $T=76470 31250 0 0 $X=76310 $Y=31090
X1425 145 M1M2_PR_DigitalLDOLogic_gds $T=76470 32610 0 0 $X=76310 $Y=32450
X1426 19 M1M2_PR_DigitalLDOLogic_gds $T=79230 11190 0 0 $X=79070 $Y=11030
X1427 78 M1M2_PR_DigitalLDOLogic_gds $T=79230 16970 0 0 $X=79070 $Y=16810
X1428 125 M1M2_PR_DigitalLDOLogic_gds $T=79230 17650 0 0 $X=79070 $Y=17490
X1429 125 M1M2_PR_DigitalLDOLogic_gds $T=79230 19010 0 0 $X=79070 $Y=18850
X1430 78 M1M2_PR_DigitalLDOLogic_gds $T=79230 20370 0 0 $X=79070 $Y=20210
X1431 14 M1M2_PR_DigitalLDOLogic_gds $T=79230 22410 0 0 $X=79070 $Y=22250
X1432 126 M1M2_PR_DigitalLDOLogic_gds $T=79230 24450 0 0 $X=79070 $Y=24290
X1433 126 M1M2_PR_DigitalLDOLogic_gds $T=79230 29550 0 0 $X=79070 $Y=29390
X1434 79 M1M2_PR_DigitalLDOLogic_gds $T=79230 30230 0 0 $X=79070 $Y=30070
X1435 96 M1M2_PR_DigitalLDOLogic_gds $T=81990 11530 0 0 $X=81830 $Y=11370
X1436 96 M1M2_PR_DigitalLDOLogic_gds $T=81990 16290 0 0 $X=81830 $Y=16130
X1437 95 M1M2_PR_DigitalLDOLogic_gds $T=81990 17650 0 0 $X=81830 $Y=17490
X1438 95 M1M2_PR_DigitalLDOLogic_gds $T=81990 19010 0 0 $X=81830 $Y=18850
X1439 79 M1M2_PR_DigitalLDOLogic_gds $T=81990 19690 0 0 $X=81830 $Y=19530
X1440 81 M1M2_PR_DigitalLDOLogic_gds $T=81990 23090 0 0 $X=81830 $Y=22930
X1441 78 M1M2_PR_DigitalLDOLogic_gds $T=81990 30910 0 0 $X=81830 $Y=30750
X1442 78 M1M2_PR_DigitalLDOLogic_gds $T=81990 32270 0 0 $X=81830 $Y=32110
X1443 79 M1M2_PR_DigitalLDOLogic_gds $T=82375 13910 0 0 $X=82215 $Y=13750
X1444 78 M1M2_PR_DigitalLDOLogic_gds $T=84750 16290 0 0 $X=84590 $Y=16130
X1445 93 M1M2_PR_DigitalLDOLogic_gds $T=84750 18670 0 0 $X=84590 $Y=18510
X1446 124 M1M2_PR_DigitalLDOLogic_gds $T=84750 20370 0 0 $X=84590 $Y=20210
X1447 124 M1M2_PR_DigitalLDOLogic_gds $T=84750 21390 0 0 $X=84590 $Y=21230
X1448 93 M1M2_PR_DigitalLDOLogic_gds $T=84750 24110 0 0 $X=84590 $Y=23950
X1449 127 M1M2_PR_DigitalLDOLogic_gds $T=84750 27510 0 0 $X=84590 $Y=27350
X1450 127 M1M2_PR_DigitalLDOLogic_gds $T=84750 29550 0 0 $X=84590 $Y=29390
X1451 78 M1M2_PR_DigitalLDOLogic_gds $T=84750 30570 0 0 $X=84590 $Y=30410
X1452 78 M1M2_PR_DigitalLDOLogic_gds $T=84750 32270 0 0 $X=84590 $Y=32110
X1453 20 M1M2_PR_DigitalLDOLogic_gds $T=86130 650 0 0 $X=85970 $Y=490
X1454 21 M1M2_PR_DigitalLDOLogic_gds $T=87510 10510 0 0 $X=87350 $Y=10350
X1455 96 M1M2_PR_DigitalLDOLogic_gds $T=87510 11870 0 0 $X=87350 $Y=11710
X1456 79 M1M2_PR_DigitalLDOLogic_gds $T=87510 14930 0 0 $X=87350 $Y=14770
X1457 79 M1M2_PR_DigitalLDOLogic_gds $T=87510 15950 0 0 $X=87350 $Y=15790
X1458 79 M1M2_PR_DigitalLDOLogic_gds $T=87510 16970 0 0 $X=87350 $Y=16810
X1459 96 M1M2_PR_DigitalLDOLogic_gds $T=87510 18670 0 0 $X=87350 $Y=18510
X1460 145 M1M2_PR_DigitalLDOLogic_gds $T=87510 19690 0 0 $X=87350 $Y=19530
X1461 145 M1M2_PR_DigitalLDOLogic_gds $T=87510 31250 0 0 $X=87350 $Y=31090
X1462 97 M1M2_PR_DigitalLDOLogic_gds $T=90270 11530 0 0 $X=90110 $Y=11370
X1463 97 M1M2_PR_DigitalLDOLogic_gds $T=90270 14590 0 0 $X=90110 $Y=14430
X1464 97 M1M2_PR_DigitalLDOLogic_gds $T=90270 19010 0 0 $X=90110 $Y=18850
X1465 97 M1M2_PR_DigitalLDOLogic_gds $T=90270 21390 0 0 $X=90110 $Y=21230
X1466 81 M1M2_PR_DigitalLDOLogic_gds $T=90270 22410 0 0 $X=90110 $Y=22250
X1467 81 M1M2_PR_DigitalLDOLogic_gds $T=90270 24790 0 0 $X=90110 $Y=24630
X1468 98 M1M2_PR_DigitalLDOLogic_gds $T=90270 28530 0 0 $X=90110 $Y=28370
X1469 98 M1M2_PR_DigitalLDOLogic_gds $T=90270 29890 0 0 $X=90110 $Y=29730
X1470 20 M1M2_PR_DigitalLDOLogic_gds $T=93030 650 0 0 $X=92870 $Y=490
X1471 20 M1M2_PR_DigitalLDOLogic_gds $T=93030 11190 0 0 $X=92870 $Y=11030
X1472 78 M1M2_PR_DigitalLDOLogic_gds $T=93030 13230 0 0 $X=92870 $Y=13070
X1473 78 M1M2_PR_DigitalLDOLogic_gds $T=93030 16630 0 0 $X=92870 $Y=16470
X1474 129 M1M2_PR_DigitalLDOLogic_gds $T=93030 17650 0 0 $X=92870 $Y=17490
X1475 129 M1M2_PR_DigitalLDOLogic_gds $T=93030 19010 0 0 $X=92870 $Y=18850
X1476 81 M1M2_PR_DigitalLDOLogic_gds $T=93030 19690 0 0 $X=92870 $Y=19530
X1477 81 M1M2_PR_DigitalLDOLogic_gds $T=93030 22410 0 0 $X=92870 $Y=22250
X1478 127 M1M2_PR_DigitalLDOLogic_gds $T=93030 23090 0 0 $X=92870 $Y=22930
X1479 127 M1M2_PR_DigitalLDOLogic_gds $T=93030 27170 0 0 $X=92870 $Y=27010
X1480 79 M1M2_PR_DigitalLDOLogic_gds $T=93030 27850 0 0 $X=92870 $Y=27690
X1481 79 M1M2_PR_DigitalLDOLogic_gds $T=93030 29890 0 0 $X=92870 $Y=29730
X1482 22 M1M2_PR_DigitalLDOLogic_gds $T=95790 11190 0 0 $X=95630 $Y=11030
X1483 128 M1M2_PR_DigitalLDOLogic_gds $T=95790 13230 0 0 $X=95630 $Y=13070
X1484 145 M1M2_PR_DigitalLDOLogic_gds $T=95790 13910 0 0 $X=95630 $Y=13750
X1485 145 M1M2_PR_DigitalLDOLogic_gds $T=95790 16970 0 0 $X=95630 $Y=16810
X1486 145 M1M2_PR_DigitalLDOLogic_gds $T=95790 19010 0 0 $X=95630 $Y=18850
X1487 96 M1M2_PR_DigitalLDOLogic_gds $T=95790 20370 0 0 $X=95630 $Y=20210
X1488 128 M1M2_PR_DigitalLDOLogic_gds $T=95790 24110 0 0 $X=95630 $Y=23950
X1489 96 M1M2_PR_DigitalLDOLogic_gds $T=95790 29550 0 0 $X=95630 $Y=29390
X1490 101 M1M2_PR_DigitalLDOLogic_gds $T=95790 30230 0 0 $X=95630 $Y=30070
X1491 98 M1M2_PR_DigitalLDOLogic_gds $T=98550 11530 0 0 $X=98390 $Y=11370
X1492 98 M1M2_PR_DigitalLDOLogic_gds $T=98550 13230 0 0 $X=98390 $Y=13070
X1493 98 M1M2_PR_DigitalLDOLogic_gds $T=98550 24110 0 0 $X=98390 $Y=23950
X1494 98 M1M2_PR_DigitalLDOLogic_gds $T=98550 28190 0 0 $X=98390 $Y=28030
X1495 23 M1M2_PR_DigitalLDOLogic_gds $T=101310 16290 0 0 $X=101150 $Y=16130
X1496 100 M1M2_PR_DigitalLDOLogic_gds $T=101310 16970 0 0 $X=101150 $Y=16810
X1497 100 M1M2_PR_DigitalLDOLogic_gds $T=101310 21390 0 0 $X=101150 $Y=21230
X1498 130 M1M2_PR_DigitalLDOLogic_gds $T=101310 22750 0 0 $X=101150 $Y=22590
X1499 130 M1M2_PR_DigitalLDOLogic_gds $T=101310 29550 0 0 $X=101150 $Y=29390
X1500 24 M1M2_PR_DigitalLDOLogic_gds $T=104070 14250 0 0 $X=103910 $Y=14090
X1501 79 M1M2_PR_DigitalLDOLogic_gds $T=104070 15950 0 0 $X=103910 $Y=15790
X1502 79 M1M2_PR_DigitalLDOLogic_gds $T=104070 17650 0 0 $X=103910 $Y=17490
X1503 25 M1M2_PR_DigitalLDOLogic_gds $T=106830 19010 0 0 $X=106670 $Y=18850
X1504 78 M1M2_PR_DigitalLDOLogic_gds $T=109590 15950 0 0 $X=109430 $Y=15790
X1505 79 M1M2_PR_DigitalLDOLogic_gds $T=109590 17650 0 0 $X=109430 $Y=17490
X1506 79 M1M2_PR_DigitalLDOLogic_gds $T=109590 24790 0 0 $X=109430 $Y=24630
X1507 79 M1M2_PR_DigitalLDOLogic_gds $T=109590 27850 0 0 $X=109430 $Y=27690
X1508 101 M1M2_PR_DigitalLDOLogic_gds $T=109590 29550 0 0 $X=109430 $Y=29390
X1509 99 M1M2_PR_DigitalLDOLogic_gds $T=112350 13910 0 0 $X=112190 $Y=13750
X1510 78 M1M2_PR_DigitalLDOLogic_gds $T=112350 15950 0 0 $X=112190 $Y=15790
X1511 78 M1M2_PR_DigitalLDOLogic_gds $T=112350 16970 0 0 $X=112190 $Y=16810
X1512 131 M1M2_PR_DigitalLDOLogic_gds $T=112350 17650 0 0 $X=112190 $Y=17490
X1513 131 M1M2_PR_DigitalLDOLogic_gds $T=112350 22750 0 0 $X=112190 $Y=22590
X1514 78 M1M2_PR_DigitalLDOLogic_gds $T=112350 24110 0 0 $X=112190 $Y=23950
X1515 145 M1M2_PR_DigitalLDOLogic_gds $T=112350 25810 0 0 $X=112190 $Y=25650
X1516 79 M1M2_PR_DigitalLDOLogic_gds $T=112350 27850 0 0 $X=112190 $Y=27690
X1517 79 M1M2_PR_DigitalLDOLogic_gds $T=112350 30230 0 0 $X=112190 $Y=30070
X1518 145 M1M2_PR_DigitalLDOLogic_gds $T=112350 30910 0 0 $X=112190 $Y=30750
X1519 145 M1M2_PR_DigitalLDOLogic_gds $T=112350 32270 0 0 $X=112190 $Y=32110
X1520 26 M1M2_PR_DigitalLDOLogic_gds $T=115110 14250 0 0 $X=114950 $Y=14090
X1521 99 M1M2_PR_DigitalLDOLogic_gds $T=115110 18670 0 0 $X=114950 $Y=18510
X1522 101 M1M2_PR_DigitalLDOLogic_gds $T=115110 19350 0 0 $X=114950 $Y=19190
X1523 101 M1M2_PR_DigitalLDOLogic_gds $T=115110 21390 0 0 $X=114950 $Y=21230
X1524 101 M1M2_PR_DigitalLDOLogic_gds $T=115110 29550 0 0 $X=114950 $Y=29390
X1525 102 M1M2_PR_DigitalLDOLogic_gds $T=117870 12210 0 0 $X=117710 $Y=12050
X1526 102 M1M2_PR_DigitalLDOLogic_gds $T=117870 13910 0 0 $X=117710 $Y=13750
X1527 145 M1M2_PR_DigitalLDOLogic_gds $T=117870 16970 0 0 $X=117710 $Y=16810
X1528 145 M1M2_PR_DigitalLDOLogic_gds $T=117870 19010 0 0 $X=117710 $Y=18850
X1529 82 M1M2_PR_DigitalLDOLogic_gds $T=117870 19690 0 0 $X=117710 $Y=19530
X1530 82 M1M2_PR_DigitalLDOLogic_gds $T=117870 22410 0 0 $X=117710 $Y=22250
X1531 82 M1M2_PR_DigitalLDOLogic_gds $T=117870 24790 0 0 $X=117710 $Y=24630
X1532 85 M1M2_PR_DigitalLDOLogic_gds $T=117870 25810 0 0 $X=117710 $Y=25650
X1533 85 M1M2_PR_DigitalLDOLogic_gds $T=117870 28190 0 0 $X=117710 $Y=28030
X1534 85 M1M2_PR_DigitalLDOLogic_gds $T=117870 38390 0 0 $X=117710 $Y=38230
X1535 79 M1M2_PR_DigitalLDOLogic_gds $T=118270 14590 0 0 $X=118110 $Y=14430
X1536 79 M1M2_PR_DigitalLDOLogic_gds $T=118270 16290 0 0 $X=118110 $Y=16130
X1537 132 M1M2_PR_DigitalLDOLogic_gds $T=120630 13230 0 0 $X=120470 $Y=13070
X1538 28 M1M2_PR_DigitalLDOLogic_gds $T=120630 16630 0 0 $X=120470 $Y=16470
X1539 132 M1M2_PR_DigitalLDOLogic_gds $T=120630 19010 0 0 $X=120470 $Y=18850
X1540 78 M1M2_PR_DigitalLDOLogic_gds $T=120630 27170 0 0 $X=120470 $Y=27010
X1541 78 M1M2_PR_DigitalLDOLogic_gds $T=120630 27850 0 0 $X=120470 $Y=27690
X1542 78 M1M2_PR_DigitalLDOLogic_gds $T=120630 30230 0 0 $X=120470 $Y=30070
X1543 27 M1M2_PR_DigitalLDOLogic_gds $T=123390 11190 0 0 $X=123230 $Y=11030
X1544 102 M1M2_PR_DigitalLDOLogic_gds $T=123390 12210 0 0 $X=123230 $Y=12050
X1545 102 M1M2_PR_DigitalLDOLogic_gds $T=123390 13570 0 0 $X=123230 $Y=13410
X1546 79 M1M2_PR_DigitalLDOLogic_gds $T=123390 14930 0 0 $X=123230 $Y=14770
X1547 79 M1M2_PR_DigitalLDOLogic_gds $T=123390 16290 0 0 $X=123230 $Y=16130
X1548 99 M1M2_PR_DigitalLDOLogic_gds $T=123390 17310 0 0 $X=123230 $Y=17150
X1549 99 M1M2_PR_DigitalLDOLogic_gds $T=123390 18670 0 0 $X=123230 $Y=18510
X1550 145 M1M2_PR_DigitalLDOLogic_gds $T=123390 19350 0 0 $X=123230 $Y=19190
X1551 82 M1M2_PR_DigitalLDOLogic_gds $T=123390 22410 0 0 $X=123230 $Y=22250
X1552 82 M1M2_PR_DigitalLDOLogic_gds $T=123390 27510 0 0 $X=123230 $Y=27350
X1553 145 M1M2_PR_DigitalLDOLogic_gds $T=123390 28190 0 0 $X=123230 $Y=28030
X1554 145 M1M2_PR_DigitalLDOLogic_gds $T=123390 30230 0 0 $X=123230 $Y=30070
X1555 145 M1M2_PR_DigitalLDOLogic_gds $T=123390 32270 0 0 $X=123230 $Y=32110
X1556 103 M1M2_PR_DigitalLDOLogic_gds $T=126150 11530 0 0 $X=125990 $Y=11370
X1557 103 M1M2_PR_DigitalLDOLogic_gds $T=126150 16290 0 0 $X=125990 $Y=16130
X1558 78 M1M2_PR_DigitalLDOLogic_gds $T=126150 16970 0 0 $X=125990 $Y=16810
X1559 104 M1M2_PR_DigitalLDOLogic_gds $T=126150 17650 0 0 $X=125990 $Y=17490
X1560 104 M1M2_PR_DigitalLDOLogic_gds $T=126150 21390 0 0 $X=125990 $Y=21230
X1561 134 M1M2_PR_DigitalLDOLogic_gds $T=126150 22750 0 0 $X=125990 $Y=22590
X1562 113 M1M2_PR_DigitalLDOLogic_gds $T=126150 24790 0 0 $X=125990 $Y=24630
X1563 113 M1M2_PR_DigitalLDOLogic_gds $T=126150 26830 0 0 $X=125990 $Y=26670
X1564 134 M1M2_PR_DigitalLDOLogic_gds $T=126150 29550 0 0 $X=125990 $Y=29390
X1565 78 M1M2_PR_DigitalLDOLogic_gds $T=126150 30570 0 0 $X=125990 $Y=30410
X1566 145 M1M2_PR_DigitalLDOLogic_gds $T=128910 13910 0 0 $X=128750 $Y=13750
X1567 79 M1M2_PR_DigitalLDOLogic_gds $T=128910 14590 0 0 $X=128750 $Y=14430
X1568 145 M1M2_PR_DigitalLDOLogic_gds $T=128910 16970 0 0 $X=128750 $Y=16810
X1569 79 M1M2_PR_DigitalLDOLogic_gds $T=128910 18670 0 0 $X=128750 $Y=18510
X1570 145 M1M2_PR_DigitalLDOLogic_gds $T=128910 19350 0 0 $X=128750 $Y=19190
X1571 82 M1M2_PR_DigitalLDOLogic_gds $T=128910 20030 0 0 $X=128750 $Y=19870
X1572 82 M1M2_PR_DigitalLDOLogic_gds $T=128910 22410 0 0 $X=128750 $Y=22250
X1573 145 M1M2_PR_DigitalLDOLogic_gds $T=128910 24110 0 0 $X=128750 $Y=23950
X1574 78 M1M2_PR_DigitalLDOLogic_gds $T=131670 14250 0 0 $X=131510 $Y=14090
X1575 78 M1M2_PR_DigitalLDOLogic_gds $T=131670 16970 0 0 $X=131510 $Y=16810
X1576 136 M1M2_PR_DigitalLDOLogic_gds $T=131670 17650 0 0 $X=131510 $Y=17490
X1577 136 M1M2_PR_DigitalLDOLogic_gds $T=131670 19010 0 0 $X=131510 $Y=18850
X1578 104 M1M2_PR_DigitalLDOLogic_gds $T=131670 21390 0 0 $X=131510 $Y=21230
X1579 14 M1M2_PR_DigitalLDOLogic_gds $T=131670 22410 0 0 $X=131510 $Y=22250
X1580 104 M1M2_PR_DigitalLDOLogic_gds $T=131670 25130 0 0 $X=131510 $Y=24970
X1581 112 M1M2_PR_DigitalLDOLogic_gds $T=131670 27850 0 0 $X=131510 $Y=27690
X1582 30 M1M2_PR_DigitalLDOLogic_gds $T=134430 14250 0 0 $X=134270 $Y=14090
X1583 105 M1M2_PR_DigitalLDOLogic_gds $T=134430 14930 0 0 $X=134270 $Y=14770
X1584 105 M1M2_PR_DigitalLDOLogic_gds $T=134430 16630 0 0 $X=134270 $Y=16470
X1585 105 M1M2_PR_DigitalLDOLogic_gds $T=134430 20370 0 0 $X=134270 $Y=20210
X1586 82 M1M2_PR_DigitalLDOLogic_gds $T=134430 23090 0 0 $X=134270 $Y=22930
X1587 82 M1M2_PR_DigitalLDOLogic_gds $T=134430 27510 0 0 $X=134270 $Y=27350
X1588 31 M1M2_PR_DigitalLDOLogic_gds $T=137190 11190 0 0 $X=137030 $Y=11030
X1589 102 M1M2_PR_DigitalLDOLogic_gds $T=137190 13570 0 0 $X=137030 $Y=13410
X1590 102 M1M2_PR_DigitalLDOLogic_gds $T=137190 17650 0 0 $X=137030 $Y=17490
X1591 102 M1M2_PR_DigitalLDOLogic_gds $T=137190 18670 0 0 $X=137030 $Y=18510
X1592 137 M1M2_PR_DigitalLDOLogic_gds $T=137190 22750 0 0 $X=137030 $Y=22590
X1593 137 M1M2_PR_DigitalLDOLogic_gds $T=137190 24110 0 0 $X=137030 $Y=23950
X1594 145 M1M2_PR_DigitalLDOLogic_gds $T=137190 24790 0 0 $X=137030 $Y=24630
X1595 138 M1M2_PR_DigitalLDOLogic_gds $T=137190 28190 0 0 $X=137030 $Y=28030
X1596 138 M1M2_PR_DigitalLDOLogic_gds $T=137190 29550 0 0 $X=137030 $Y=29390
X1597 145 M1M2_PR_DigitalLDOLogic_gds $T=137190 30230 0 0 $X=137030 $Y=30070
X1598 106 M1M2_PR_DigitalLDOLogic_gds $T=139950 11530 0 0 $X=139790 $Y=11370
X1599 140 M1M2_PR_DigitalLDOLogic_gds $T=139950 17650 0 0 $X=139790 $Y=17490
X1600 106 M1M2_PR_DigitalLDOLogic_gds $T=139950 23090 0 0 $X=139790 $Y=22930
X1601 106 M1M2_PR_DigitalLDOLogic_gds $T=139950 29890 0 0 $X=139790 $Y=29730
X1602 32 M1M2_PR_DigitalLDOLogic_gds $T=142710 14250 0 0 $X=142550 $Y=14090
X1603 78 M1M2_PR_DigitalLDOLogic_gds $T=142710 16290 0 0 $X=142550 $Y=16130
X1604 79 M1M2_PR_DigitalLDOLogic_gds $T=142710 16970 0 0 $X=142550 $Y=16810
X1605 145 M1M2_PR_DigitalLDOLogic_gds $T=142710 17650 0 0 $X=142550 $Y=17490
X1606 145 M1M2_PR_DigitalLDOLogic_gds $T=142710 18670 0 0 $X=142550 $Y=18510
X1607 79 M1M2_PR_DigitalLDOLogic_gds $T=142710 19350 0 0 $X=142550 $Y=19190
X1608 78 M1M2_PR_DigitalLDOLogic_gds $T=142710 20030 0 0 $X=142550 $Y=19870
X1609 79 M1M2_PR_DigitalLDOLogic_gds $T=142710 24790 0 0 $X=142550 $Y=24630
X1610 78 M1M2_PR_DigitalLDOLogic_gds $T=142710 25470 0 0 $X=142550 $Y=25310
X1611 78 M1M2_PR_DigitalLDOLogic_gds $T=142710 27170 0 0 $X=142550 $Y=27010
X1612 78 M1M2_PR_DigitalLDOLogic_gds $T=142710 29550 0 0 $X=142550 $Y=29390
X1613 78 M1M2_PR_DigitalLDOLogic_gds $T=142710 31250 0 0 $X=142550 $Y=31090
X1614 107 M1M2_PR_DigitalLDOLogic_gds $T=145470 13910 0 0 $X=145310 $Y=13750
X1615 107 M1M2_PR_DigitalLDOLogic_gds $T=145470 16290 0 0 $X=145310 $Y=16130
X1616 143 M1M2_PR_DigitalLDOLogic_gds $T=145470 17650 0 0 $X=145310 $Y=17490
X1617 143 M1M2_PR_DigitalLDOLogic_gds $T=145470 18670 0 0 $X=145310 $Y=18510
X1618 108 M1M2_PR_DigitalLDOLogic_gds $T=145470 24450 0 0 $X=145310 $Y=24290
X1619 108 M1M2_PR_DigitalLDOLogic_gds $T=145470 26830 0 0 $X=145310 $Y=26670
X1620 109 M1M2_PR_DigitalLDOLogic_gds $T=148230 11530 0 0 $X=148070 $Y=11370
X1621 139 M1M2_PR_DigitalLDOLogic_gds $T=148230 17650 0 0 $X=148070 $Y=17490
X1622 139 M1M2_PR_DigitalLDOLogic_gds $T=148230 19010 0 0 $X=148070 $Y=18850
X1623 109 M1M2_PR_DigitalLDOLogic_gds $T=148230 19690 0 0 $X=148070 $Y=19530
X1624 145 M1M2_PR_DigitalLDOLogic_gds $T=148230 22410 0 0 $X=148070 $Y=22250
X1625 145 M1M2_PR_DigitalLDOLogic_gds $T=148230 24110 0 0 $X=148070 $Y=23950
X1626 140 M1M2_PR_DigitalLDOLogic_gds $T=150990 16630 0 0 $X=150830 $Y=16470
X1627 33 M1M2_PR_DigitalLDOLogic_gds $T=150990 25130 0 0 $X=150830 $Y=24970
X1628 79 M1M2_PR_DigitalLDOLogic_gds $T=150990 25810 0 0 $X=150830 $Y=25650
X1629 79 M1M2_PR_DigitalLDOLogic_gds $T=150990 27850 0 0 $X=150830 $Y=27690
X1630 79 M1M2_PR_DigitalLDOLogic_gds $T=150990 29890 0 0 $X=150830 $Y=29730
X1631 34 M1M2_PR_DigitalLDOLogic_gds $T=153750 11190 0 0 $X=153590 $Y=11030
X1632 83 M1M2_PR_DigitalLDOLogic_gds $T=153750 16970 0 0 $X=153590 $Y=16810
X1633 83 M1M2_PR_DigitalLDOLogic_gds $T=153750 19350 0 0 $X=153590 $Y=19190
X1634 83 M1M2_PR_DigitalLDOLogic_gds $T=153750 22070 0 0 $X=153590 $Y=21910
X1635 141 M1M2_PR_DigitalLDOLogic_gds $T=153750 22750 0 0 $X=153590 $Y=22590
X1636 141 M1M2_PR_DigitalLDOLogic_gds $T=153750 24110 0 0 $X=153590 $Y=23950
X1637 78 M1M2_PR_DigitalLDOLogic_gds $T=153750 25470 0 0 $X=153590 $Y=25310
X1638 78 M1M2_PR_DigitalLDOLogic_gds $T=153750 26830 0 0 $X=153590 $Y=26670
X1639 110 M1M2_PR_DigitalLDOLogic_gds $T=156510 16970 0 0 $X=156350 $Y=16810
X1640 110 M1M2_PR_DigitalLDOLogic_gds $T=156510 23090 0 0 $X=156350 $Y=22930
X1641 110 M1M2_PR_DigitalLDOLogic_gds $T=156510 28190 0 0 $X=156350 $Y=28030
X1642 110 M1M2_PR_DigitalLDOLogic_gds $T=156510 30230 0 0 $X=156350 $Y=30070
X1643 145 M1M2_PR_DigitalLDOLogic_gds $T=159270 13910 0 0 $X=159110 $Y=13750
X1644 145 M1M2_PR_DigitalLDOLogic_gds $T=159270 22410 0 0 $X=159110 $Y=22250
X1645 145 M1M2_PR_DigitalLDOLogic_gds $T=159270 27850 0 0 $X=159110 $Y=27690
X1646 35 M1M2_PR_DigitalLDOLogic_gds $T=162030 11190 0 0 $X=161870 $Y=11030
X1647 83 M1M2_PR_DigitalLDOLogic_gds $T=162030 22410 0 0 $X=161870 $Y=22250
X1648 142 M1M2_PR_DigitalLDOLogic_gds $T=162030 23090 0 0 $X=161870 $Y=22930
X1649 142 M1M2_PR_DigitalLDOLogic_gds $T=162030 26830 0 0 $X=161870 $Y=26670
X1650 36 M1M2_PR_DigitalLDOLogic_gds $T=164790 16630 0 0 $X=164630 $Y=16470
X1651 83 M1M2_PR_DigitalLDOLogic_gds $T=164790 19350 0 0 $X=164630 $Y=19190
X1652 112 M1M2_PR_DigitalLDOLogic_gds $T=164790 23090 0 0 $X=164630 $Y=22930
X1653 112 M1M2_PR_DigitalLDOLogic_gds $T=164790 24110 0 0 $X=164630 $Y=23950
X1654 111 M1M2_PR_DigitalLDOLogic_gds $T=167550 12210 0 0 $X=167390 $Y=12050
X1655 111 M1M2_PR_DigitalLDOLogic_gds $T=167550 13570 0 0 $X=167390 $Y=13410
X1656 77 M1M2_PR_DigitalLDOLogic_gds $T=167550 14930 0 0 $X=167390 $Y=14770
X1657 77 M1M2_PR_DigitalLDOLogic_gds $T=167550 18670 0 0 $X=167390 $Y=18510
X1658 79 M1M2_PR_DigitalLDOLogic_gds $T=167550 20370 0 0 $X=167390 $Y=20210
X1659 79 M1M2_PR_DigitalLDOLogic_gds $T=167550 24450 0 0 $X=167390 $Y=24290
X1660 78 M1M2_PR_DigitalLDOLogic_gds $T=167550 25470 0 0 $X=167390 $Y=25310
X1661 78 M1M2_PR_DigitalLDOLogic_gds $T=167550 26830 0 0 $X=167390 $Y=26670
X1662 29 M1M2_PR_DigitalLDOLogic_gds $T=170310 13910 0 0 $X=170150 $Y=13750
X1663 83 M1M2_PR_DigitalLDOLogic_gds $T=170310 17310 0 0 $X=170150 $Y=17150
X1664 83 M1M2_PR_DigitalLDOLogic_gds $T=170310 21730 0 0 $X=170150 $Y=21570
X1665 14 M1M2_PR_DigitalLDOLogic_gds $T=170310 22410 0 0 $X=170150 $Y=22250
X1666 29 M1M2_PR_DigitalLDOLogic_gds $T=170310 23090 0 0 $X=170150 $Y=22930
X1667 29 M1M2_PR_DigitalLDOLogic_gds $T=170310 32950 0 0 $X=170150 $Y=32790
X1668 109 M1M2_PR_DigitalLDOLogic_gds $T=173070 10510 0 0 $X=172910 $Y=10350
X1669 37 M1M2_PR_DigitalLDOLogic_gds $T=173070 13910 0 0 $X=172910 $Y=13750
X1670 37 M1M2_PR_DigitalLDOLogic_gds $T=173070 19350 0 0 $X=172910 $Y=19190
X1671 109 M1M2_PR_DigitalLDOLogic_gds $T=173070 20030 0 0 $X=172910 $Y=19870
X1672 78 M1M2_PR_DigitalLDOLogic_gds $T=173070 22750 0 0 $X=172910 $Y=22590
X1673 109 M1M2_PR_DigitalLDOLogic_gds $T=173070 24110 0 0 $X=172910 $Y=23950
X1674 78 M1M2_PR_DigitalLDOLogic_gds $T=173070 24790 0 0 $X=172910 $Y=24630
X1675 37 M1M2_PR_DigitalLDOLogic_gds $T=173530 9490 0 0 $X=173370 $Y=9330
X1676 107 M1M2_PR_DigitalLDOLogic_gds $T=175830 14590 0 0 $X=175670 $Y=14430
X1677 107 M1M2_PR_DigitalLDOLogic_gds $T=175830 15950 0 0 $X=175670 $Y=15790
X1678 112 M1M2_PR_DigitalLDOLogic_gds $T=175830 16970 0 0 $X=175670 $Y=16810
X1679 112 M1M2_PR_DigitalLDOLogic_gds $T=175830 21390 0 0 $X=175670 $Y=21230
X1680 144 M1M2_PR_DigitalLDOLogic_gds $T=175830 22750 0 0 $X=175670 $Y=22590
X1681 144 M1M2_PR_DigitalLDOLogic_gds $T=175830 24110 0 0 $X=175670 $Y=23950
X1682 38 M1M2_PR_DigitalLDOLogic_gds $T=178590 16630 0 0 $X=178430 $Y=16470
X1683 37 M1M2_PR_DigitalLDOLogic_gds $T=180430 9490 0 0 $X=180270 $Y=9330
X1684 113 M1M2_PR_DigitalLDOLogic_gds $T=181350 24790 0 0 $X=181190 $Y=24630
X1685 113 M1M2_PR_DigitalLDOLogic_gds $T=181350 28190 0 0 $X=181190 $Y=28030
X1686 111 M1M2_PR_DigitalLDOLogic_gds $T=184110 13570 0 0 $X=183950 $Y=13410
X1687 111 M1M2_PR_DigitalLDOLogic_gds $T=184110 21390 0 0 $X=183950 $Y=21230
X1688 39 M1M2_PR_DigitalLDOLogic_gds $T=186870 24450 0 0 $X=186710 $Y=24290
X1689 3 M2M3_PR_DigitalLDOLogic_gds $T=15750 1630 0 0 $X=15585 $Y=1445
X1690 6 M2M3_PR_DigitalLDOLogic_gds $T=26790 1020 0 0 $X=26625 $Y=835
X1691 8 M2M3_PR_DigitalLDOLogic_gds $T=35070 1020 0 0 $X=34905 $Y=835
X1692 79 M2M3_PR_DigitalLDOLogic_gds $T=43350 15050 0 0 $X=43185 $Y=14865
X1693 10 M2M3_PR_DigitalLDOLogic_gds $T=46570 8950 0 0 $X=46405 $Y=8765
X1694 12 M2M3_PR_DigitalLDOLogic_gds $T=48870 10170 0 0 $X=48705 $Y=9985
X1695 80 M2M3_PR_DigitalLDOLogic_gds $T=48870 22980 0 0 $X=48705 $Y=22795
X1696 79 M2M3_PR_DigitalLDOLogic_gds $T=51630 14440 0 0 $X=51465 $Y=14255
X1697 145 M2M3_PR_DigitalLDOLogic_gds $T=54390 27250 0 0 $X=54225 $Y=27065
X1698 78 M2M3_PR_DigitalLDOLogic_gds $T=59910 15050 0 0 $X=59745 $Y=14865
X1699 80 M2M3_PR_DigitalLDOLogic_gds $T=59910 22980 0 0 $X=59745 $Y=22795
X1700 10 M2M3_PR_DigitalLDOLogic_gds $T=62670 13830 0 0 $X=62505 $Y=13645
X1701 15 M2M3_PR_DigitalLDOLogic_gds $T=65430 1020 0 0 $X=65265 $Y=835
X1702 81 M2M3_PR_DigitalLDOLogic_gds $T=65430 26030 0 0 $X=65265 $Y=25845
X1703 145 M2M3_PR_DigitalLDOLogic_gds $T=65430 27250 0 0 $X=65265 $Y=27065
X1704 18 M2M3_PR_DigitalLDOLogic_gds $T=73710 10780 0 0 $X=73545 $Y=10595
X1705 81 M2M3_PR_DigitalLDOLogic_gds $T=73710 26030 0 0 $X=73545 $Y=25845
X1706 79 M2M3_PR_DigitalLDOLogic_gds $T=73710 30300 0 0 $X=73545 $Y=30115
X1707 17 M2M3_PR_DigitalLDOLogic_gds $T=76470 3460 0 0 $X=76305 $Y=3275
X1708 18 M2M3_PR_DigitalLDOLogic_gds $T=76470 18100 0 0 $X=76305 $Y=17915
X1709 78 M2M3_PR_DigitalLDOLogic_gds $T=79230 15050 0 0 $X=79065 $Y=14865
X1710 14 M2M3_PR_DigitalLDOLogic_gds $T=79230 22370 0 0 $X=79065 $Y=22185
X1711 79 M2M3_PR_DigitalLDOLogic_gds $T=79230 30300 0 0 $X=79065 $Y=30115
X1712 81 M2M3_PR_DigitalLDOLogic_gds $T=81990 26030 0 0 $X=81825 $Y=25845
X1713 78 M2M3_PR_DigitalLDOLogic_gds $T=84750 15050 0 0 $X=84585 $Y=14865
X1714 21 M2M3_PR_DigitalLDOLogic_gds $T=87510 10170 0 0 $X=87345 $Y=9985
X1715 78 M2M3_PR_DigitalLDOLogic_gds $T=93030 15050 0 0 $X=92865 $Y=14865
X1716 79 M2M3_PR_DigitalLDOLogic_gds $T=93030 30910 0 0 $X=92865 $Y=30725
X1717 101 M2M3_PR_DigitalLDOLogic_gds $T=95790 30300 0 0 $X=95625 $Y=30115
X1718 23 M2M3_PR_DigitalLDOLogic_gds $T=101310 2850 0 0 $X=101145 $Y=2665
X1719 25 M2M3_PR_DigitalLDOLogic_gds $T=107290 8950 0 0 $X=107125 $Y=8765
X1720 78 M2M3_PR_DigitalLDOLogic_gds $T=109590 15050 0 0 $X=109425 $Y=14865
X1721 101 M2M3_PR_DigitalLDOLogic_gds $T=109590 30300 0 0 $X=109425 $Y=30115
X1722 99 M2M3_PR_DigitalLDOLogic_gds $T=112350 15050 0 0 $X=112185 $Y=14865
X1723 99 M2M3_PR_DigitalLDOLogic_gds $T=115110 15050 0 0 $X=114945 $Y=14865
X1724 28 M2M3_PR_DigitalLDOLogic_gds $T=120630 14440 0 0 $X=120465 $Y=14255
X1725 145 M2M3_PR_DigitalLDOLogic_gds $T=128910 18100 0 0 $X=128745 $Y=17915
X1726 78 M2M3_PR_DigitalLDOLogic_gds $T=131670 15050 0 0 $X=131505 $Y=14865
X1727 14 M2M3_PR_DigitalLDOLogic_gds $T=131670 22370 0 0 $X=131505 $Y=22185
X1728 112 M2M3_PR_DigitalLDOLogic_gds $T=131670 26030 0 0 $X=131505 $Y=25845
X1729 31 M2M3_PR_DigitalLDOLogic_gds $T=137190 1020 0 0 $X=137025 $Y=835
X1730 140 M2M3_PR_DigitalLDOLogic_gds $T=140410 9560 0 0 $X=140245 $Y=9375
X1731 78 M2M3_PR_DigitalLDOLogic_gds $T=142710 15050 0 0 $X=142545 $Y=14865
X1732 145 M2M3_PR_DigitalLDOLogic_gds $T=142710 18710 0 0 $X=142545 $Y=18525
X1733 140 M2M3_PR_DigitalLDOLogic_gds $T=150530 9560 0 0 $X=150365 $Y=9375
X1734 33 M2M3_PR_DigitalLDOLogic_gds $T=151450 8950 0 0 $X=151285 $Y=8765
X1735 83 M2M3_PR_DigitalLDOLogic_gds $T=153750 18710 0 0 $X=153585 $Y=18525
X1736 83 M2M3_PR_DigitalLDOLogic_gds $T=162030 18710 0 0 $X=161865 $Y=18525
X1737 36 M2M3_PR_DigitalLDOLogic_gds $T=164790 3460 0 0 $X=164625 $Y=3275
X1738 83 M2M3_PR_DigitalLDOLogic_gds $T=164790 18710 0 0 $X=164625 $Y=18525
X1739 112 M2M3_PR_DigitalLDOLogic_gds $T=164790 26030 0 0 $X=164625 $Y=25845
X1740 83 M2M3_PR_DigitalLDOLogic_gds $T=170310 18710 0 0 $X=170145 $Y=18525
X1741 14 M2M3_PR_DigitalLDOLogic_gds $T=170310 22370 0 0 $X=170145 $Y=22185
X1742 38 M2M3_PR_DigitalLDOLogic_gds $T=178590 4070 0 0 $X=178425 $Y=3885
X1743 39 M2M3_PR_DigitalLDOLogic_gds $T=186870 5290 0 0 $X=186705 $Y=5105
X1744 14 M2M3_PR_DigitalLDOLogic_gds $T=189630 1020 0 0 $X=189465 $Y=835
X1745 3 M3M4_PR_DigitalLDOLogic_gds $T=10230 1630 0 0 $X=10040 $Y=1465
X1746 6 M3M4_PR_DigitalLDOLogic_gds $T=23340 1020 0 0 $X=23150 $Y=855
X1747 8 M3M4_PR_DigitalLDOLogic_gds $T=36450 1020 0 0 $X=36260 $Y=855
X1748 12 M3M4_PR_DigitalLDOLogic_gds $T=48870 10170 0 0 $X=48680 $Y=10005
X1749 10 M3M4_PR_DigitalLDOLogic_gds $T=60600 8950 0 0 $X=60410 $Y=8785
X1750 10 M3M4_PR_DigitalLDOLogic_gds $T=60600 13830 0 0 $X=60410 $Y=13665
X1751 15 M3M4_PR_DigitalLDOLogic_gds $T=61980 1020 0 0 $X=61790 $Y=855
X1752 17 M3M4_PR_DigitalLDOLogic_gds $T=74400 3460 0 0 $X=74210 $Y=3295
X1753 18 M3M4_PR_DigitalLDOLogic_gds $T=76470 10780 0 0 $X=76280 $Y=10615
X1754 18 M3M4_PR_DigitalLDOLogic_gds $T=76470 18100 0 0 $X=76280 $Y=17935
X1755 21 M3M4_PR_DigitalLDOLogic_gds $T=87510 10170 0 0 $X=87320 $Y=10005
X1756 23 M3M4_PR_DigitalLDOLogic_gds $T=99930 2850 0 0 $X=99740 $Y=2685
X1757 25 M3M4_PR_DigitalLDOLogic_gds $T=113040 8950 0 0 $X=112850 $Y=8785
X1758 28 M3M4_PR_DigitalLDOLogic_gds $T=126150 14440 0 0 $X=125960 $Y=14275
X1759 31 M3M4_PR_DigitalLDOLogic_gds $T=138570 1020 0 0 $X=138380 $Y=855
X1760 33 M3M4_PR_DigitalLDOLogic_gds $T=151680 8950 0 0 $X=151490 $Y=8785
X1761 36 M3M4_PR_DigitalLDOLogic_gds $T=164100 3460 0 0 $X=163910 $Y=3295
X1762 14 M3M4_PR_DigitalLDOLogic_gds $T=171000 1020 0 0 $X=170810 $Y=855
X1763 14 M3M4_PR_DigitalLDOLogic_gds $T=171000 22370 0 0 $X=170810 $Y=22205
X1764 38 M3M4_PR_DigitalLDOLogic_gds $T=177210 4070 0 0 $X=177020 $Y=3905
X1765 39 M3M4_PR_DigitalLDOLogic_gds $T=189630 5290 0 0 $X=189440 $Y=5125
X1766 2 DigitalLDOLogic_VIA0 $T=11150 12720 0 0 $X=10900 $Y=12480
X1767 2 DigitalLDOLogic_VIA0 $T=11150 18160 0 0 $X=10900 $Y=17920
X1768 2 DigitalLDOLogic_VIA0 $T=11150 23600 0 0 $X=10900 $Y=23360
X1769 2 DigitalLDOLogic_VIA0 $T=11150 29040 0 0 $X=10900 $Y=28800
X1770 2 DigitalLDOLogic_VIA0 $T=11150 34480 0 0 $X=10900 $Y=34240
X1771 2 DigitalLDOLogic_VIA0 $T=11150 39920 0 0 $X=10900 $Y=39680
X1772 2 DigitalLDOLogic_VIA0 $T=11150 45360 0 0 $X=10900 $Y=45120
X1773 2 DigitalLDOLogic_VIA0 $T=11150 50800 0 0 $X=10900 $Y=50560
X1774 2 DigitalLDOLogic_VIA0 $T=11150 56240 0 0 $X=10900 $Y=56000
X1775 1 DigitalLDOLogic_VIA0 $T=12070 15440 0 0 $X=11820 $Y=15200
X1776 1 DigitalLDOLogic_VIA0 $T=12070 20880 0 0 $X=11820 $Y=20640
X1777 1 DigitalLDOLogic_VIA0 $T=12070 26320 0 0 $X=11820 $Y=26080
X1778 1 DigitalLDOLogic_VIA0 $T=12070 31760 0 0 $X=11820 $Y=31520
X1779 1 DigitalLDOLogic_VIA0 $T=12070 37200 0 0 $X=11820 $Y=36960
X1780 1 DigitalLDOLogic_VIA0 $T=12070 42640 0 0 $X=11820 $Y=42400
X1781 1 DigitalLDOLogic_VIA0 $T=12070 48080 0 0 $X=11820 $Y=47840
X1782 1 DigitalLDOLogic_VIA0 $T=12070 53520 0 0 $X=11820 $Y=53280
X1783 1 DigitalLDOLogic_VIA0 $T=12070 58960 0 0 $X=11820 $Y=58720
X1784 2 DigitalLDOLogic_VIA0 $T=13910 12720 0 0 $X=13660 $Y=12480
X1785 2 DigitalLDOLogic_VIA0 $T=13910 18160 0 0 $X=13660 $Y=17920
X1786 2 DigitalLDOLogic_VIA0 $T=13910 23600 0 0 $X=13660 $Y=23360
X1787 2 DigitalLDOLogic_VIA0 $T=13910 29040 0 0 $X=13660 $Y=28800
X1788 2 DigitalLDOLogic_VIA0 $T=13910 34480 0 0 $X=13660 $Y=34240
X1789 2 DigitalLDOLogic_VIA0 $T=13910 39920 0 0 $X=13660 $Y=39680
X1790 2 DigitalLDOLogic_VIA0 $T=13910 45360 0 0 $X=13660 $Y=45120
X1791 2 DigitalLDOLogic_VIA0 $T=13910 50800 0 0 $X=13660 $Y=50560
X1792 2 DigitalLDOLogic_VIA0 $T=13910 56240 0 0 $X=13660 $Y=56000
X1793 1 DigitalLDOLogic_VIA0 $T=14830 15440 0 0 $X=14580 $Y=15200
X1794 1 DigitalLDOLogic_VIA0 $T=14830 20880 0 0 $X=14580 $Y=20640
X1795 1 DigitalLDOLogic_VIA0 $T=14830 26320 0 0 $X=14580 $Y=26080
X1796 1 DigitalLDOLogic_VIA0 $T=14830 31760 0 0 $X=14580 $Y=31520
X1797 1 DigitalLDOLogic_VIA0 $T=14830 37200 0 0 $X=14580 $Y=36960
X1798 1 DigitalLDOLogic_VIA0 $T=14830 42640 0 0 $X=14580 $Y=42400
X1799 1 DigitalLDOLogic_VIA0 $T=14830 48080 0 0 $X=14580 $Y=47840
X1800 1 DigitalLDOLogic_VIA0 $T=14830 53520 0 0 $X=14580 $Y=53280
X1801 1 DigitalLDOLogic_VIA0 $T=14830 58960 0 0 $X=14580 $Y=58720
X1802 2 DigitalLDOLogic_VIA0 $T=16670 12720 0 0 $X=16420 $Y=12480
X1803 2 DigitalLDOLogic_VIA0 $T=16670 18160 0 0 $X=16420 $Y=17920
X1804 2 DigitalLDOLogic_VIA0 $T=16670 23600 0 0 $X=16420 $Y=23360
X1805 2 DigitalLDOLogic_VIA0 $T=16670 29040 0 0 $X=16420 $Y=28800
X1806 2 DigitalLDOLogic_VIA0 $T=16670 34480 0 0 $X=16420 $Y=34240
X1807 2 DigitalLDOLogic_VIA0 $T=16670 39920 0 0 $X=16420 $Y=39680
X1808 2 DigitalLDOLogic_VIA0 $T=16670 45360 0 0 $X=16420 $Y=45120
X1809 2 DigitalLDOLogic_VIA0 $T=16670 50800 0 0 $X=16420 $Y=50560
X1810 2 DigitalLDOLogic_VIA0 $T=16670 56240 0 0 $X=16420 $Y=56000
X1811 1 DigitalLDOLogic_VIA0 $T=17590 15440 0 0 $X=17340 $Y=15200
X1812 1 DigitalLDOLogic_VIA0 $T=17590 20880 0 0 $X=17340 $Y=20640
X1813 1 DigitalLDOLogic_VIA0 $T=17590 26320 0 0 $X=17340 $Y=26080
X1814 1 DigitalLDOLogic_VIA0 $T=17590 31760 0 0 $X=17340 $Y=31520
X1815 1 DigitalLDOLogic_VIA0 $T=17590 37200 0 0 $X=17340 $Y=36960
X1816 1 DigitalLDOLogic_VIA0 $T=17590 42640 0 0 $X=17340 $Y=42400
X1817 1 DigitalLDOLogic_VIA0 $T=17590 48080 0 0 $X=17340 $Y=47840
X1818 1 DigitalLDOLogic_VIA0 $T=17590 53520 0 0 $X=17340 $Y=53280
X1819 1 DigitalLDOLogic_VIA0 $T=17590 58960 0 0 $X=17340 $Y=58720
X1820 2 DigitalLDOLogic_VIA0 $T=19430 12720 0 0 $X=19180 $Y=12480
X1821 2 DigitalLDOLogic_VIA0 $T=19430 18160 0 0 $X=19180 $Y=17920
X1822 2 DigitalLDOLogic_VIA0 $T=19430 23600 0 0 $X=19180 $Y=23360
X1823 2 DigitalLDOLogic_VIA0 $T=19430 29040 0 0 $X=19180 $Y=28800
X1824 2 DigitalLDOLogic_VIA0 $T=19430 34480 0 0 $X=19180 $Y=34240
X1825 2 DigitalLDOLogic_VIA0 $T=19430 39920 0 0 $X=19180 $Y=39680
X1826 2 DigitalLDOLogic_VIA0 $T=19430 45360 0 0 $X=19180 $Y=45120
X1827 2 DigitalLDOLogic_VIA0 $T=19430 50800 0 0 $X=19180 $Y=50560
X1828 2 DigitalLDOLogic_VIA0 $T=19430 56240 0 0 $X=19180 $Y=56000
X1829 1 DigitalLDOLogic_VIA0 $T=20350 15440 0 0 $X=20100 $Y=15200
X1830 1 DigitalLDOLogic_VIA0 $T=20350 20880 0 0 $X=20100 $Y=20640
X1831 1 DigitalLDOLogic_VIA0 $T=20350 26320 0 0 $X=20100 $Y=26080
X1832 1 DigitalLDOLogic_VIA0 $T=20350 31760 0 0 $X=20100 $Y=31520
X1833 1 DigitalLDOLogic_VIA0 $T=20350 37200 0 0 $X=20100 $Y=36960
X1834 1 DigitalLDOLogic_VIA0 $T=20350 42640 0 0 $X=20100 $Y=42400
X1835 1 DigitalLDOLogic_VIA0 $T=20350 48080 0 0 $X=20100 $Y=47840
X1836 1 DigitalLDOLogic_VIA0 $T=20350 53520 0 0 $X=20100 $Y=53280
X1837 1 DigitalLDOLogic_VIA0 $T=20350 58960 0 0 $X=20100 $Y=58720
X1838 2 DigitalLDOLogic_VIA0 $T=22190 12720 0 0 $X=21940 $Y=12480
X1839 2 DigitalLDOLogic_VIA0 $T=22190 18160 0 0 $X=21940 $Y=17920
X1840 2 DigitalLDOLogic_VIA0 $T=22190 23600 0 0 $X=21940 $Y=23360
X1841 2 DigitalLDOLogic_VIA0 $T=22190 29040 0 0 $X=21940 $Y=28800
X1842 2 DigitalLDOLogic_VIA0 $T=22190 34480 0 0 $X=21940 $Y=34240
X1843 2 DigitalLDOLogic_VIA0 $T=22190 39920 0 0 $X=21940 $Y=39680
X1844 2 DigitalLDOLogic_VIA0 $T=22190 45360 0 0 $X=21940 $Y=45120
X1845 2 DigitalLDOLogic_VIA0 $T=22190 50800 0 0 $X=21940 $Y=50560
X1846 2 DigitalLDOLogic_VIA0 $T=22190 56240 0 0 $X=21940 $Y=56000
X1847 1 DigitalLDOLogic_VIA0 $T=23110 15440 0 0 $X=22860 $Y=15200
X1848 1 DigitalLDOLogic_VIA0 $T=23110 20880 0 0 $X=22860 $Y=20640
X1849 1 DigitalLDOLogic_VIA0 $T=23110 26320 0 0 $X=22860 $Y=26080
X1850 1 DigitalLDOLogic_VIA0 $T=23110 31760 0 0 $X=22860 $Y=31520
X1851 1 DigitalLDOLogic_VIA0 $T=23110 37200 0 0 $X=22860 $Y=36960
X1852 1 DigitalLDOLogic_VIA0 $T=23110 42640 0 0 $X=22860 $Y=42400
X1853 1 DigitalLDOLogic_VIA0 $T=23110 48080 0 0 $X=22860 $Y=47840
X1854 1 DigitalLDOLogic_VIA0 $T=23110 53520 0 0 $X=22860 $Y=53280
X1855 1 DigitalLDOLogic_VIA0 $T=23110 58960 0 0 $X=22860 $Y=58720
X1856 2 DigitalLDOLogic_VIA0 $T=24950 12720 0 0 $X=24700 $Y=12480
X1857 2 DigitalLDOLogic_VIA0 $T=24950 18160 0 0 $X=24700 $Y=17920
X1858 2 DigitalLDOLogic_VIA0 $T=24950 23600 0 0 $X=24700 $Y=23360
X1859 2 DigitalLDOLogic_VIA0 $T=24950 29040 0 0 $X=24700 $Y=28800
X1860 2 DigitalLDOLogic_VIA0 $T=24950 34480 0 0 $X=24700 $Y=34240
X1861 2 DigitalLDOLogic_VIA0 $T=24950 39920 0 0 $X=24700 $Y=39680
X1862 2 DigitalLDOLogic_VIA0 $T=24950 45360 0 0 $X=24700 $Y=45120
X1863 2 DigitalLDOLogic_VIA0 $T=24950 50800 0 0 $X=24700 $Y=50560
X1864 2 DigitalLDOLogic_VIA0 $T=24950 56240 0 0 $X=24700 $Y=56000
X1865 1 DigitalLDOLogic_VIA0 $T=25870 15440 0 0 $X=25620 $Y=15200
X1866 1 DigitalLDOLogic_VIA0 $T=25870 20880 0 0 $X=25620 $Y=20640
X1867 1 DigitalLDOLogic_VIA0 $T=25870 26320 0 0 $X=25620 $Y=26080
X1868 1 DigitalLDOLogic_VIA0 $T=25870 31760 0 0 $X=25620 $Y=31520
X1869 1 DigitalLDOLogic_VIA0 $T=25870 37200 0 0 $X=25620 $Y=36960
X1870 1 DigitalLDOLogic_VIA0 $T=25870 42640 0 0 $X=25620 $Y=42400
X1871 1 DigitalLDOLogic_VIA0 $T=25870 48080 0 0 $X=25620 $Y=47840
X1872 1 DigitalLDOLogic_VIA0 $T=25870 53520 0 0 $X=25620 $Y=53280
X1873 1 DigitalLDOLogic_VIA0 $T=25870 58960 0 0 $X=25620 $Y=58720
X1874 2 DigitalLDOLogic_VIA0 $T=27710 12720 0 0 $X=27460 $Y=12480
X1875 2 DigitalLDOLogic_VIA0 $T=27710 18160 0 0 $X=27460 $Y=17920
X1876 2 DigitalLDOLogic_VIA0 $T=27710 23600 0 0 $X=27460 $Y=23360
X1877 2 DigitalLDOLogic_VIA0 $T=27710 29040 0 0 $X=27460 $Y=28800
X1878 2 DigitalLDOLogic_VIA0 $T=27710 34480 0 0 $X=27460 $Y=34240
X1879 2 DigitalLDOLogic_VIA0 $T=27710 39920 0 0 $X=27460 $Y=39680
X1880 2 DigitalLDOLogic_VIA0 $T=27710 45360 0 0 $X=27460 $Y=45120
X1881 2 DigitalLDOLogic_VIA0 $T=27710 50800 0 0 $X=27460 $Y=50560
X1882 2 DigitalLDOLogic_VIA0 $T=27710 56240 0 0 $X=27460 $Y=56000
X1883 1 DigitalLDOLogic_VIA0 $T=28630 15440 0 0 $X=28380 $Y=15200
X1884 1 DigitalLDOLogic_VIA0 $T=28630 20880 0 0 $X=28380 $Y=20640
X1885 1 DigitalLDOLogic_VIA0 $T=28630 26320 0 0 $X=28380 $Y=26080
X1886 1 DigitalLDOLogic_VIA0 $T=28630 31760 0 0 $X=28380 $Y=31520
X1887 1 DigitalLDOLogic_VIA0 $T=28630 37200 0 0 $X=28380 $Y=36960
X1888 1 DigitalLDOLogic_VIA0 $T=28630 42640 0 0 $X=28380 $Y=42400
X1889 1 DigitalLDOLogic_VIA0 $T=28630 48080 0 0 $X=28380 $Y=47840
X1890 1 DigitalLDOLogic_VIA0 $T=28630 53520 0 0 $X=28380 $Y=53280
X1891 1 DigitalLDOLogic_VIA0 $T=28630 58960 0 0 $X=28380 $Y=58720
X1892 2 DigitalLDOLogic_VIA0 $T=30470 12720 0 0 $X=30220 $Y=12480
X1893 2 DigitalLDOLogic_VIA0 $T=30470 18160 0 0 $X=30220 $Y=17920
X1894 2 DigitalLDOLogic_VIA0 $T=30470 23600 0 0 $X=30220 $Y=23360
X1895 2 DigitalLDOLogic_VIA0 $T=30470 29040 0 0 $X=30220 $Y=28800
X1896 2 DigitalLDOLogic_VIA0 $T=30470 34480 0 0 $X=30220 $Y=34240
X1897 2 DigitalLDOLogic_VIA0 $T=30470 39920 0 0 $X=30220 $Y=39680
X1898 2 DigitalLDOLogic_VIA0 $T=30470 45360 0 0 $X=30220 $Y=45120
X1899 2 DigitalLDOLogic_VIA0 $T=30470 50800 0 0 $X=30220 $Y=50560
X1900 2 DigitalLDOLogic_VIA0 $T=30470 56240 0 0 $X=30220 $Y=56000
X1901 1 DigitalLDOLogic_VIA0 $T=31390 15440 0 0 $X=31140 $Y=15200
X1902 1 DigitalLDOLogic_VIA0 $T=31390 20880 0 0 $X=31140 $Y=20640
X1903 1 DigitalLDOLogic_VIA0 $T=31390 26320 0 0 $X=31140 $Y=26080
X1904 1 DigitalLDOLogic_VIA0 $T=31390 31760 0 0 $X=31140 $Y=31520
X1905 1 DigitalLDOLogic_VIA0 $T=31390 37200 0 0 $X=31140 $Y=36960
X1906 1 DigitalLDOLogic_VIA0 $T=31390 42640 0 0 $X=31140 $Y=42400
X1907 1 DigitalLDOLogic_VIA0 $T=31390 48080 0 0 $X=31140 $Y=47840
X1908 1 DigitalLDOLogic_VIA0 $T=31390 53520 0 0 $X=31140 $Y=53280
X1909 1 DigitalLDOLogic_VIA0 $T=31390 58960 0 0 $X=31140 $Y=58720
X1910 2 DigitalLDOLogic_VIA0 $T=33230 12720 0 0 $X=32980 $Y=12480
X1911 2 DigitalLDOLogic_VIA0 $T=33230 18160 0 0 $X=32980 $Y=17920
X1912 2 DigitalLDOLogic_VIA0 $T=33230 23600 0 0 $X=32980 $Y=23360
X1913 2 DigitalLDOLogic_VIA0 $T=33230 29040 0 0 $X=32980 $Y=28800
X1914 2 DigitalLDOLogic_VIA0 $T=33230 34480 0 0 $X=32980 $Y=34240
X1915 2 DigitalLDOLogic_VIA0 $T=33230 39920 0 0 $X=32980 $Y=39680
X1916 2 DigitalLDOLogic_VIA0 $T=33230 45360 0 0 $X=32980 $Y=45120
X1917 2 DigitalLDOLogic_VIA0 $T=33230 50800 0 0 $X=32980 $Y=50560
X1918 2 DigitalLDOLogic_VIA0 $T=33230 56240 0 0 $X=32980 $Y=56000
X1919 1 DigitalLDOLogic_VIA0 $T=34150 15440 0 0 $X=33900 $Y=15200
X1920 1 DigitalLDOLogic_VIA0 $T=34150 20880 0 0 $X=33900 $Y=20640
X1921 1 DigitalLDOLogic_VIA0 $T=34150 26320 0 0 $X=33900 $Y=26080
X1922 1 DigitalLDOLogic_VIA0 $T=34150 31760 0 0 $X=33900 $Y=31520
X1923 1 DigitalLDOLogic_VIA0 $T=34150 37200 0 0 $X=33900 $Y=36960
X1924 1 DigitalLDOLogic_VIA0 $T=34150 42640 0 0 $X=33900 $Y=42400
X1925 1 DigitalLDOLogic_VIA0 $T=34150 48080 0 0 $X=33900 $Y=47840
X1926 1 DigitalLDOLogic_VIA0 $T=34150 53520 0 0 $X=33900 $Y=53280
X1927 1 DigitalLDOLogic_VIA0 $T=34150 58960 0 0 $X=33900 $Y=58720
X1928 2 DigitalLDOLogic_VIA0 $T=35990 12720 0 0 $X=35740 $Y=12480
X1929 2 DigitalLDOLogic_VIA0 $T=35990 18160 0 0 $X=35740 $Y=17920
X1930 2 DigitalLDOLogic_VIA0 $T=35990 23600 0 0 $X=35740 $Y=23360
X1931 2 DigitalLDOLogic_VIA0 $T=35990 29040 0 0 $X=35740 $Y=28800
X1932 2 DigitalLDOLogic_VIA0 $T=35990 34480 0 0 $X=35740 $Y=34240
X1933 2 DigitalLDOLogic_VIA0 $T=35990 39920 0 0 $X=35740 $Y=39680
X1934 2 DigitalLDOLogic_VIA0 $T=35990 45360 0 0 $X=35740 $Y=45120
X1935 2 DigitalLDOLogic_VIA0 $T=35990 50800 0 0 $X=35740 $Y=50560
X1936 2 DigitalLDOLogic_VIA0 $T=35990 56240 0 0 $X=35740 $Y=56000
X1937 1 DigitalLDOLogic_VIA0 $T=36910 15440 0 0 $X=36660 $Y=15200
X1938 1 DigitalLDOLogic_VIA0 $T=36910 20880 0 0 $X=36660 $Y=20640
X1939 1 DigitalLDOLogic_VIA0 $T=36910 26320 0 0 $X=36660 $Y=26080
X1940 1 DigitalLDOLogic_VIA0 $T=36910 31760 0 0 $X=36660 $Y=31520
X1941 1 DigitalLDOLogic_VIA0 $T=36910 37200 0 0 $X=36660 $Y=36960
X1942 1 DigitalLDOLogic_VIA0 $T=36910 42640 0 0 $X=36660 $Y=42400
X1943 1 DigitalLDOLogic_VIA0 $T=36910 48080 0 0 $X=36660 $Y=47840
X1944 1 DigitalLDOLogic_VIA0 $T=36910 53520 0 0 $X=36660 $Y=53280
X1945 1 DigitalLDOLogic_VIA0 $T=36910 58960 0 0 $X=36660 $Y=58720
X1946 2 DigitalLDOLogic_VIA0 $T=38750 12720 0 0 $X=38500 $Y=12480
X1947 2 DigitalLDOLogic_VIA0 $T=38750 18160 0 0 $X=38500 $Y=17920
X1948 2 DigitalLDOLogic_VIA0 $T=38750 23600 0 0 $X=38500 $Y=23360
X1949 2 DigitalLDOLogic_VIA0 $T=38750 29040 0 0 $X=38500 $Y=28800
X1950 2 DigitalLDOLogic_VIA0 $T=38750 34480 0 0 $X=38500 $Y=34240
X1951 2 DigitalLDOLogic_VIA0 $T=38750 39920 0 0 $X=38500 $Y=39680
X1952 2 DigitalLDOLogic_VIA0 $T=38750 45360 0 0 $X=38500 $Y=45120
X1953 2 DigitalLDOLogic_VIA0 $T=38750 50800 0 0 $X=38500 $Y=50560
X1954 2 DigitalLDOLogic_VIA0 $T=38750 56240 0 0 $X=38500 $Y=56000
X1955 1 DigitalLDOLogic_VIA0 $T=39670 15440 0 0 $X=39420 $Y=15200
X1956 1 DigitalLDOLogic_VIA0 $T=39670 20880 0 0 $X=39420 $Y=20640
X1957 1 DigitalLDOLogic_VIA0 $T=39670 26320 0 0 $X=39420 $Y=26080
X1958 1 DigitalLDOLogic_VIA0 $T=39670 31760 0 0 $X=39420 $Y=31520
X1959 1 DigitalLDOLogic_VIA0 $T=39670 37200 0 0 $X=39420 $Y=36960
X1960 1 DigitalLDOLogic_VIA0 $T=39670 42640 0 0 $X=39420 $Y=42400
X1961 1 DigitalLDOLogic_VIA0 $T=39670 48080 0 0 $X=39420 $Y=47840
X1962 1 DigitalLDOLogic_VIA0 $T=39670 53520 0 0 $X=39420 $Y=53280
X1963 1 DigitalLDOLogic_VIA0 $T=39670 58960 0 0 $X=39420 $Y=58720
X1964 2 DigitalLDOLogic_VIA0 $T=41510 12720 0 0 $X=41260 $Y=12480
X1965 2 DigitalLDOLogic_VIA0 $T=41510 18160 0 0 $X=41260 $Y=17920
X1966 2 DigitalLDOLogic_VIA0 $T=41510 23600 0 0 $X=41260 $Y=23360
X1967 2 DigitalLDOLogic_VIA0 $T=41510 29040 0 0 $X=41260 $Y=28800
X1968 2 DigitalLDOLogic_VIA0 $T=41510 34480 0 0 $X=41260 $Y=34240
X1969 2 DigitalLDOLogic_VIA0 $T=41510 39920 0 0 $X=41260 $Y=39680
X1970 2 DigitalLDOLogic_VIA0 $T=41510 45360 0 0 $X=41260 $Y=45120
X1971 2 DigitalLDOLogic_VIA0 $T=41510 50800 0 0 $X=41260 $Y=50560
X1972 2 DigitalLDOLogic_VIA0 $T=41510 56240 0 0 $X=41260 $Y=56000
X1973 1 DigitalLDOLogic_VIA0 $T=42430 15440 0 0 $X=42180 $Y=15200
X1974 1 DigitalLDOLogic_VIA0 $T=42430 20880 0 0 $X=42180 $Y=20640
X1975 1 DigitalLDOLogic_VIA0 $T=42430 26320 0 0 $X=42180 $Y=26080
X1976 1 DigitalLDOLogic_VIA0 $T=42430 31760 0 0 $X=42180 $Y=31520
X1977 1 DigitalLDOLogic_VIA0 $T=42430 37200 0 0 $X=42180 $Y=36960
X1978 1 DigitalLDOLogic_VIA0 $T=42430 42640 0 0 $X=42180 $Y=42400
X1979 1 DigitalLDOLogic_VIA0 $T=42430 48080 0 0 $X=42180 $Y=47840
X1980 1 DigitalLDOLogic_VIA0 $T=42430 53520 0 0 $X=42180 $Y=53280
X1981 1 DigitalLDOLogic_VIA0 $T=42430 58960 0 0 $X=42180 $Y=58720
X1982 2 DigitalLDOLogic_VIA0 $T=44270 12720 0 0 $X=44020 $Y=12480
X1983 2 DigitalLDOLogic_VIA0 $T=44270 18160 0 0 $X=44020 $Y=17920
X1984 2 DigitalLDOLogic_VIA0 $T=44270 23600 0 0 $X=44020 $Y=23360
X1985 2 DigitalLDOLogic_VIA0 $T=44270 29040 0 0 $X=44020 $Y=28800
X1986 2 DigitalLDOLogic_VIA0 $T=44270 34480 0 0 $X=44020 $Y=34240
X1987 2 DigitalLDOLogic_VIA0 $T=44270 39920 0 0 $X=44020 $Y=39680
X1988 2 DigitalLDOLogic_VIA0 $T=44270 45360 0 0 $X=44020 $Y=45120
X1989 2 DigitalLDOLogic_VIA0 $T=44270 50800 0 0 $X=44020 $Y=50560
X1990 2 DigitalLDOLogic_VIA0 $T=44270 56240 0 0 $X=44020 $Y=56000
X1991 1 DigitalLDOLogic_VIA0 $T=45190 15440 0 0 $X=44940 $Y=15200
X1992 1 DigitalLDOLogic_VIA0 $T=45190 20880 0 0 $X=44940 $Y=20640
X1993 1 DigitalLDOLogic_VIA0 $T=45190 26320 0 0 $X=44940 $Y=26080
X1994 1 DigitalLDOLogic_VIA0 $T=45190 31760 0 0 $X=44940 $Y=31520
X1995 1 DigitalLDOLogic_VIA0 $T=45190 37200 0 0 $X=44940 $Y=36960
X1996 1 DigitalLDOLogic_VIA0 $T=45190 42640 0 0 $X=44940 $Y=42400
X1997 1 DigitalLDOLogic_VIA0 $T=45190 48080 0 0 $X=44940 $Y=47840
X1998 1 DigitalLDOLogic_VIA0 $T=45190 53520 0 0 $X=44940 $Y=53280
X1999 1 DigitalLDOLogic_VIA0 $T=45190 58960 0 0 $X=44940 $Y=58720
X2000 2 DigitalLDOLogic_VIA0 $T=47030 12720 0 0 $X=46780 $Y=12480
X2001 2 DigitalLDOLogic_VIA0 $T=47030 18160 0 0 $X=46780 $Y=17920
X2002 2 DigitalLDOLogic_VIA0 $T=47030 23600 0 0 $X=46780 $Y=23360
X2003 2 DigitalLDOLogic_VIA0 $T=47030 29040 0 0 $X=46780 $Y=28800
X2004 2 DigitalLDOLogic_VIA0 $T=47030 34480 0 0 $X=46780 $Y=34240
X2005 2 DigitalLDOLogic_VIA0 $T=47030 39920 0 0 $X=46780 $Y=39680
X2006 2 DigitalLDOLogic_VIA0 $T=47030 45360 0 0 $X=46780 $Y=45120
X2007 2 DigitalLDOLogic_VIA0 $T=47030 50800 0 0 $X=46780 $Y=50560
X2008 2 DigitalLDOLogic_VIA0 $T=47030 56240 0 0 $X=46780 $Y=56000
X2009 1 DigitalLDOLogic_VIA0 $T=47950 15440 0 0 $X=47700 $Y=15200
X2010 1 DigitalLDOLogic_VIA0 $T=47950 20880 0 0 $X=47700 $Y=20640
X2011 1 DigitalLDOLogic_VIA0 $T=47950 26320 0 0 $X=47700 $Y=26080
X2012 1 DigitalLDOLogic_VIA0 $T=47950 31760 0 0 $X=47700 $Y=31520
X2013 1 DigitalLDOLogic_VIA0 $T=47950 37200 0 0 $X=47700 $Y=36960
X2014 1 DigitalLDOLogic_VIA0 $T=47950 42640 0 0 $X=47700 $Y=42400
X2015 1 DigitalLDOLogic_VIA0 $T=47950 48080 0 0 $X=47700 $Y=47840
X2016 1 DigitalLDOLogic_VIA0 $T=47950 53520 0 0 $X=47700 $Y=53280
X2017 1 DigitalLDOLogic_VIA0 $T=47950 58960 0 0 $X=47700 $Y=58720
X2018 2 DigitalLDOLogic_VIA0 $T=49790 12720 0 0 $X=49540 $Y=12480
X2019 2 DigitalLDOLogic_VIA0 $T=49790 18160 0 0 $X=49540 $Y=17920
X2020 2 DigitalLDOLogic_VIA0 $T=49790 23600 0 0 $X=49540 $Y=23360
X2021 2 DigitalLDOLogic_VIA0 $T=49790 29040 0 0 $X=49540 $Y=28800
X2022 2 DigitalLDOLogic_VIA0 $T=49790 34480 0 0 $X=49540 $Y=34240
X2023 2 DigitalLDOLogic_VIA0 $T=49790 39920 0 0 $X=49540 $Y=39680
X2024 2 DigitalLDOLogic_VIA0 $T=49790 45360 0 0 $X=49540 $Y=45120
X2025 2 DigitalLDOLogic_VIA0 $T=49790 50800 0 0 $X=49540 $Y=50560
X2026 2 DigitalLDOLogic_VIA0 $T=49790 56240 0 0 $X=49540 $Y=56000
X2027 1 DigitalLDOLogic_VIA0 $T=50710 15440 0 0 $X=50460 $Y=15200
X2028 1 DigitalLDOLogic_VIA0 $T=50710 20880 0 0 $X=50460 $Y=20640
X2029 1 DigitalLDOLogic_VIA0 $T=50710 26320 0 0 $X=50460 $Y=26080
X2030 1 DigitalLDOLogic_VIA0 $T=50710 31760 0 0 $X=50460 $Y=31520
X2031 1 DigitalLDOLogic_VIA0 $T=50710 37200 0 0 $X=50460 $Y=36960
X2032 1 DigitalLDOLogic_VIA0 $T=50710 42640 0 0 $X=50460 $Y=42400
X2033 1 DigitalLDOLogic_VIA0 $T=50710 48080 0 0 $X=50460 $Y=47840
X2034 1 DigitalLDOLogic_VIA0 $T=50710 53520 0 0 $X=50460 $Y=53280
X2035 1 DigitalLDOLogic_VIA0 $T=50710 58960 0 0 $X=50460 $Y=58720
X2036 2 DigitalLDOLogic_VIA0 $T=52550 12720 0 0 $X=52300 $Y=12480
X2037 2 DigitalLDOLogic_VIA0 $T=52550 18160 0 0 $X=52300 $Y=17920
X2038 2 DigitalLDOLogic_VIA0 $T=52550 23600 0 0 $X=52300 $Y=23360
X2039 2 DigitalLDOLogic_VIA0 $T=52550 29040 0 0 $X=52300 $Y=28800
X2040 2 DigitalLDOLogic_VIA0 $T=52550 34480 0 0 $X=52300 $Y=34240
X2041 2 DigitalLDOLogic_VIA0 $T=52550 39920 0 0 $X=52300 $Y=39680
X2042 2 DigitalLDOLogic_VIA0 $T=52550 45360 0 0 $X=52300 $Y=45120
X2043 2 DigitalLDOLogic_VIA0 $T=52550 50800 0 0 $X=52300 $Y=50560
X2044 2 DigitalLDOLogic_VIA0 $T=52550 56240 0 0 $X=52300 $Y=56000
X2045 1 DigitalLDOLogic_VIA0 $T=53470 15440 0 0 $X=53220 $Y=15200
X2046 1 DigitalLDOLogic_VIA0 $T=53470 20880 0 0 $X=53220 $Y=20640
X2047 1 DigitalLDOLogic_VIA0 $T=53470 26320 0 0 $X=53220 $Y=26080
X2048 1 DigitalLDOLogic_VIA0 $T=53470 31760 0 0 $X=53220 $Y=31520
X2049 1 DigitalLDOLogic_VIA0 $T=53470 37200 0 0 $X=53220 $Y=36960
X2050 1 DigitalLDOLogic_VIA0 $T=53470 42640 0 0 $X=53220 $Y=42400
X2051 1 DigitalLDOLogic_VIA0 $T=53470 48080 0 0 $X=53220 $Y=47840
X2052 1 DigitalLDOLogic_VIA0 $T=53470 53520 0 0 $X=53220 $Y=53280
X2053 1 DigitalLDOLogic_VIA0 $T=53470 58960 0 0 $X=53220 $Y=58720
X2054 2 DigitalLDOLogic_VIA0 $T=55310 12720 0 0 $X=55060 $Y=12480
X2055 2 DigitalLDOLogic_VIA0 $T=55310 18160 0 0 $X=55060 $Y=17920
X2056 2 DigitalLDOLogic_VIA0 $T=55310 23600 0 0 $X=55060 $Y=23360
X2057 2 DigitalLDOLogic_VIA0 $T=55310 29040 0 0 $X=55060 $Y=28800
X2058 2 DigitalLDOLogic_VIA0 $T=55310 34480 0 0 $X=55060 $Y=34240
X2059 2 DigitalLDOLogic_VIA0 $T=55310 39920 0 0 $X=55060 $Y=39680
X2060 2 DigitalLDOLogic_VIA0 $T=55310 45360 0 0 $X=55060 $Y=45120
X2061 2 DigitalLDOLogic_VIA0 $T=55310 50800 0 0 $X=55060 $Y=50560
X2062 2 DigitalLDOLogic_VIA0 $T=55310 56240 0 0 $X=55060 $Y=56000
X2063 1 DigitalLDOLogic_VIA0 $T=56230 15440 0 0 $X=55980 $Y=15200
X2064 1 DigitalLDOLogic_VIA0 $T=56230 20880 0 0 $X=55980 $Y=20640
X2065 1 DigitalLDOLogic_VIA0 $T=56230 26320 0 0 $X=55980 $Y=26080
X2066 1 DigitalLDOLogic_VIA0 $T=56230 31760 0 0 $X=55980 $Y=31520
X2067 1 DigitalLDOLogic_VIA0 $T=56230 37200 0 0 $X=55980 $Y=36960
X2068 1 DigitalLDOLogic_VIA0 $T=56230 42640 0 0 $X=55980 $Y=42400
X2069 1 DigitalLDOLogic_VIA0 $T=56230 48080 0 0 $X=55980 $Y=47840
X2070 1 DigitalLDOLogic_VIA0 $T=56230 53520 0 0 $X=55980 $Y=53280
X2071 1 DigitalLDOLogic_VIA0 $T=56230 58960 0 0 $X=55980 $Y=58720
X2072 2 DigitalLDOLogic_VIA0 $T=58070 12720 0 0 $X=57820 $Y=12480
X2073 2 DigitalLDOLogic_VIA0 $T=58070 18160 0 0 $X=57820 $Y=17920
X2074 2 DigitalLDOLogic_VIA0 $T=58070 23600 0 0 $X=57820 $Y=23360
X2075 2 DigitalLDOLogic_VIA0 $T=58070 29040 0 0 $X=57820 $Y=28800
X2076 2 DigitalLDOLogic_VIA0 $T=58070 34480 0 0 $X=57820 $Y=34240
X2077 2 DigitalLDOLogic_VIA0 $T=58070 39920 0 0 $X=57820 $Y=39680
X2078 2 DigitalLDOLogic_VIA0 $T=58070 45360 0 0 $X=57820 $Y=45120
X2079 2 DigitalLDOLogic_VIA0 $T=58070 50800 0 0 $X=57820 $Y=50560
X2080 2 DigitalLDOLogic_VIA0 $T=58070 56240 0 0 $X=57820 $Y=56000
X2081 1 DigitalLDOLogic_VIA0 $T=58990 15440 0 0 $X=58740 $Y=15200
X2082 1 DigitalLDOLogic_VIA0 $T=58990 20880 0 0 $X=58740 $Y=20640
X2083 1 DigitalLDOLogic_VIA0 $T=58990 26320 0 0 $X=58740 $Y=26080
X2084 1 DigitalLDOLogic_VIA0 $T=58990 31760 0 0 $X=58740 $Y=31520
X2085 1 DigitalLDOLogic_VIA0 $T=58990 37200 0 0 $X=58740 $Y=36960
X2086 1 DigitalLDOLogic_VIA0 $T=58990 42640 0 0 $X=58740 $Y=42400
X2087 1 DigitalLDOLogic_VIA0 $T=58990 48080 0 0 $X=58740 $Y=47840
X2088 1 DigitalLDOLogic_VIA0 $T=58990 53520 0 0 $X=58740 $Y=53280
X2089 1 DigitalLDOLogic_VIA0 $T=58990 58960 0 0 $X=58740 $Y=58720
X2090 2 DigitalLDOLogic_VIA0 $T=60830 12720 0 0 $X=60580 $Y=12480
X2091 2 DigitalLDOLogic_VIA0 $T=60830 18160 0 0 $X=60580 $Y=17920
X2092 2 DigitalLDOLogic_VIA0 $T=60830 23600 0 0 $X=60580 $Y=23360
X2093 2 DigitalLDOLogic_VIA0 $T=60830 29040 0 0 $X=60580 $Y=28800
X2094 2 DigitalLDOLogic_VIA0 $T=60830 34480 0 0 $X=60580 $Y=34240
X2095 2 DigitalLDOLogic_VIA0 $T=60830 39920 0 0 $X=60580 $Y=39680
X2096 2 DigitalLDOLogic_VIA0 $T=60830 45360 0 0 $X=60580 $Y=45120
X2097 2 DigitalLDOLogic_VIA0 $T=60830 50800 0 0 $X=60580 $Y=50560
X2098 2 DigitalLDOLogic_VIA0 $T=60830 56240 0 0 $X=60580 $Y=56000
X2099 1 DigitalLDOLogic_VIA0 $T=61750 15440 0 0 $X=61500 $Y=15200
X2100 1 DigitalLDOLogic_VIA0 $T=61750 20880 0 0 $X=61500 $Y=20640
X2101 1 DigitalLDOLogic_VIA0 $T=61750 26320 0 0 $X=61500 $Y=26080
X2102 1 DigitalLDOLogic_VIA0 $T=61750 31760 0 0 $X=61500 $Y=31520
X2103 1 DigitalLDOLogic_VIA0 $T=61750 37200 0 0 $X=61500 $Y=36960
X2104 1 DigitalLDOLogic_VIA0 $T=61750 42640 0 0 $X=61500 $Y=42400
X2105 1 DigitalLDOLogic_VIA0 $T=61750 48080 0 0 $X=61500 $Y=47840
X2106 1 DigitalLDOLogic_VIA0 $T=61750 53520 0 0 $X=61500 $Y=53280
X2107 1 DigitalLDOLogic_VIA0 $T=61750 58960 0 0 $X=61500 $Y=58720
X2108 2 DigitalLDOLogic_VIA0 $T=63590 12720 0 0 $X=63340 $Y=12480
X2109 2 DigitalLDOLogic_VIA0 $T=63590 18160 0 0 $X=63340 $Y=17920
X2110 2 DigitalLDOLogic_VIA0 $T=63590 23600 0 0 $X=63340 $Y=23360
X2111 2 DigitalLDOLogic_VIA0 $T=63590 29040 0 0 $X=63340 $Y=28800
X2112 2 DigitalLDOLogic_VIA0 $T=63590 34480 0 0 $X=63340 $Y=34240
X2113 2 DigitalLDOLogic_VIA0 $T=63590 39920 0 0 $X=63340 $Y=39680
X2114 2 DigitalLDOLogic_VIA0 $T=63590 45360 0 0 $X=63340 $Y=45120
X2115 2 DigitalLDOLogic_VIA0 $T=63590 50800 0 0 $X=63340 $Y=50560
X2116 2 DigitalLDOLogic_VIA0 $T=63590 56240 0 0 $X=63340 $Y=56000
X2117 1 DigitalLDOLogic_VIA0 $T=64510 15440 0 0 $X=64260 $Y=15200
X2118 1 DigitalLDOLogic_VIA0 $T=64510 20880 0 0 $X=64260 $Y=20640
X2119 1 DigitalLDOLogic_VIA0 $T=64510 26320 0 0 $X=64260 $Y=26080
X2120 1 DigitalLDOLogic_VIA0 $T=64510 31760 0 0 $X=64260 $Y=31520
X2121 1 DigitalLDOLogic_VIA0 $T=64510 37200 0 0 $X=64260 $Y=36960
X2122 1 DigitalLDOLogic_VIA0 $T=64510 42640 0 0 $X=64260 $Y=42400
X2123 1 DigitalLDOLogic_VIA0 $T=64510 48080 0 0 $X=64260 $Y=47840
X2124 1 DigitalLDOLogic_VIA0 $T=64510 53520 0 0 $X=64260 $Y=53280
X2125 1 DigitalLDOLogic_VIA0 $T=64510 58960 0 0 $X=64260 $Y=58720
X2126 2 DigitalLDOLogic_VIA0 $T=66350 12720 0 0 $X=66100 $Y=12480
X2127 2 DigitalLDOLogic_VIA0 $T=66350 18160 0 0 $X=66100 $Y=17920
X2128 2 DigitalLDOLogic_VIA0 $T=66350 23600 0 0 $X=66100 $Y=23360
X2129 2 DigitalLDOLogic_VIA0 $T=66350 29040 0 0 $X=66100 $Y=28800
X2130 2 DigitalLDOLogic_VIA0 $T=66350 34480 0 0 $X=66100 $Y=34240
X2131 2 DigitalLDOLogic_VIA0 $T=66350 39920 0 0 $X=66100 $Y=39680
X2132 2 DigitalLDOLogic_VIA0 $T=66350 45360 0 0 $X=66100 $Y=45120
X2133 2 DigitalLDOLogic_VIA0 $T=66350 50800 0 0 $X=66100 $Y=50560
X2134 2 DigitalLDOLogic_VIA0 $T=66350 56240 0 0 $X=66100 $Y=56000
X2135 1 DigitalLDOLogic_VIA0 $T=67270 15440 0 0 $X=67020 $Y=15200
X2136 1 DigitalLDOLogic_VIA0 $T=67270 20880 0 0 $X=67020 $Y=20640
X2137 1 DigitalLDOLogic_VIA0 $T=67270 26320 0 0 $X=67020 $Y=26080
X2138 1 DigitalLDOLogic_VIA0 $T=67270 31760 0 0 $X=67020 $Y=31520
X2139 1 DigitalLDOLogic_VIA0 $T=67270 37200 0 0 $X=67020 $Y=36960
X2140 1 DigitalLDOLogic_VIA0 $T=67270 42640 0 0 $X=67020 $Y=42400
X2141 1 DigitalLDOLogic_VIA0 $T=67270 48080 0 0 $X=67020 $Y=47840
X2142 1 DigitalLDOLogic_VIA0 $T=67270 53520 0 0 $X=67020 $Y=53280
X2143 1 DigitalLDOLogic_VIA0 $T=67270 58960 0 0 $X=67020 $Y=58720
X2144 2 DigitalLDOLogic_VIA0 $T=69110 12720 0 0 $X=68860 $Y=12480
X2145 2 DigitalLDOLogic_VIA0 $T=69110 18160 0 0 $X=68860 $Y=17920
X2146 2 DigitalLDOLogic_VIA0 $T=69110 23600 0 0 $X=68860 $Y=23360
X2147 2 DigitalLDOLogic_VIA0 $T=69110 29040 0 0 $X=68860 $Y=28800
X2148 2 DigitalLDOLogic_VIA0 $T=69110 34480 0 0 $X=68860 $Y=34240
X2149 2 DigitalLDOLogic_VIA0 $T=69110 39920 0 0 $X=68860 $Y=39680
X2150 2 DigitalLDOLogic_VIA0 $T=69110 45360 0 0 $X=68860 $Y=45120
X2151 2 DigitalLDOLogic_VIA0 $T=69110 50800 0 0 $X=68860 $Y=50560
X2152 2 DigitalLDOLogic_VIA0 $T=69110 56240 0 0 $X=68860 $Y=56000
X2153 1 DigitalLDOLogic_VIA0 $T=70030 15440 0 0 $X=69780 $Y=15200
X2154 1 DigitalLDOLogic_VIA0 $T=70030 20880 0 0 $X=69780 $Y=20640
X2155 1 DigitalLDOLogic_VIA0 $T=70030 26320 0 0 $X=69780 $Y=26080
X2156 1 DigitalLDOLogic_VIA0 $T=70030 31760 0 0 $X=69780 $Y=31520
X2157 1 DigitalLDOLogic_VIA0 $T=70030 37200 0 0 $X=69780 $Y=36960
X2158 1 DigitalLDOLogic_VIA0 $T=70030 42640 0 0 $X=69780 $Y=42400
X2159 1 DigitalLDOLogic_VIA0 $T=70030 48080 0 0 $X=69780 $Y=47840
X2160 1 DigitalLDOLogic_VIA0 $T=70030 53520 0 0 $X=69780 $Y=53280
X2161 1 DigitalLDOLogic_VIA0 $T=70030 58960 0 0 $X=69780 $Y=58720
X2162 2 DigitalLDOLogic_VIA0 $T=71870 12720 0 0 $X=71620 $Y=12480
X2163 2 DigitalLDOLogic_VIA0 $T=71870 18160 0 0 $X=71620 $Y=17920
X2164 2 DigitalLDOLogic_VIA0 $T=71870 23600 0 0 $X=71620 $Y=23360
X2165 2 DigitalLDOLogic_VIA0 $T=71870 29040 0 0 $X=71620 $Y=28800
X2166 2 DigitalLDOLogic_VIA0 $T=71870 34480 0 0 $X=71620 $Y=34240
X2167 2 DigitalLDOLogic_VIA0 $T=71870 39920 0 0 $X=71620 $Y=39680
X2168 2 DigitalLDOLogic_VIA0 $T=71870 45360 0 0 $X=71620 $Y=45120
X2169 2 DigitalLDOLogic_VIA0 $T=71870 50800 0 0 $X=71620 $Y=50560
X2170 2 DigitalLDOLogic_VIA0 $T=71870 56240 0 0 $X=71620 $Y=56000
X2171 1 DigitalLDOLogic_VIA0 $T=72790 15440 0 0 $X=72540 $Y=15200
X2172 1 DigitalLDOLogic_VIA0 $T=72790 20880 0 0 $X=72540 $Y=20640
X2173 1 DigitalLDOLogic_VIA0 $T=72790 26320 0 0 $X=72540 $Y=26080
X2174 1 DigitalLDOLogic_VIA0 $T=72790 31760 0 0 $X=72540 $Y=31520
X2175 1 DigitalLDOLogic_VIA0 $T=72790 37200 0 0 $X=72540 $Y=36960
X2176 1 DigitalLDOLogic_VIA0 $T=72790 42640 0 0 $X=72540 $Y=42400
X2177 1 DigitalLDOLogic_VIA0 $T=72790 48080 0 0 $X=72540 $Y=47840
X2178 1 DigitalLDOLogic_VIA0 $T=72790 53520 0 0 $X=72540 $Y=53280
X2179 1 DigitalLDOLogic_VIA0 $T=72790 58960 0 0 $X=72540 $Y=58720
X2180 2 DigitalLDOLogic_VIA0 $T=74630 12720 0 0 $X=74380 $Y=12480
X2181 2 DigitalLDOLogic_VIA0 $T=74630 18160 0 0 $X=74380 $Y=17920
X2182 2 DigitalLDOLogic_VIA0 $T=74630 23600 0 0 $X=74380 $Y=23360
X2183 2 DigitalLDOLogic_VIA0 $T=74630 29040 0 0 $X=74380 $Y=28800
X2184 2 DigitalLDOLogic_VIA0 $T=74630 34480 0 0 $X=74380 $Y=34240
X2185 2 DigitalLDOLogic_VIA0 $T=74630 39920 0 0 $X=74380 $Y=39680
X2186 2 DigitalLDOLogic_VIA0 $T=74630 45360 0 0 $X=74380 $Y=45120
X2187 2 DigitalLDOLogic_VIA0 $T=74630 50800 0 0 $X=74380 $Y=50560
X2188 2 DigitalLDOLogic_VIA0 $T=74630 56240 0 0 $X=74380 $Y=56000
X2189 1 DigitalLDOLogic_VIA0 $T=75550 15440 0 0 $X=75300 $Y=15200
X2190 1 DigitalLDOLogic_VIA0 $T=75550 20880 0 0 $X=75300 $Y=20640
X2191 1 DigitalLDOLogic_VIA0 $T=75550 26320 0 0 $X=75300 $Y=26080
X2192 1 DigitalLDOLogic_VIA0 $T=75550 31760 0 0 $X=75300 $Y=31520
X2193 1 DigitalLDOLogic_VIA0 $T=75550 37200 0 0 $X=75300 $Y=36960
X2194 1 DigitalLDOLogic_VIA0 $T=75550 42640 0 0 $X=75300 $Y=42400
X2195 1 DigitalLDOLogic_VIA0 $T=75550 48080 0 0 $X=75300 $Y=47840
X2196 1 DigitalLDOLogic_VIA0 $T=75550 53520 0 0 $X=75300 $Y=53280
X2197 1 DigitalLDOLogic_VIA0 $T=75550 58960 0 0 $X=75300 $Y=58720
X2198 2 DigitalLDOLogic_VIA0 $T=77390 12720 0 0 $X=77140 $Y=12480
X2199 2 DigitalLDOLogic_VIA0 $T=77390 18160 0 0 $X=77140 $Y=17920
X2200 2 DigitalLDOLogic_VIA0 $T=77390 23600 0 0 $X=77140 $Y=23360
X2201 2 DigitalLDOLogic_VIA0 $T=77390 29040 0 0 $X=77140 $Y=28800
X2202 2 DigitalLDOLogic_VIA0 $T=77390 34480 0 0 $X=77140 $Y=34240
X2203 2 DigitalLDOLogic_VIA0 $T=77390 39920 0 0 $X=77140 $Y=39680
X2204 2 DigitalLDOLogic_VIA0 $T=77390 45360 0 0 $X=77140 $Y=45120
X2205 2 DigitalLDOLogic_VIA0 $T=77390 50800 0 0 $X=77140 $Y=50560
X2206 2 DigitalLDOLogic_VIA0 $T=77390 56240 0 0 $X=77140 $Y=56000
X2207 1 DigitalLDOLogic_VIA0 $T=78310 15440 0 0 $X=78060 $Y=15200
X2208 1 DigitalLDOLogic_VIA0 $T=78310 20880 0 0 $X=78060 $Y=20640
X2209 1 DigitalLDOLogic_VIA0 $T=78310 26320 0 0 $X=78060 $Y=26080
X2210 1 DigitalLDOLogic_VIA0 $T=78310 31760 0 0 $X=78060 $Y=31520
X2211 1 DigitalLDOLogic_VIA0 $T=78310 37200 0 0 $X=78060 $Y=36960
X2212 1 DigitalLDOLogic_VIA0 $T=78310 42640 0 0 $X=78060 $Y=42400
X2213 1 DigitalLDOLogic_VIA0 $T=78310 48080 0 0 $X=78060 $Y=47840
X2214 1 DigitalLDOLogic_VIA0 $T=78310 53520 0 0 $X=78060 $Y=53280
X2215 1 DigitalLDOLogic_VIA0 $T=78310 58960 0 0 $X=78060 $Y=58720
X2216 2 DigitalLDOLogic_VIA0 $T=80150 12720 0 0 $X=79900 $Y=12480
X2217 2 DigitalLDOLogic_VIA0 $T=80150 18160 0 0 $X=79900 $Y=17920
X2218 2 DigitalLDOLogic_VIA0 $T=80150 23600 0 0 $X=79900 $Y=23360
X2219 2 DigitalLDOLogic_VIA0 $T=80150 29040 0 0 $X=79900 $Y=28800
X2220 2 DigitalLDOLogic_VIA0 $T=80150 34480 0 0 $X=79900 $Y=34240
X2221 2 DigitalLDOLogic_VIA0 $T=80150 39920 0 0 $X=79900 $Y=39680
X2222 2 DigitalLDOLogic_VIA0 $T=80150 45360 0 0 $X=79900 $Y=45120
X2223 2 DigitalLDOLogic_VIA0 $T=80150 50800 0 0 $X=79900 $Y=50560
X2224 2 DigitalLDOLogic_VIA0 $T=80150 56240 0 0 $X=79900 $Y=56000
X2225 1 DigitalLDOLogic_VIA0 $T=81070 15440 0 0 $X=80820 $Y=15200
X2226 1 DigitalLDOLogic_VIA0 $T=81070 20880 0 0 $X=80820 $Y=20640
X2227 1 DigitalLDOLogic_VIA0 $T=81070 26320 0 0 $X=80820 $Y=26080
X2228 1 DigitalLDOLogic_VIA0 $T=81070 31760 0 0 $X=80820 $Y=31520
X2229 1 DigitalLDOLogic_VIA0 $T=81070 37200 0 0 $X=80820 $Y=36960
X2230 1 DigitalLDOLogic_VIA0 $T=81070 42640 0 0 $X=80820 $Y=42400
X2231 1 DigitalLDOLogic_VIA0 $T=81070 48080 0 0 $X=80820 $Y=47840
X2232 1 DigitalLDOLogic_VIA0 $T=81070 53520 0 0 $X=80820 $Y=53280
X2233 1 DigitalLDOLogic_VIA0 $T=81070 58960 0 0 $X=80820 $Y=58720
X2234 2 DigitalLDOLogic_VIA0 $T=82910 12720 0 0 $X=82660 $Y=12480
X2235 2 DigitalLDOLogic_VIA0 $T=82910 18160 0 0 $X=82660 $Y=17920
X2236 2 DigitalLDOLogic_VIA0 $T=82910 23600 0 0 $X=82660 $Y=23360
X2237 2 DigitalLDOLogic_VIA0 $T=82910 29040 0 0 $X=82660 $Y=28800
X2238 2 DigitalLDOLogic_VIA0 $T=82910 34480 0 0 $X=82660 $Y=34240
X2239 2 DigitalLDOLogic_VIA0 $T=82910 39920 0 0 $X=82660 $Y=39680
X2240 2 DigitalLDOLogic_VIA0 $T=82910 45360 0 0 $X=82660 $Y=45120
X2241 2 DigitalLDOLogic_VIA0 $T=82910 50800 0 0 $X=82660 $Y=50560
X2242 2 DigitalLDOLogic_VIA0 $T=82910 56240 0 0 $X=82660 $Y=56000
X2243 1 DigitalLDOLogic_VIA0 $T=83830 15440 0 0 $X=83580 $Y=15200
X2244 1 DigitalLDOLogic_VIA0 $T=83830 20880 0 0 $X=83580 $Y=20640
X2245 1 DigitalLDOLogic_VIA0 $T=83830 26320 0 0 $X=83580 $Y=26080
X2246 1 DigitalLDOLogic_VIA0 $T=83830 31760 0 0 $X=83580 $Y=31520
X2247 1 DigitalLDOLogic_VIA0 $T=83830 37200 0 0 $X=83580 $Y=36960
X2248 1 DigitalLDOLogic_VIA0 $T=83830 42640 0 0 $X=83580 $Y=42400
X2249 1 DigitalLDOLogic_VIA0 $T=83830 48080 0 0 $X=83580 $Y=47840
X2250 1 DigitalLDOLogic_VIA0 $T=83830 53520 0 0 $X=83580 $Y=53280
X2251 1 DigitalLDOLogic_VIA0 $T=83830 58960 0 0 $X=83580 $Y=58720
X2252 2 DigitalLDOLogic_VIA0 $T=85670 12720 0 0 $X=85420 $Y=12480
X2253 2 DigitalLDOLogic_VIA0 $T=85670 18160 0 0 $X=85420 $Y=17920
X2254 2 DigitalLDOLogic_VIA0 $T=85670 23600 0 0 $X=85420 $Y=23360
X2255 2 DigitalLDOLogic_VIA0 $T=85670 29040 0 0 $X=85420 $Y=28800
X2256 2 DigitalLDOLogic_VIA0 $T=85670 34480 0 0 $X=85420 $Y=34240
X2257 2 DigitalLDOLogic_VIA0 $T=85670 39920 0 0 $X=85420 $Y=39680
X2258 2 DigitalLDOLogic_VIA0 $T=85670 45360 0 0 $X=85420 $Y=45120
X2259 2 DigitalLDOLogic_VIA0 $T=85670 50800 0 0 $X=85420 $Y=50560
X2260 2 DigitalLDOLogic_VIA0 $T=85670 56240 0 0 $X=85420 $Y=56000
X2261 1 DigitalLDOLogic_VIA0 $T=86590 15440 0 0 $X=86340 $Y=15200
X2262 1 DigitalLDOLogic_VIA0 $T=86590 20880 0 0 $X=86340 $Y=20640
X2263 1 DigitalLDOLogic_VIA0 $T=86590 26320 0 0 $X=86340 $Y=26080
X2264 1 DigitalLDOLogic_VIA0 $T=86590 31760 0 0 $X=86340 $Y=31520
X2265 1 DigitalLDOLogic_VIA0 $T=86590 37200 0 0 $X=86340 $Y=36960
X2266 1 DigitalLDOLogic_VIA0 $T=86590 42640 0 0 $X=86340 $Y=42400
X2267 1 DigitalLDOLogic_VIA0 $T=86590 48080 0 0 $X=86340 $Y=47840
X2268 1 DigitalLDOLogic_VIA0 $T=86590 53520 0 0 $X=86340 $Y=53280
X2269 1 DigitalLDOLogic_VIA0 $T=86590 58960 0 0 $X=86340 $Y=58720
X2270 2 DigitalLDOLogic_VIA0 $T=88430 12720 0 0 $X=88180 $Y=12480
X2271 2 DigitalLDOLogic_VIA0 $T=88430 18160 0 0 $X=88180 $Y=17920
X2272 2 DigitalLDOLogic_VIA0 $T=88430 23600 0 0 $X=88180 $Y=23360
X2273 2 DigitalLDOLogic_VIA0 $T=88430 29040 0 0 $X=88180 $Y=28800
X2274 2 DigitalLDOLogic_VIA0 $T=88430 34480 0 0 $X=88180 $Y=34240
X2275 2 DigitalLDOLogic_VIA0 $T=88430 39920 0 0 $X=88180 $Y=39680
X2276 2 DigitalLDOLogic_VIA0 $T=88430 45360 0 0 $X=88180 $Y=45120
X2277 2 DigitalLDOLogic_VIA0 $T=88430 50800 0 0 $X=88180 $Y=50560
X2278 2 DigitalLDOLogic_VIA0 $T=88430 56240 0 0 $X=88180 $Y=56000
X2279 1 DigitalLDOLogic_VIA0 $T=89350 15440 0 0 $X=89100 $Y=15200
X2280 1 DigitalLDOLogic_VIA0 $T=89350 20880 0 0 $X=89100 $Y=20640
X2281 1 DigitalLDOLogic_VIA0 $T=89350 26320 0 0 $X=89100 $Y=26080
X2282 1 DigitalLDOLogic_VIA0 $T=89350 31760 0 0 $X=89100 $Y=31520
X2283 1 DigitalLDOLogic_VIA0 $T=89350 37200 0 0 $X=89100 $Y=36960
X2284 1 DigitalLDOLogic_VIA0 $T=89350 42640 0 0 $X=89100 $Y=42400
X2285 1 DigitalLDOLogic_VIA0 $T=89350 48080 0 0 $X=89100 $Y=47840
X2286 1 DigitalLDOLogic_VIA0 $T=89350 53520 0 0 $X=89100 $Y=53280
X2287 1 DigitalLDOLogic_VIA0 $T=89350 58960 0 0 $X=89100 $Y=58720
X2288 2 DigitalLDOLogic_VIA0 $T=91190 12720 0 0 $X=90940 $Y=12480
X2289 2 DigitalLDOLogic_VIA0 $T=91190 18160 0 0 $X=90940 $Y=17920
X2290 2 DigitalLDOLogic_VIA0 $T=91190 23600 0 0 $X=90940 $Y=23360
X2291 2 DigitalLDOLogic_VIA0 $T=91190 29040 0 0 $X=90940 $Y=28800
X2292 2 DigitalLDOLogic_VIA0 $T=91190 34480 0 0 $X=90940 $Y=34240
X2293 2 DigitalLDOLogic_VIA0 $T=91190 39920 0 0 $X=90940 $Y=39680
X2294 2 DigitalLDOLogic_VIA0 $T=91190 45360 0 0 $X=90940 $Y=45120
X2295 2 DigitalLDOLogic_VIA0 $T=91190 50800 0 0 $X=90940 $Y=50560
X2296 2 DigitalLDOLogic_VIA0 $T=91190 56240 0 0 $X=90940 $Y=56000
X2297 1 DigitalLDOLogic_VIA0 $T=92110 15440 0 0 $X=91860 $Y=15200
X2298 1 DigitalLDOLogic_VIA0 $T=92110 20880 0 0 $X=91860 $Y=20640
X2299 1 DigitalLDOLogic_VIA0 $T=92110 26320 0 0 $X=91860 $Y=26080
X2300 1 DigitalLDOLogic_VIA0 $T=92110 31760 0 0 $X=91860 $Y=31520
X2301 1 DigitalLDOLogic_VIA0 $T=92110 37200 0 0 $X=91860 $Y=36960
X2302 1 DigitalLDOLogic_VIA0 $T=92110 42640 0 0 $X=91860 $Y=42400
X2303 1 DigitalLDOLogic_VIA0 $T=92110 48080 0 0 $X=91860 $Y=47840
X2304 1 DigitalLDOLogic_VIA0 $T=92110 53520 0 0 $X=91860 $Y=53280
X2305 1 DigitalLDOLogic_VIA0 $T=92110 58960 0 0 $X=91860 $Y=58720
X2306 2 DigitalLDOLogic_VIA0 $T=93950 12720 0 0 $X=93700 $Y=12480
X2307 2 DigitalLDOLogic_VIA0 $T=93950 18160 0 0 $X=93700 $Y=17920
X2308 2 DigitalLDOLogic_VIA0 $T=93950 23600 0 0 $X=93700 $Y=23360
X2309 2 DigitalLDOLogic_VIA0 $T=93950 29040 0 0 $X=93700 $Y=28800
X2310 2 DigitalLDOLogic_VIA0 $T=93950 34480 0 0 $X=93700 $Y=34240
X2311 2 DigitalLDOLogic_VIA0 $T=93950 39920 0 0 $X=93700 $Y=39680
X2312 2 DigitalLDOLogic_VIA0 $T=93950 45360 0 0 $X=93700 $Y=45120
X2313 2 DigitalLDOLogic_VIA0 $T=93950 50800 0 0 $X=93700 $Y=50560
X2314 2 DigitalLDOLogic_VIA0 $T=93950 56240 0 0 $X=93700 $Y=56000
X2315 1 DigitalLDOLogic_VIA0 $T=94870 15440 0 0 $X=94620 $Y=15200
X2316 1 DigitalLDOLogic_VIA0 $T=94870 20880 0 0 $X=94620 $Y=20640
X2317 1 DigitalLDOLogic_VIA0 $T=94870 26320 0 0 $X=94620 $Y=26080
X2318 1 DigitalLDOLogic_VIA0 $T=94870 31760 0 0 $X=94620 $Y=31520
X2319 1 DigitalLDOLogic_VIA0 $T=94870 37200 0 0 $X=94620 $Y=36960
X2320 1 DigitalLDOLogic_VIA0 $T=94870 42640 0 0 $X=94620 $Y=42400
X2321 1 DigitalLDOLogic_VIA0 $T=94870 48080 0 0 $X=94620 $Y=47840
X2322 1 DigitalLDOLogic_VIA0 $T=94870 53520 0 0 $X=94620 $Y=53280
X2323 1 DigitalLDOLogic_VIA0 $T=94870 58960 0 0 $X=94620 $Y=58720
X2324 2 DigitalLDOLogic_VIA0 $T=96710 12720 0 0 $X=96460 $Y=12480
X2325 2 DigitalLDOLogic_VIA0 $T=96710 18160 0 0 $X=96460 $Y=17920
X2326 2 DigitalLDOLogic_VIA0 $T=96710 23600 0 0 $X=96460 $Y=23360
X2327 2 DigitalLDOLogic_VIA0 $T=96710 29040 0 0 $X=96460 $Y=28800
X2328 2 DigitalLDOLogic_VIA0 $T=96710 34480 0 0 $X=96460 $Y=34240
X2329 2 DigitalLDOLogic_VIA0 $T=96710 39920 0 0 $X=96460 $Y=39680
X2330 2 DigitalLDOLogic_VIA0 $T=96710 45360 0 0 $X=96460 $Y=45120
X2331 2 DigitalLDOLogic_VIA0 $T=96710 50800 0 0 $X=96460 $Y=50560
X2332 2 DigitalLDOLogic_VIA0 $T=96710 56240 0 0 $X=96460 $Y=56000
X2333 1 DigitalLDOLogic_VIA0 $T=97630 15440 0 0 $X=97380 $Y=15200
X2334 1 DigitalLDOLogic_VIA0 $T=97630 20880 0 0 $X=97380 $Y=20640
X2335 1 DigitalLDOLogic_VIA0 $T=97630 26320 0 0 $X=97380 $Y=26080
X2336 1 DigitalLDOLogic_VIA0 $T=97630 31760 0 0 $X=97380 $Y=31520
X2337 1 DigitalLDOLogic_VIA0 $T=97630 37200 0 0 $X=97380 $Y=36960
X2338 1 DigitalLDOLogic_VIA0 $T=97630 42640 0 0 $X=97380 $Y=42400
X2339 1 DigitalLDOLogic_VIA0 $T=97630 48080 0 0 $X=97380 $Y=47840
X2340 1 DigitalLDOLogic_VIA0 $T=97630 53520 0 0 $X=97380 $Y=53280
X2341 1 DigitalLDOLogic_VIA0 $T=97630 58960 0 0 $X=97380 $Y=58720
X2342 2 DigitalLDOLogic_VIA0 $T=99470 12720 0 0 $X=99220 $Y=12480
X2343 2 DigitalLDOLogic_VIA0 $T=99470 18160 0 0 $X=99220 $Y=17920
X2344 2 DigitalLDOLogic_VIA0 $T=99470 23600 0 0 $X=99220 $Y=23360
X2345 2 DigitalLDOLogic_VIA0 $T=99470 29040 0 0 $X=99220 $Y=28800
X2346 2 DigitalLDOLogic_VIA0 $T=99470 34480 0 0 $X=99220 $Y=34240
X2347 2 DigitalLDOLogic_VIA0 $T=99470 39920 0 0 $X=99220 $Y=39680
X2348 2 DigitalLDOLogic_VIA0 $T=99470 45360 0 0 $X=99220 $Y=45120
X2349 2 DigitalLDOLogic_VIA0 $T=99470 50800 0 0 $X=99220 $Y=50560
X2350 2 DigitalLDOLogic_VIA0 $T=99470 56240 0 0 $X=99220 $Y=56000
X2351 1 DigitalLDOLogic_VIA0 $T=100390 15440 0 0 $X=100140 $Y=15200
X2352 1 DigitalLDOLogic_VIA0 $T=100390 20880 0 0 $X=100140 $Y=20640
X2353 1 DigitalLDOLogic_VIA0 $T=100390 26320 0 0 $X=100140 $Y=26080
X2354 1 DigitalLDOLogic_VIA0 $T=100390 31760 0 0 $X=100140 $Y=31520
X2355 1 DigitalLDOLogic_VIA0 $T=100390 37200 0 0 $X=100140 $Y=36960
X2356 1 DigitalLDOLogic_VIA0 $T=100390 42640 0 0 $X=100140 $Y=42400
X2357 1 DigitalLDOLogic_VIA0 $T=100390 48080 0 0 $X=100140 $Y=47840
X2358 1 DigitalLDOLogic_VIA0 $T=100390 53520 0 0 $X=100140 $Y=53280
X2359 1 DigitalLDOLogic_VIA0 $T=100390 58960 0 0 $X=100140 $Y=58720
X2360 2 DigitalLDOLogic_VIA0 $T=102230 12720 0 0 $X=101980 $Y=12480
X2361 2 DigitalLDOLogic_VIA0 $T=102230 18160 0 0 $X=101980 $Y=17920
X2362 2 DigitalLDOLogic_VIA0 $T=102230 23600 0 0 $X=101980 $Y=23360
X2363 2 DigitalLDOLogic_VIA0 $T=102230 29040 0 0 $X=101980 $Y=28800
X2364 2 DigitalLDOLogic_VIA0 $T=102230 34480 0 0 $X=101980 $Y=34240
X2365 2 DigitalLDOLogic_VIA0 $T=102230 39920 0 0 $X=101980 $Y=39680
X2366 2 DigitalLDOLogic_VIA0 $T=102230 45360 0 0 $X=101980 $Y=45120
X2367 2 DigitalLDOLogic_VIA0 $T=102230 50800 0 0 $X=101980 $Y=50560
X2368 2 DigitalLDOLogic_VIA0 $T=102230 56240 0 0 $X=101980 $Y=56000
X2369 1 DigitalLDOLogic_VIA0 $T=103150 15440 0 0 $X=102900 $Y=15200
X2370 1 DigitalLDOLogic_VIA0 $T=103150 20880 0 0 $X=102900 $Y=20640
X2371 1 DigitalLDOLogic_VIA0 $T=103150 26320 0 0 $X=102900 $Y=26080
X2372 1 DigitalLDOLogic_VIA0 $T=103150 31760 0 0 $X=102900 $Y=31520
X2373 1 DigitalLDOLogic_VIA0 $T=103150 37200 0 0 $X=102900 $Y=36960
X2374 1 DigitalLDOLogic_VIA0 $T=103150 42640 0 0 $X=102900 $Y=42400
X2375 1 DigitalLDOLogic_VIA0 $T=103150 48080 0 0 $X=102900 $Y=47840
X2376 1 DigitalLDOLogic_VIA0 $T=103150 53520 0 0 $X=102900 $Y=53280
X2377 1 DigitalLDOLogic_VIA0 $T=103150 58960 0 0 $X=102900 $Y=58720
X2378 2 DigitalLDOLogic_VIA0 $T=104990 12720 0 0 $X=104740 $Y=12480
X2379 2 DigitalLDOLogic_VIA0 $T=104990 18160 0 0 $X=104740 $Y=17920
X2380 2 DigitalLDOLogic_VIA0 $T=104990 23600 0 0 $X=104740 $Y=23360
X2381 2 DigitalLDOLogic_VIA0 $T=104990 29040 0 0 $X=104740 $Y=28800
X2382 2 DigitalLDOLogic_VIA0 $T=104990 34480 0 0 $X=104740 $Y=34240
X2383 2 DigitalLDOLogic_VIA0 $T=104990 39920 0 0 $X=104740 $Y=39680
X2384 2 DigitalLDOLogic_VIA0 $T=104990 45360 0 0 $X=104740 $Y=45120
X2385 2 DigitalLDOLogic_VIA0 $T=104990 50800 0 0 $X=104740 $Y=50560
X2386 2 DigitalLDOLogic_VIA0 $T=104990 56240 0 0 $X=104740 $Y=56000
X2387 1 DigitalLDOLogic_VIA0 $T=105910 15440 0 0 $X=105660 $Y=15200
X2388 1 DigitalLDOLogic_VIA0 $T=105910 20880 0 0 $X=105660 $Y=20640
X2389 1 DigitalLDOLogic_VIA0 $T=105910 26320 0 0 $X=105660 $Y=26080
X2390 1 DigitalLDOLogic_VIA0 $T=105910 31760 0 0 $X=105660 $Y=31520
X2391 1 DigitalLDOLogic_VIA0 $T=105910 37200 0 0 $X=105660 $Y=36960
X2392 1 DigitalLDOLogic_VIA0 $T=105910 42640 0 0 $X=105660 $Y=42400
X2393 1 DigitalLDOLogic_VIA0 $T=105910 48080 0 0 $X=105660 $Y=47840
X2394 1 DigitalLDOLogic_VIA0 $T=105910 53520 0 0 $X=105660 $Y=53280
X2395 1 DigitalLDOLogic_VIA0 $T=105910 58960 0 0 $X=105660 $Y=58720
X2396 2 DigitalLDOLogic_VIA0 $T=107750 12720 0 0 $X=107500 $Y=12480
X2397 2 DigitalLDOLogic_VIA0 $T=107750 18160 0 0 $X=107500 $Y=17920
X2398 2 DigitalLDOLogic_VIA0 $T=107750 23600 0 0 $X=107500 $Y=23360
X2399 2 DigitalLDOLogic_VIA0 $T=107750 29040 0 0 $X=107500 $Y=28800
X2400 2 DigitalLDOLogic_VIA0 $T=107750 34480 0 0 $X=107500 $Y=34240
X2401 2 DigitalLDOLogic_VIA0 $T=107750 39920 0 0 $X=107500 $Y=39680
X2402 2 DigitalLDOLogic_VIA0 $T=107750 45360 0 0 $X=107500 $Y=45120
X2403 2 DigitalLDOLogic_VIA0 $T=107750 50800 0 0 $X=107500 $Y=50560
X2404 2 DigitalLDOLogic_VIA0 $T=107750 56240 0 0 $X=107500 $Y=56000
X2405 1 DigitalLDOLogic_VIA0 $T=108670 15440 0 0 $X=108420 $Y=15200
X2406 1 DigitalLDOLogic_VIA0 $T=108670 20880 0 0 $X=108420 $Y=20640
X2407 1 DigitalLDOLogic_VIA0 $T=108670 26320 0 0 $X=108420 $Y=26080
X2408 1 DigitalLDOLogic_VIA0 $T=108670 31760 0 0 $X=108420 $Y=31520
X2409 1 DigitalLDOLogic_VIA0 $T=108670 37200 0 0 $X=108420 $Y=36960
X2410 1 DigitalLDOLogic_VIA0 $T=108670 42640 0 0 $X=108420 $Y=42400
X2411 1 DigitalLDOLogic_VIA0 $T=108670 48080 0 0 $X=108420 $Y=47840
X2412 1 DigitalLDOLogic_VIA0 $T=108670 53520 0 0 $X=108420 $Y=53280
X2413 1 DigitalLDOLogic_VIA0 $T=108670 58960 0 0 $X=108420 $Y=58720
X2414 2 DigitalLDOLogic_VIA0 $T=110510 12720 0 0 $X=110260 $Y=12480
X2415 2 DigitalLDOLogic_VIA0 $T=110510 18160 0 0 $X=110260 $Y=17920
X2416 2 DigitalLDOLogic_VIA0 $T=110510 23600 0 0 $X=110260 $Y=23360
X2417 2 DigitalLDOLogic_VIA0 $T=110510 29040 0 0 $X=110260 $Y=28800
X2418 2 DigitalLDOLogic_VIA0 $T=110510 34480 0 0 $X=110260 $Y=34240
X2419 2 DigitalLDOLogic_VIA0 $T=110510 39920 0 0 $X=110260 $Y=39680
X2420 2 DigitalLDOLogic_VIA0 $T=110510 45360 0 0 $X=110260 $Y=45120
X2421 2 DigitalLDOLogic_VIA0 $T=110510 50800 0 0 $X=110260 $Y=50560
X2422 2 DigitalLDOLogic_VIA0 $T=110510 56240 0 0 $X=110260 $Y=56000
X2423 1 DigitalLDOLogic_VIA0 $T=111430 15440 0 0 $X=111180 $Y=15200
X2424 1 DigitalLDOLogic_VIA0 $T=111430 20880 0 0 $X=111180 $Y=20640
X2425 1 DigitalLDOLogic_VIA0 $T=111430 26320 0 0 $X=111180 $Y=26080
X2426 1 DigitalLDOLogic_VIA0 $T=111430 31760 0 0 $X=111180 $Y=31520
X2427 1 DigitalLDOLogic_VIA0 $T=111430 37200 0 0 $X=111180 $Y=36960
X2428 1 DigitalLDOLogic_VIA0 $T=111430 42640 0 0 $X=111180 $Y=42400
X2429 1 DigitalLDOLogic_VIA0 $T=111430 48080 0 0 $X=111180 $Y=47840
X2430 1 DigitalLDOLogic_VIA0 $T=111430 53520 0 0 $X=111180 $Y=53280
X2431 1 DigitalLDOLogic_VIA0 $T=111430 58960 0 0 $X=111180 $Y=58720
X2432 2 DigitalLDOLogic_VIA0 $T=113270 12720 0 0 $X=113020 $Y=12480
X2433 2 DigitalLDOLogic_VIA0 $T=113270 18160 0 0 $X=113020 $Y=17920
X2434 2 DigitalLDOLogic_VIA0 $T=113270 23600 0 0 $X=113020 $Y=23360
X2435 2 DigitalLDOLogic_VIA0 $T=113270 29040 0 0 $X=113020 $Y=28800
X2436 2 DigitalLDOLogic_VIA0 $T=113270 34480 0 0 $X=113020 $Y=34240
X2437 2 DigitalLDOLogic_VIA0 $T=113270 39920 0 0 $X=113020 $Y=39680
X2438 2 DigitalLDOLogic_VIA0 $T=113270 45360 0 0 $X=113020 $Y=45120
X2439 2 DigitalLDOLogic_VIA0 $T=113270 50800 0 0 $X=113020 $Y=50560
X2440 2 DigitalLDOLogic_VIA0 $T=113270 56240 0 0 $X=113020 $Y=56000
X2441 1 DigitalLDOLogic_VIA0 $T=114190 15440 0 0 $X=113940 $Y=15200
X2442 1 DigitalLDOLogic_VIA0 $T=114190 20880 0 0 $X=113940 $Y=20640
X2443 1 DigitalLDOLogic_VIA0 $T=114190 26320 0 0 $X=113940 $Y=26080
X2444 1 DigitalLDOLogic_VIA0 $T=114190 31760 0 0 $X=113940 $Y=31520
X2445 1 DigitalLDOLogic_VIA0 $T=114190 37200 0 0 $X=113940 $Y=36960
X2446 1 DigitalLDOLogic_VIA0 $T=114190 42640 0 0 $X=113940 $Y=42400
X2447 1 DigitalLDOLogic_VIA0 $T=114190 48080 0 0 $X=113940 $Y=47840
X2448 1 DigitalLDOLogic_VIA0 $T=114190 53520 0 0 $X=113940 $Y=53280
X2449 1 DigitalLDOLogic_VIA0 $T=114190 58960 0 0 $X=113940 $Y=58720
X2450 2 DigitalLDOLogic_VIA0 $T=116030 12720 0 0 $X=115780 $Y=12480
X2451 2 DigitalLDOLogic_VIA0 $T=116030 18160 0 0 $X=115780 $Y=17920
X2452 2 DigitalLDOLogic_VIA0 $T=116030 23600 0 0 $X=115780 $Y=23360
X2453 2 DigitalLDOLogic_VIA0 $T=116030 29040 0 0 $X=115780 $Y=28800
X2454 2 DigitalLDOLogic_VIA0 $T=116030 34480 0 0 $X=115780 $Y=34240
X2455 2 DigitalLDOLogic_VIA0 $T=116030 39920 0 0 $X=115780 $Y=39680
X2456 2 DigitalLDOLogic_VIA0 $T=116030 45360 0 0 $X=115780 $Y=45120
X2457 2 DigitalLDOLogic_VIA0 $T=116030 50800 0 0 $X=115780 $Y=50560
X2458 2 DigitalLDOLogic_VIA0 $T=116030 56240 0 0 $X=115780 $Y=56000
X2459 1 DigitalLDOLogic_VIA0 $T=116950 15440 0 0 $X=116700 $Y=15200
X2460 1 DigitalLDOLogic_VIA0 $T=116950 20880 0 0 $X=116700 $Y=20640
X2461 1 DigitalLDOLogic_VIA0 $T=116950 26320 0 0 $X=116700 $Y=26080
X2462 1 DigitalLDOLogic_VIA0 $T=116950 31760 0 0 $X=116700 $Y=31520
X2463 1 DigitalLDOLogic_VIA0 $T=116950 37200 0 0 $X=116700 $Y=36960
X2464 1 DigitalLDOLogic_VIA0 $T=116950 42640 0 0 $X=116700 $Y=42400
X2465 1 DigitalLDOLogic_VIA0 $T=116950 48080 0 0 $X=116700 $Y=47840
X2466 1 DigitalLDOLogic_VIA0 $T=116950 53520 0 0 $X=116700 $Y=53280
X2467 1 DigitalLDOLogic_VIA0 $T=116950 58960 0 0 $X=116700 $Y=58720
X2468 2 DigitalLDOLogic_VIA0 $T=118790 12720 0 0 $X=118540 $Y=12480
X2469 2 DigitalLDOLogic_VIA0 $T=118790 18160 0 0 $X=118540 $Y=17920
X2470 2 DigitalLDOLogic_VIA0 $T=118790 23600 0 0 $X=118540 $Y=23360
X2471 2 DigitalLDOLogic_VIA0 $T=118790 29040 0 0 $X=118540 $Y=28800
X2472 2 DigitalLDOLogic_VIA0 $T=118790 34480 0 0 $X=118540 $Y=34240
X2473 2 DigitalLDOLogic_VIA0 $T=118790 39920 0 0 $X=118540 $Y=39680
X2474 2 DigitalLDOLogic_VIA0 $T=118790 45360 0 0 $X=118540 $Y=45120
X2475 2 DigitalLDOLogic_VIA0 $T=118790 50800 0 0 $X=118540 $Y=50560
X2476 2 DigitalLDOLogic_VIA0 $T=118790 56240 0 0 $X=118540 $Y=56000
X2477 1 DigitalLDOLogic_VIA0 $T=119710 15440 0 0 $X=119460 $Y=15200
X2478 1 DigitalLDOLogic_VIA0 $T=119710 20880 0 0 $X=119460 $Y=20640
X2479 1 DigitalLDOLogic_VIA0 $T=119710 26320 0 0 $X=119460 $Y=26080
X2480 1 DigitalLDOLogic_VIA0 $T=119710 31760 0 0 $X=119460 $Y=31520
X2481 1 DigitalLDOLogic_VIA0 $T=119710 37200 0 0 $X=119460 $Y=36960
X2482 1 DigitalLDOLogic_VIA0 $T=119710 42640 0 0 $X=119460 $Y=42400
X2483 1 DigitalLDOLogic_VIA0 $T=119710 48080 0 0 $X=119460 $Y=47840
X2484 1 DigitalLDOLogic_VIA0 $T=119710 53520 0 0 $X=119460 $Y=53280
X2485 1 DigitalLDOLogic_VIA0 $T=119710 58960 0 0 $X=119460 $Y=58720
X2486 2 DigitalLDOLogic_VIA0 $T=121550 12720 0 0 $X=121300 $Y=12480
X2487 2 DigitalLDOLogic_VIA0 $T=121550 18160 0 0 $X=121300 $Y=17920
X2488 2 DigitalLDOLogic_VIA0 $T=121550 23600 0 0 $X=121300 $Y=23360
X2489 2 DigitalLDOLogic_VIA0 $T=121550 29040 0 0 $X=121300 $Y=28800
X2490 2 DigitalLDOLogic_VIA0 $T=121550 34480 0 0 $X=121300 $Y=34240
X2491 2 DigitalLDOLogic_VIA0 $T=121550 39920 0 0 $X=121300 $Y=39680
X2492 2 DigitalLDOLogic_VIA0 $T=121550 45360 0 0 $X=121300 $Y=45120
X2493 2 DigitalLDOLogic_VIA0 $T=121550 50800 0 0 $X=121300 $Y=50560
X2494 2 DigitalLDOLogic_VIA0 $T=121550 56240 0 0 $X=121300 $Y=56000
X2495 1 DigitalLDOLogic_VIA0 $T=122470 15440 0 0 $X=122220 $Y=15200
X2496 1 DigitalLDOLogic_VIA0 $T=122470 20880 0 0 $X=122220 $Y=20640
X2497 1 DigitalLDOLogic_VIA0 $T=122470 26320 0 0 $X=122220 $Y=26080
X2498 1 DigitalLDOLogic_VIA0 $T=122470 31760 0 0 $X=122220 $Y=31520
X2499 1 DigitalLDOLogic_VIA0 $T=122470 37200 0 0 $X=122220 $Y=36960
X2500 1 DigitalLDOLogic_VIA0 $T=122470 42640 0 0 $X=122220 $Y=42400
X2501 1 DigitalLDOLogic_VIA0 $T=122470 48080 0 0 $X=122220 $Y=47840
X2502 1 DigitalLDOLogic_VIA0 $T=122470 53520 0 0 $X=122220 $Y=53280
X2503 1 DigitalLDOLogic_VIA0 $T=122470 58960 0 0 $X=122220 $Y=58720
X2504 2 DigitalLDOLogic_VIA0 $T=124310 12720 0 0 $X=124060 $Y=12480
X2505 2 DigitalLDOLogic_VIA0 $T=124310 18160 0 0 $X=124060 $Y=17920
X2506 2 DigitalLDOLogic_VIA0 $T=124310 23600 0 0 $X=124060 $Y=23360
X2507 2 DigitalLDOLogic_VIA0 $T=124310 29040 0 0 $X=124060 $Y=28800
X2508 2 DigitalLDOLogic_VIA0 $T=124310 34480 0 0 $X=124060 $Y=34240
X2509 2 DigitalLDOLogic_VIA0 $T=124310 39920 0 0 $X=124060 $Y=39680
X2510 2 DigitalLDOLogic_VIA0 $T=124310 45360 0 0 $X=124060 $Y=45120
X2511 2 DigitalLDOLogic_VIA0 $T=124310 50800 0 0 $X=124060 $Y=50560
X2512 2 DigitalLDOLogic_VIA0 $T=124310 56240 0 0 $X=124060 $Y=56000
X2513 1 DigitalLDOLogic_VIA0 $T=125230 15440 0 0 $X=124980 $Y=15200
X2514 1 DigitalLDOLogic_VIA0 $T=125230 20880 0 0 $X=124980 $Y=20640
X2515 1 DigitalLDOLogic_VIA0 $T=125230 26320 0 0 $X=124980 $Y=26080
X2516 1 DigitalLDOLogic_VIA0 $T=125230 31760 0 0 $X=124980 $Y=31520
X2517 1 DigitalLDOLogic_VIA0 $T=125230 37200 0 0 $X=124980 $Y=36960
X2518 1 DigitalLDOLogic_VIA0 $T=125230 42640 0 0 $X=124980 $Y=42400
X2519 1 DigitalLDOLogic_VIA0 $T=125230 48080 0 0 $X=124980 $Y=47840
X2520 1 DigitalLDOLogic_VIA0 $T=125230 53520 0 0 $X=124980 $Y=53280
X2521 1 DigitalLDOLogic_VIA0 $T=125230 58960 0 0 $X=124980 $Y=58720
X2522 2 DigitalLDOLogic_VIA0 $T=127070 12720 0 0 $X=126820 $Y=12480
X2523 2 DigitalLDOLogic_VIA0 $T=127070 18160 0 0 $X=126820 $Y=17920
X2524 2 DigitalLDOLogic_VIA0 $T=127070 23600 0 0 $X=126820 $Y=23360
X2525 2 DigitalLDOLogic_VIA0 $T=127070 29040 0 0 $X=126820 $Y=28800
X2526 2 DigitalLDOLogic_VIA0 $T=127070 34480 0 0 $X=126820 $Y=34240
X2527 2 DigitalLDOLogic_VIA0 $T=127070 39920 0 0 $X=126820 $Y=39680
X2528 2 DigitalLDOLogic_VIA0 $T=127070 45360 0 0 $X=126820 $Y=45120
X2529 2 DigitalLDOLogic_VIA0 $T=127070 50800 0 0 $X=126820 $Y=50560
X2530 2 DigitalLDOLogic_VIA0 $T=127070 56240 0 0 $X=126820 $Y=56000
X2531 1 DigitalLDOLogic_VIA0 $T=127990 15440 0 0 $X=127740 $Y=15200
X2532 1 DigitalLDOLogic_VIA0 $T=127990 20880 0 0 $X=127740 $Y=20640
X2533 1 DigitalLDOLogic_VIA0 $T=127990 26320 0 0 $X=127740 $Y=26080
X2534 1 DigitalLDOLogic_VIA0 $T=127990 31760 0 0 $X=127740 $Y=31520
X2535 1 DigitalLDOLogic_VIA0 $T=127990 37200 0 0 $X=127740 $Y=36960
X2536 1 DigitalLDOLogic_VIA0 $T=127990 42640 0 0 $X=127740 $Y=42400
X2537 1 DigitalLDOLogic_VIA0 $T=127990 48080 0 0 $X=127740 $Y=47840
X2538 1 DigitalLDOLogic_VIA0 $T=127990 53520 0 0 $X=127740 $Y=53280
X2539 1 DigitalLDOLogic_VIA0 $T=127990 58960 0 0 $X=127740 $Y=58720
X2540 2 DigitalLDOLogic_VIA0 $T=129830 12720 0 0 $X=129580 $Y=12480
X2541 2 DigitalLDOLogic_VIA0 $T=129830 18160 0 0 $X=129580 $Y=17920
X2542 2 DigitalLDOLogic_VIA0 $T=129830 23600 0 0 $X=129580 $Y=23360
X2543 2 DigitalLDOLogic_VIA0 $T=129830 29040 0 0 $X=129580 $Y=28800
X2544 2 DigitalLDOLogic_VIA0 $T=129830 34480 0 0 $X=129580 $Y=34240
X2545 2 DigitalLDOLogic_VIA0 $T=129830 39920 0 0 $X=129580 $Y=39680
X2546 2 DigitalLDOLogic_VIA0 $T=129830 45360 0 0 $X=129580 $Y=45120
X2547 2 DigitalLDOLogic_VIA0 $T=129830 50800 0 0 $X=129580 $Y=50560
X2548 2 DigitalLDOLogic_VIA0 $T=129830 56240 0 0 $X=129580 $Y=56000
X2549 1 DigitalLDOLogic_VIA0 $T=130750 15440 0 0 $X=130500 $Y=15200
X2550 1 DigitalLDOLogic_VIA0 $T=130750 20880 0 0 $X=130500 $Y=20640
X2551 1 DigitalLDOLogic_VIA0 $T=130750 26320 0 0 $X=130500 $Y=26080
X2552 1 DigitalLDOLogic_VIA0 $T=130750 31760 0 0 $X=130500 $Y=31520
X2553 1 DigitalLDOLogic_VIA0 $T=130750 37200 0 0 $X=130500 $Y=36960
X2554 1 DigitalLDOLogic_VIA0 $T=130750 42640 0 0 $X=130500 $Y=42400
X2555 1 DigitalLDOLogic_VIA0 $T=130750 48080 0 0 $X=130500 $Y=47840
X2556 1 DigitalLDOLogic_VIA0 $T=130750 53520 0 0 $X=130500 $Y=53280
X2557 1 DigitalLDOLogic_VIA0 $T=130750 58960 0 0 $X=130500 $Y=58720
X2558 2 DigitalLDOLogic_VIA0 $T=132590 12720 0 0 $X=132340 $Y=12480
X2559 2 DigitalLDOLogic_VIA0 $T=132590 18160 0 0 $X=132340 $Y=17920
X2560 2 DigitalLDOLogic_VIA0 $T=132590 23600 0 0 $X=132340 $Y=23360
X2561 2 DigitalLDOLogic_VIA0 $T=132590 29040 0 0 $X=132340 $Y=28800
X2562 2 DigitalLDOLogic_VIA0 $T=132590 34480 0 0 $X=132340 $Y=34240
X2563 2 DigitalLDOLogic_VIA0 $T=132590 39920 0 0 $X=132340 $Y=39680
X2564 2 DigitalLDOLogic_VIA0 $T=132590 45360 0 0 $X=132340 $Y=45120
X2565 2 DigitalLDOLogic_VIA0 $T=132590 50800 0 0 $X=132340 $Y=50560
X2566 2 DigitalLDOLogic_VIA0 $T=132590 56240 0 0 $X=132340 $Y=56000
X2567 1 DigitalLDOLogic_VIA0 $T=133510 15440 0 0 $X=133260 $Y=15200
X2568 1 DigitalLDOLogic_VIA0 $T=133510 20880 0 0 $X=133260 $Y=20640
X2569 1 DigitalLDOLogic_VIA0 $T=133510 26320 0 0 $X=133260 $Y=26080
X2570 1 DigitalLDOLogic_VIA0 $T=133510 31760 0 0 $X=133260 $Y=31520
X2571 1 DigitalLDOLogic_VIA0 $T=133510 37200 0 0 $X=133260 $Y=36960
X2572 1 DigitalLDOLogic_VIA0 $T=133510 42640 0 0 $X=133260 $Y=42400
X2573 1 DigitalLDOLogic_VIA0 $T=133510 48080 0 0 $X=133260 $Y=47840
X2574 1 DigitalLDOLogic_VIA0 $T=133510 53520 0 0 $X=133260 $Y=53280
X2575 1 DigitalLDOLogic_VIA0 $T=133510 58960 0 0 $X=133260 $Y=58720
X2576 2 DigitalLDOLogic_VIA0 $T=135350 12720 0 0 $X=135100 $Y=12480
X2577 2 DigitalLDOLogic_VIA0 $T=135350 18160 0 0 $X=135100 $Y=17920
X2578 2 DigitalLDOLogic_VIA0 $T=135350 23600 0 0 $X=135100 $Y=23360
X2579 2 DigitalLDOLogic_VIA0 $T=135350 29040 0 0 $X=135100 $Y=28800
X2580 2 DigitalLDOLogic_VIA0 $T=135350 34480 0 0 $X=135100 $Y=34240
X2581 2 DigitalLDOLogic_VIA0 $T=135350 39920 0 0 $X=135100 $Y=39680
X2582 2 DigitalLDOLogic_VIA0 $T=135350 45360 0 0 $X=135100 $Y=45120
X2583 2 DigitalLDOLogic_VIA0 $T=135350 50800 0 0 $X=135100 $Y=50560
X2584 2 DigitalLDOLogic_VIA0 $T=135350 56240 0 0 $X=135100 $Y=56000
X2585 1 DigitalLDOLogic_VIA0 $T=136270 15440 0 0 $X=136020 $Y=15200
X2586 1 DigitalLDOLogic_VIA0 $T=136270 20880 0 0 $X=136020 $Y=20640
X2587 1 DigitalLDOLogic_VIA0 $T=136270 26320 0 0 $X=136020 $Y=26080
X2588 1 DigitalLDOLogic_VIA0 $T=136270 31760 0 0 $X=136020 $Y=31520
X2589 1 DigitalLDOLogic_VIA0 $T=136270 37200 0 0 $X=136020 $Y=36960
X2590 1 DigitalLDOLogic_VIA0 $T=136270 42640 0 0 $X=136020 $Y=42400
X2591 1 DigitalLDOLogic_VIA0 $T=136270 48080 0 0 $X=136020 $Y=47840
X2592 1 DigitalLDOLogic_VIA0 $T=136270 53520 0 0 $X=136020 $Y=53280
X2593 1 DigitalLDOLogic_VIA0 $T=136270 58960 0 0 $X=136020 $Y=58720
X2594 2 DigitalLDOLogic_VIA0 $T=138110 12720 0 0 $X=137860 $Y=12480
X2595 2 DigitalLDOLogic_VIA0 $T=138110 18160 0 0 $X=137860 $Y=17920
X2596 2 DigitalLDOLogic_VIA0 $T=138110 23600 0 0 $X=137860 $Y=23360
X2597 2 DigitalLDOLogic_VIA0 $T=138110 29040 0 0 $X=137860 $Y=28800
X2598 2 DigitalLDOLogic_VIA0 $T=138110 34480 0 0 $X=137860 $Y=34240
X2599 2 DigitalLDOLogic_VIA0 $T=138110 39920 0 0 $X=137860 $Y=39680
X2600 2 DigitalLDOLogic_VIA0 $T=138110 45360 0 0 $X=137860 $Y=45120
X2601 2 DigitalLDOLogic_VIA0 $T=138110 50800 0 0 $X=137860 $Y=50560
X2602 2 DigitalLDOLogic_VIA0 $T=138110 56240 0 0 $X=137860 $Y=56000
X2603 1 DigitalLDOLogic_VIA0 $T=139030 15440 0 0 $X=138780 $Y=15200
X2604 1 DigitalLDOLogic_VIA0 $T=139030 20880 0 0 $X=138780 $Y=20640
X2605 1 DigitalLDOLogic_VIA0 $T=139030 26320 0 0 $X=138780 $Y=26080
X2606 1 DigitalLDOLogic_VIA0 $T=139030 31760 0 0 $X=138780 $Y=31520
X2607 1 DigitalLDOLogic_VIA0 $T=139030 37200 0 0 $X=138780 $Y=36960
X2608 1 DigitalLDOLogic_VIA0 $T=139030 42640 0 0 $X=138780 $Y=42400
X2609 1 DigitalLDOLogic_VIA0 $T=139030 48080 0 0 $X=138780 $Y=47840
X2610 1 DigitalLDOLogic_VIA0 $T=139030 53520 0 0 $X=138780 $Y=53280
X2611 1 DigitalLDOLogic_VIA0 $T=139030 58960 0 0 $X=138780 $Y=58720
X2612 2 DigitalLDOLogic_VIA0 $T=140870 12720 0 0 $X=140620 $Y=12480
X2613 2 DigitalLDOLogic_VIA0 $T=140870 18160 0 0 $X=140620 $Y=17920
X2614 2 DigitalLDOLogic_VIA0 $T=140870 23600 0 0 $X=140620 $Y=23360
X2615 2 DigitalLDOLogic_VIA0 $T=140870 29040 0 0 $X=140620 $Y=28800
X2616 2 DigitalLDOLogic_VIA0 $T=140870 34480 0 0 $X=140620 $Y=34240
X2617 2 DigitalLDOLogic_VIA0 $T=140870 39920 0 0 $X=140620 $Y=39680
X2618 2 DigitalLDOLogic_VIA0 $T=140870 45360 0 0 $X=140620 $Y=45120
X2619 2 DigitalLDOLogic_VIA0 $T=140870 50800 0 0 $X=140620 $Y=50560
X2620 2 DigitalLDOLogic_VIA0 $T=140870 56240 0 0 $X=140620 $Y=56000
X2621 1 DigitalLDOLogic_VIA0 $T=141790 15440 0 0 $X=141540 $Y=15200
X2622 1 DigitalLDOLogic_VIA0 $T=141790 20880 0 0 $X=141540 $Y=20640
X2623 1 DigitalLDOLogic_VIA0 $T=141790 26320 0 0 $X=141540 $Y=26080
X2624 1 DigitalLDOLogic_VIA0 $T=141790 31760 0 0 $X=141540 $Y=31520
X2625 1 DigitalLDOLogic_VIA0 $T=141790 37200 0 0 $X=141540 $Y=36960
X2626 1 DigitalLDOLogic_VIA0 $T=141790 42640 0 0 $X=141540 $Y=42400
X2627 1 DigitalLDOLogic_VIA0 $T=141790 48080 0 0 $X=141540 $Y=47840
X2628 1 DigitalLDOLogic_VIA0 $T=141790 53520 0 0 $X=141540 $Y=53280
X2629 1 DigitalLDOLogic_VIA0 $T=141790 58960 0 0 $X=141540 $Y=58720
X2630 2 DigitalLDOLogic_VIA0 $T=143630 12720 0 0 $X=143380 $Y=12480
X2631 2 DigitalLDOLogic_VIA0 $T=143630 18160 0 0 $X=143380 $Y=17920
X2632 2 DigitalLDOLogic_VIA0 $T=143630 23600 0 0 $X=143380 $Y=23360
X2633 2 DigitalLDOLogic_VIA0 $T=143630 29040 0 0 $X=143380 $Y=28800
X2634 2 DigitalLDOLogic_VIA0 $T=143630 34480 0 0 $X=143380 $Y=34240
X2635 2 DigitalLDOLogic_VIA0 $T=143630 39920 0 0 $X=143380 $Y=39680
X2636 2 DigitalLDOLogic_VIA0 $T=143630 45360 0 0 $X=143380 $Y=45120
X2637 2 DigitalLDOLogic_VIA0 $T=143630 50800 0 0 $X=143380 $Y=50560
X2638 2 DigitalLDOLogic_VIA0 $T=143630 56240 0 0 $X=143380 $Y=56000
X2639 1 DigitalLDOLogic_VIA0 $T=144550 15440 0 0 $X=144300 $Y=15200
X2640 1 DigitalLDOLogic_VIA0 $T=144550 20880 0 0 $X=144300 $Y=20640
X2641 1 DigitalLDOLogic_VIA0 $T=144550 26320 0 0 $X=144300 $Y=26080
X2642 1 DigitalLDOLogic_VIA0 $T=144550 31760 0 0 $X=144300 $Y=31520
X2643 1 DigitalLDOLogic_VIA0 $T=144550 37200 0 0 $X=144300 $Y=36960
X2644 1 DigitalLDOLogic_VIA0 $T=144550 42640 0 0 $X=144300 $Y=42400
X2645 1 DigitalLDOLogic_VIA0 $T=144550 48080 0 0 $X=144300 $Y=47840
X2646 1 DigitalLDOLogic_VIA0 $T=144550 53520 0 0 $X=144300 $Y=53280
X2647 1 DigitalLDOLogic_VIA0 $T=144550 58960 0 0 $X=144300 $Y=58720
X2648 2 DigitalLDOLogic_VIA0 $T=146390 12720 0 0 $X=146140 $Y=12480
X2649 2 DigitalLDOLogic_VIA0 $T=146390 18160 0 0 $X=146140 $Y=17920
X2650 2 DigitalLDOLogic_VIA0 $T=146390 23600 0 0 $X=146140 $Y=23360
X2651 2 DigitalLDOLogic_VIA0 $T=146390 29040 0 0 $X=146140 $Y=28800
X2652 2 DigitalLDOLogic_VIA0 $T=146390 34480 0 0 $X=146140 $Y=34240
X2653 2 DigitalLDOLogic_VIA0 $T=146390 39920 0 0 $X=146140 $Y=39680
X2654 2 DigitalLDOLogic_VIA0 $T=146390 45360 0 0 $X=146140 $Y=45120
X2655 2 DigitalLDOLogic_VIA0 $T=146390 50800 0 0 $X=146140 $Y=50560
X2656 2 DigitalLDOLogic_VIA0 $T=146390 56240 0 0 $X=146140 $Y=56000
X2657 1 DigitalLDOLogic_VIA0 $T=147310 15440 0 0 $X=147060 $Y=15200
X2658 1 DigitalLDOLogic_VIA0 $T=147310 20880 0 0 $X=147060 $Y=20640
X2659 1 DigitalLDOLogic_VIA0 $T=147310 26320 0 0 $X=147060 $Y=26080
X2660 1 DigitalLDOLogic_VIA0 $T=147310 31760 0 0 $X=147060 $Y=31520
X2661 1 DigitalLDOLogic_VIA0 $T=147310 37200 0 0 $X=147060 $Y=36960
X2662 1 DigitalLDOLogic_VIA0 $T=147310 42640 0 0 $X=147060 $Y=42400
X2663 1 DigitalLDOLogic_VIA0 $T=147310 48080 0 0 $X=147060 $Y=47840
X2664 1 DigitalLDOLogic_VIA0 $T=147310 53520 0 0 $X=147060 $Y=53280
X2665 1 DigitalLDOLogic_VIA0 $T=147310 58960 0 0 $X=147060 $Y=58720
X2666 2 DigitalLDOLogic_VIA0 $T=149150 12720 0 0 $X=148900 $Y=12480
X2667 2 DigitalLDOLogic_VIA0 $T=149150 18160 0 0 $X=148900 $Y=17920
X2668 2 DigitalLDOLogic_VIA0 $T=149150 23600 0 0 $X=148900 $Y=23360
X2669 2 DigitalLDOLogic_VIA0 $T=149150 29040 0 0 $X=148900 $Y=28800
X2670 2 DigitalLDOLogic_VIA0 $T=149150 34480 0 0 $X=148900 $Y=34240
X2671 2 DigitalLDOLogic_VIA0 $T=149150 39920 0 0 $X=148900 $Y=39680
X2672 2 DigitalLDOLogic_VIA0 $T=149150 45360 0 0 $X=148900 $Y=45120
X2673 2 DigitalLDOLogic_VIA0 $T=149150 50800 0 0 $X=148900 $Y=50560
X2674 2 DigitalLDOLogic_VIA0 $T=149150 56240 0 0 $X=148900 $Y=56000
X2675 1 DigitalLDOLogic_VIA0 $T=150070 15440 0 0 $X=149820 $Y=15200
X2676 1 DigitalLDOLogic_VIA0 $T=150070 20880 0 0 $X=149820 $Y=20640
X2677 1 DigitalLDOLogic_VIA0 $T=150070 26320 0 0 $X=149820 $Y=26080
X2678 1 DigitalLDOLogic_VIA0 $T=150070 31760 0 0 $X=149820 $Y=31520
X2679 1 DigitalLDOLogic_VIA0 $T=150070 37200 0 0 $X=149820 $Y=36960
X2680 1 DigitalLDOLogic_VIA0 $T=150070 42640 0 0 $X=149820 $Y=42400
X2681 1 DigitalLDOLogic_VIA0 $T=150070 48080 0 0 $X=149820 $Y=47840
X2682 1 DigitalLDOLogic_VIA0 $T=150070 53520 0 0 $X=149820 $Y=53280
X2683 1 DigitalLDOLogic_VIA0 $T=150070 58960 0 0 $X=149820 $Y=58720
X2684 2 DigitalLDOLogic_VIA0 $T=151910 12720 0 0 $X=151660 $Y=12480
X2685 2 DigitalLDOLogic_VIA0 $T=151910 18160 0 0 $X=151660 $Y=17920
X2686 2 DigitalLDOLogic_VIA0 $T=151910 23600 0 0 $X=151660 $Y=23360
X2687 2 DigitalLDOLogic_VIA0 $T=151910 29040 0 0 $X=151660 $Y=28800
X2688 2 DigitalLDOLogic_VIA0 $T=151910 34480 0 0 $X=151660 $Y=34240
X2689 2 DigitalLDOLogic_VIA0 $T=151910 39920 0 0 $X=151660 $Y=39680
X2690 2 DigitalLDOLogic_VIA0 $T=151910 45360 0 0 $X=151660 $Y=45120
X2691 2 DigitalLDOLogic_VIA0 $T=151910 50800 0 0 $X=151660 $Y=50560
X2692 2 DigitalLDOLogic_VIA0 $T=151910 56240 0 0 $X=151660 $Y=56000
X2693 1 DigitalLDOLogic_VIA0 $T=152830 15440 0 0 $X=152580 $Y=15200
X2694 1 DigitalLDOLogic_VIA0 $T=152830 20880 0 0 $X=152580 $Y=20640
X2695 1 DigitalLDOLogic_VIA0 $T=152830 26320 0 0 $X=152580 $Y=26080
X2696 1 DigitalLDOLogic_VIA0 $T=152830 31760 0 0 $X=152580 $Y=31520
X2697 1 DigitalLDOLogic_VIA0 $T=152830 37200 0 0 $X=152580 $Y=36960
X2698 1 DigitalLDOLogic_VIA0 $T=152830 42640 0 0 $X=152580 $Y=42400
X2699 1 DigitalLDOLogic_VIA0 $T=152830 48080 0 0 $X=152580 $Y=47840
X2700 1 DigitalLDOLogic_VIA0 $T=152830 53520 0 0 $X=152580 $Y=53280
X2701 1 DigitalLDOLogic_VIA0 $T=152830 58960 0 0 $X=152580 $Y=58720
X2702 2 DigitalLDOLogic_VIA0 $T=154670 12720 0 0 $X=154420 $Y=12480
X2703 2 DigitalLDOLogic_VIA0 $T=154670 18160 0 0 $X=154420 $Y=17920
X2704 2 DigitalLDOLogic_VIA0 $T=154670 23600 0 0 $X=154420 $Y=23360
X2705 2 DigitalLDOLogic_VIA0 $T=154670 29040 0 0 $X=154420 $Y=28800
X2706 2 DigitalLDOLogic_VIA0 $T=154670 34480 0 0 $X=154420 $Y=34240
X2707 2 DigitalLDOLogic_VIA0 $T=154670 39920 0 0 $X=154420 $Y=39680
X2708 2 DigitalLDOLogic_VIA0 $T=154670 45360 0 0 $X=154420 $Y=45120
X2709 2 DigitalLDOLogic_VIA0 $T=154670 50800 0 0 $X=154420 $Y=50560
X2710 2 DigitalLDOLogic_VIA0 $T=154670 56240 0 0 $X=154420 $Y=56000
X2711 1 DigitalLDOLogic_VIA0 $T=155590 15440 0 0 $X=155340 $Y=15200
X2712 1 DigitalLDOLogic_VIA0 $T=155590 20880 0 0 $X=155340 $Y=20640
X2713 1 DigitalLDOLogic_VIA0 $T=155590 26320 0 0 $X=155340 $Y=26080
X2714 1 DigitalLDOLogic_VIA0 $T=155590 31760 0 0 $X=155340 $Y=31520
X2715 1 DigitalLDOLogic_VIA0 $T=155590 37200 0 0 $X=155340 $Y=36960
X2716 1 DigitalLDOLogic_VIA0 $T=155590 42640 0 0 $X=155340 $Y=42400
X2717 1 DigitalLDOLogic_VIA0 $T=155590 48080 0 0 $X=155340 $Y=47840
X2718 1 DigitalLDOLogic_VIA0 $T=155590 53520 0 0 $X=155340 $Y=53280
X2719 1 DigitalLDOLogic_VIA0 $T=155590 58960 0 0 $X=155340 $Y=58720
X2720 2 DigitalLDOLogic_VIA0 $T=157430 12720 0 0 $X=157180 $Y=12480
X2721 2 DigitalLDOLogic_VIA0 $T=157430 18160 0 0 $X=157180 $Y=17920
X2722 2 DigitalLDOLogic_VIA0 $T=157430 23600 0 0 $X=157180 $Y=23360
X2723 2 DigitalLDOLogic_VIA0 $T=157430 29040 0 0 $X=157180 $Y=28800
X2724 2 DigitalLDOLogic_VIA0 $T=157430 34480 0 0 $X=157180 $Y=34240
X2725 2 DigitalLDOLogic_VIA0 $T=157430 39920 0 0 $X=157180 $Y=39680
X2726 2 DigitalLDOLogic_VIA0 $T=157430 45360 0 0 $X=157180 $Y=45120
X2727 2 DigitalLDOLogic_VIA0 $T=157430 50800 0 0 $X=157180 $Y=50560
X2728 2 DigitalLDOLogic_VIA0 $T=157430 56240 0 0 $X=157180 $Y=56000
X2729 1 DigitalLDOLogic_VIA0 $T=158350 15440 0 0 $X=158100 $Y=15200
X2730 1 DigitalLDOLogic_VIA0 $T=158350 20880 0 0 $X=158100 $Y=20640
X2731 1 DigitalLDOLogic_VIA0 $T=158350 26320 0 0 $X=158100 $Y=26080
X2732 1 DigitalLDOLogic_VIA0 $T=158350 31760 0 0 $X=158100 $Y=31520
X2733 1 DigitalLDOLogic_VIA0 $T=158350 37200 0 0 $X=158100 $Y=36960
X2734 1 DigitalLDOLogic_VIA0 $T=158350 42640 0 0 $X=158100 $Y=42400
X2735 1 DigitalLDOLogic_VIA0 $T=158350 48080 0 0 $X=158100 $Y=47840
X2736 1 DigitalLDOLogic_VIA0 $T=158350 53520 0 0 $X=158100 $Y=53280
X2737 1 DigitalLDOLogic_VIA0 $T=158350 58960 0 0 $X=158100 $Y=58720
X2738 2 DigitalLDOLogic_VIA0 $T=160190 12720 0 0 $X=159940 $Y=12480
X2739 2 DigitalLDOLogic_VIA0 $T=160190 18160 0 0 $X=159940 $Y=17920
X2740 2 DigitalLDOLogic_VIA0 $T=160190 23600 0 0 $X=159940 $Y=23360
X2741 2 DigitalLDOLogic_VIA0 $T=160190 29040 0 0 $X=159940 $Y=28800
X2742 2 DigitalLDOLogic_VIA0 $T=160190 34480 0 0 $X=159940 $Y=34240
X2743 2 DigitalLDOLogic_VIA0 $T=160190 39920 0 0 $X=159940 $Y=39680
X2744 2 DigitalLDOLogic_VIA0 $T=160190 45360 0 0 $X=159940 $Y=45120
X2745 2 DigitalLDOLogic_VIA0 $T=160190 50800 0 0 $X=159940 $Y=50560
X2746 2 DigitalLDOLogic_VIA0 $T=160190 56240 0 0 $X=159940 $Y=56000
X2747 1 DigitalLDOLogic_VIA0 $T=161110 15440 0 0 $X=160860 $Y=15200
X2748 1 DigitalLDOLogic_VIA0 $T=161110 20880 0 0 $X=160860 $Y=20640
X2749 1 DigitalLDOLogic_VIA0 $T=161110 26320 0 0 $X=160860 $Y=26080
X2750 1 DigitalLDOLogic_VIA0 $T=161110 31760 0 0 $X=160860 $Y=31520
X2751 1 DigitalLDOLogic_VIA0 $T=161110 37200 0 0 $X=160860 $Y=36960
X2752 1 DigitalLDOLogic_VIA0 $T=161110 42640 0 0 $X=160860 $Y=42400
X2753 1 DigitalLDOLogic_VIA0 $T=161110 48080 0 0 $X=160860 $Y=47840
X2754 1 DigitalLDOLogic_VIA0 $T=161110 53520 0 0 $X=160860 $Y=53280
X2755 1 DigitalLDOLogic_VIA0 $T=161110 58960 0 0 $X=160860 $Y=58720
X2756 2 DigitalLDOLogic_VIA0 $T=162950 12720 0 0 $X=162700 $Y=12480
X2757 2 DigitalLDOLogic_VIA0 $T=162950 18160 0 0 $X=162700 $Y=17920
X2758 2 DigitalLDOLogic_VIA0 $T=162950 23600 0 0 $X=162700 $Y=23360
X2759 2 DigitalLDOLogic_VIA0 $T=162950 29040 0 0 $X=162700 $Y=28800
X2760 2 DigitalLDOLogic_VIA0 $T=162950 34480 0 0 $X=162700 $Y=34240
X2761 2 DigitalLDOLogic_VIA0 $T=162950 39920 0 0 $X=162700 $Y=39680
X2762 2 DigitalLDOLogic_VIA0 $T=162950 45360 0 0 $X=162700 $Y=45120
X2763 2 DigitalLDOLogic_VIA0 $T=162950 50800 0 0 $X=162700 $Y=50560
X2764 2 DigitalLDOLogic_VIA0 $T=162950 56240 0 0 $X=162700 $Y=56000
X2765 1 DigitalLDOLogic_VIA0 $T=163870 15440 0 0 $X=163620 $Y=15200
X2766 1 DigitalLDOLogic_VIA0 $T=163870 20880 0 0 $X=163620 $Y=20640
X2767 1 DigitalLDOLogic_VIA0 $T=163870 26320 0 0 $X=163620 $Y=26080
X2768 1 DigitalLDOLogic_VIA0 $T=163870 31760 0 0 $X=163620 $Y=31520
X2769 1 DigitalLDOLogic_VIA0 $T=163870 37200 0 0 $X=163620 $Y=36960
X2770 1 DigitalLDOLogic_VIA0 $T=163870 42640 0 0 $X=163620 $Y=42400
X2771 1 DigitalLDOLogic_VIA0 $T=163870 48080 0 0 $X=163620 $Y=47840
X2772 1 DigitalLDOLogic_VIA0 $T=163870 53520 0 0 $X=163620 $Y=53280
X2773 1 DigitalLDOLogic_VIA0 $T=163870 58960 0 0 $X=163620 $Y=58720
X2774 2 DigitalLDOLogic_VIA0 $T=165710 12720 0 0 $X=165460 $Y=12480
X2775 2 DigitalLDOLogic_VIA0 $T=165710 18160 0 0 $X=165460 $Y=17920
X2776 2 DigitalLDOLogic_VIA0 $T=165710 23600 0 0 $X=165460 $Y=23360
X2777 2 DigitalLDOLogic_VIA0 $T=165710 29040 0 0 $X=165460 $Y=28800
X2778 2 DigitalLDOLogic_VIA0 $T=165710 34480 0 0 $X=165460 $Y=34240
X2779 2 DigitalLDOLogic_VIA0 $T=165710 39920 0 0 $X=165460 $Y=39680
X2780 2 DigitalLDOLogic_VIA0 $T=165710 45360 0 0 $X=165460 $Y=45120
X2781 2 DigitalLDOLogic_VIA0 $T=165710 50800 0 0 $X=165460 $Y=50560
X2782 2 DigitalLDOLogic_VIA0 $T=165710 56240 0 0 $X=165460 $Y=56000
X2783 1 DigitalLDOLogic_VIA0 $T=166630 15440 0 0 $X=166380 $Y=15200
X2784 1 DigitalLDOLogic_VIA0 $T=166630 20880 0 0 $X=166380 $Y=20640
X2785 1 DigitalLDOLogic_VIA0 $T=166630 26320 0 0 $X=166380 $Y=26080
X2786 1 DigitalLDOLogic_VIA0 $T=166630 31760 0 0 $X=166380 $Y=31520
X2787 1 DigitalLDOLogic_VIA0 $T=166630 37200 0 0 $X=166380 $Y=36960
X2788 1 DigitalLDOLogic_VIA0 $T=166630 42640 0 0 $X=166380 $Y=42400
X2789 1 DigitalLDOLogic_VIA0 $T=166630 48080 0 0 $X=166380 $Y=47840
X2790 1 DigitalLDOLogic_VIA0 $T=166630 53520 0 0 $X=166380 $Y=53280
X2791 1 DigitalLDOLogic_VIA0 $T=166630 58960 0 0 $X=166380 $Y=58720
X2792 2 DigitalLDOLogic_VIA0 $T=168470 12720 0 0 $X=168220 $Y=12480
X2793 2 DigitalLDOLogic_VIA0 $T=168470 18160 0 0 $X=168220 $Y=17920
X2794 2 DigitalLDOLogic_VIA0 $T=168470 23600 0 0 $X=168220 $Y=23360
X2795 2 DigitalLDOLogic_VIA0 $T=168470 29040 0 0 $X=168220 $Y=28800
X2796 2 DigitalLDOLogic_VIA0 $T=168470 34480 0 0 $X=168220 $Y=34240
X2797 2 DigitalLDOLogic_VIA0 $T=168470 39920 0 0 $X=168220 $Y=39680
X2798 2 DigitalLDOLogic_VIA0 $T=168470 45360 0 0 $X=168220 $Y=45120
X2799 2 DigitalLDOLogic_VIA0 $T=168470 50800 0 0 $X=168220 $Y=50560
X2800 2 DigitalLDOLogic_VIA0 $T=168470 56240 0 0 $X=168220 $Y=56000
X2801 1 DigitalLDOLogic_VIA0 $T=169390 15440 0 0 $X=169140 $Y=15200
X2802 1 DigitalLDOLogic_VIA0 $T=169390 20880 0 0 $X=169140 $Y=20640
X2803 1 DigitalLDOLogic_VIA0 $T=169390 26320 0 0 $X=169140 $Y=26080
X2804 1 DigitalLDOLogic_VIA0 $T=169390 31760 0 0 $X=169140 $Y=31520
X2805 1 DigitalLDOLogic_VIA0 $T=169390 37200 0 0 $X=169140 $Y=36960
X2806 1 DigitalLDOLogic_VIA0 $T=169390 42640 0 0 $X=169140 $Y=42400
X2807 1 DigitalLDOLogic_VIA0 $T=169390 48080 0 0 $X=169140 $Y=47840
X2808 1 DigitalLDOLogic_VIA0 $T=169390 53520 0 0 $X=169140 $Y=53280
X2809 1 DigitalLDOLogic_VIA0 $T=169390 58960 0 0 $X=169140 $Y=58720
X2810 2 DigitalLDOLogic_VIA0 $T=171230 12720 0 0 $X=170980 $Y=12480
X2811 2 DigitalLDOLogic_VIA0 $T=171230 18160 0 0 $X=170980 $Y=17920
X2812 2 DigitalLDOLogic_VIA0 $T=171230 23600 0 0 $X=170980 $Y=23360
X2813 2 DigitalLDOLogic_VIA0 $T=171230 29040 0 0 $X=170980 $Y=28800
X2814 2 DigitalLDOLogic_VIA0 $T=171230 34480 0 0 $X=170980 $Y=34240
X2815 2 DigitalLDOLogic_VIA0 $T=171230 39920 0 0 $X=170980 $Y=39680
X2816 2 DigitalLDOLogic_VIA0 $T=171230 45360 0 0 $X=170980 $Y=45120
X2817 2 DigitalLDOLogic_VIA0 $T=171230 50800 0 0 $X=170980 $Y=50560
X2818 2 DigitalLDOLogic_VIA0 $T=171230 56240 0 0 $X=170980 $Y=56000
X2819 1 DigitalLDOLogic_VIA0 $T=172150 15440 0 0 $X=171900 $Y=15200
X2820 1 DigitalLDOLogic_VIA0 $T=172150 20880 0 0 $X=171900 $Y=20640
X2821 1 DigitalLDOLogic_VIA0 $T=172150 26320 0 0 $X=171900 $Y=26080
X2822 1 DigitalLDOLogic_VIA0 $T=172150 31760 0 0 $X=171900 $Y=31520
X2823 1 DigitalLDOLogic_VIA0 $T=172150 37200 0 0 $X=171900 $Y=36960
X2824 1 DigitalLDOLogic_VIA0 $T=172150 42640 0 0 $X=171900 $Y=42400
X2825 1 DigitalLDOLogic_VIA0 $T=172150 48080 0 0 $X=171900 $Y=47840
X2826 1 DigitalLDOLogic_VIA0 $T=172150 53520 0 0 $X=171900 $Y=53280
X2827 1 DigitalLDOLogic_VIA0 $T=172150 58960 0 0 $X=171900 $Y=58720
X2828 2 DigitalLDOLogic_VIA0 $T=173990 12720 0 0 $X=173740 $Y=12480
X2829 2 DigitalLDOLogic_VIA0 $T=173990 18160 0 0 $X=173740 $Y=17920
X2830 2 DigitalLDOLogic_VIA0 $T=173990 23600 0 0 $X=173740 $Y=23360
X2831 2 DigitalLDOLogic_VIA0 $T=173990 29040 0 0 $X=173740 $Y=28800
X2832 2 DigitalLDOLogic_VIA0 $T=173990 34480 0 0 $X=173740 $Y=34240
X2833 2 DigitalLDOLogic_VIA0 $T=173990 39920 0 0 $X=173740 $Y=39680
X2834 2 DigitalLDOLogic_VIA0 $T=173990 45360 0 0 $X=173740 $Y=45120
X2835 2 DigitalLDOLogic_VIA0 $T=173990 50800 0 0 $X=173740 $Y=50560
X2836 2 DigitalLDOLogic_VIA0 $T=173990 56240 0 0 $X=173740 $Y=56000
X2837 1 DigitalLDOLogic_VIA0 $T=174910 15440 0 0 $X=174660 $Y=15200
X2838 1 DigitalLDOLogic_VIA0 $T=174910 20880 0 0 $X=174660 $Y=20640
X2839 1 DigitalLDOLogic_VIA0 $T=174910 26320 0 0 $X=174660 $Y=26080
X2840 1 DigitalLDOLogic_VIA0 $T=174910 31760 0 0 $X=174660 $Y=31520
X2841 1 DigitalLDOLogic_VIA0 $T=174910 37200 0 0 $X=174660 $Y=36960
X2842 1 DigitalLDOLogic_VIA0 $T=174910 42640 0 0 $X=174660 $Y=42400
X2843 1 DigitalLDOLogic_VIA0 $T=174910 48080 0 0 $X=174660 $Y=47840
X2844 1 DigitalLDOLogic_VIA0 $T=174910 53520 0 0 $X=174660 $Y=53280
X2845 1 DigitalLDOLogic_VIA0 $T=174910 58960 0 0 $X=174660 $Y=58720
X2846 2 DigitalLDOLogic_VIA0 $T=176750 12720 0 0 $X=176500 $Y=12480
X2847 2 DigitalLDOLogic_VIA0 $T=176750 18160 0 0 $X=176500 $Y=17920
X2848 2 DigitalLDOLogic_VIA0 $T=176750 23600 0 0 $X=176500 $Y=23360
X2849 2 DigitalLDOLogic_VIA0 $T=176750 29040 0 0 $X=176500 $Y=28800
X2850 2 DigitalLDOLogic_VIA0 $T=176750 34480 0 0 $X=176500 $Y=34240
X2851 2 DigitalLDOLogic_VIA0 $T=176750 39920 0 0 $X=176500 $Y=39680
X2852 2 DigitalLDOLogic_VIA0 $T=176750 45360 0 0 $X=176500 $Y=45120
X2853 2 DigitalLDOLogic_VIA0 $T=176750 50800 0 0 $X=176500 $Y=50560
X2854 2 DigitalLDOLogic_VIA0 $T=176750 56240 0 0 $X=176500 $Y=56000
X2855 1 DigitalLDOLogic_VIA0 $T=177670 15440 0 0 $X=177420 $Y=15200
X2856 1 DigitalLDOLogic_VIA0 $T=177670 20880 0 0 $X=177420 $Y=20640
X2857 1 DigitalLDOLogic_VIA0 $T=177670 26320 0 0 $X=177420 $Y=26080
X2858 1 DigitalLDOLogic_VIA0 $T=177670 31760 0 0 $X=177420 $Y=31520
X2859 1 DigitalLDOLogic_VIA0 $T=177670 37200 0 0 $X=177420 $Y=36960
X2860 1 DigitalLDOLogic_VIA0 $T=177670 42640 0 0 $X=177420 $Y=42400
X2861 1 DigitalLDOLogic_VIA0 $T=177670 48080 0 0 $X=177420 $Y=47840
X2862 1 DigitalLDOLogic_VIA0 $T=177670 53520 0 0 $X=177420 $Y=53280
X2863 1 DigitalLDOLogic_VIA0 $T=177670 58960 0 0 $X=177420 $Y=58720
X2864 2 DigitalLDOLogic_VIA0 $T=179510 12720 0 0 $X=179260 $Y=12480
X2865 2 DigitalLDOLogic_VIA0 $T=179510 18160 0 0 $X=179260 $Y=17920
X2866 2 DigitalLDOLogic_VIA0 $T=179510 23600 0 0 $X=179260 $Y=23360
X2867 2 DigitalLDOLogic_VIA0 $T=179510 29040 0 0 $X=179260 $Y=28800
X2868 2 DigitalLDOLogic_VIA0 $T=179510 34480 0 0 $X=179260 $Y=34240
X2869 2 DigitalLDOLogic_VIA0 $T=179510 39920 0 0 $X=179260 $Y=39680
X2870 2 DigitalLDOLogic_VIA0 $T=179510 45360 0 0 $X=179260 $Y=45120
X2871 2 DigitalLDOLogic_VIA0 $T=179510 50800 0 0 $X=179260 $Y=50560
X2872 2 DigitalLDOLogic_VIA0 $T=179510 56240 0 0 $X=179260 $Y=56000
X2873 1 DigitalLDOLogic_VIA0 $T=180430 15440 0 0 $X=180180 $Y=15200
X2874 1 DigitalLDOLogic_VIA0 $T=180430 20880 0 0 $X=180180 $Y=20640
X2875 1 DigitalLDOLogic_VIA0 $T=180430 26320 0 0 $X=180180 $Y=26080
X2876 1 DigitalLDOLogic_VIA0 $T=180430 31760 0 0 $X=180180 $Y=31520
X2877 1 DigitalLDOLogic_VIA0 $T=180430 37200 0 0 $X=180180 $Y=36960
X2878 1 DigitalLDOLogic_VIA0 $T=180430 42640 0 0 $X=180180 $Y=42400
X2879 1 DigitalLDOLogic_VIA0 $T=180430 48080 0 0 $X=180180 $Y=47840
X2880 1 DigitalLDOLogic_VIA0 $T=180430 53520 0 0 $X=180180 $Y=53280
X2881 1 DigitalLDOLogic_VIA0 $T=180430 58960 0 0 $X=180180 $Y=58720
X2882 2 DigitalLDOLogic_VIA0 $T=182270 12720 0 0 $X=182020 $Y=12480
X2883 2 DigitalLDOLogic_VIA0 $T=182270 18160 0 0 $X=182020 $Y=17920
X2884 2 DigitalLDOLogic_VIA0 $T=182270 23600 0 0 $X=182020 $Y=23360
X2885 2 DigitalLDOLogic_VIA0 $T=182270 29040 0 0 $X=182020 $Y=28800
X2886 2 DigitalLDOLogic_VIA0 $T=182270 34480 0 0 $X=182020 $Y=34240
X2887 2 DigitalLDOLogic_VIA0 $T=182270 39920 0 0 $X=182020 $Y=39680
X2888 2 DigitalLDOLogic_VIA0 $T=182270 45360 0 0 $X=182020 $Y=45120
X2889 2 DigitalLDOLogic_VIA0 $T=182270 50800 0 0 $X=182020 $Y=50560
X2890 2 DigitalLDOLogic_VIA0 $T=182270 56240 0 0 $X=182020 $Y=56000
X2891 1 DigitalLDOLogic_VIA0 $T=183190 15440 0 0 $X=182940 $Y=15200
X2892 1 DigitalLDOLogic_VIA0 $T=183190 20880 0 0 $X=182940 $Y=20640
X2893 1 DigitalLDOLogic_VIA0 $T=183190 26320 0 0 $X=182940 $Y=26080
X2894 1 DigitalLDOLogic_VIA0 $T=183190 31760 0 0 $X=182940 $Y=31520
X2895 1 DigitalLDOLogic_VIA0 $T=183190 37200 0 0 $X=182940 $Y=36960
X2896 1 DigitalLDOLogic_VIA0 $T=183190 42640 0 0 $X=182940 $Y=42400
X2897 1 DigitalLDOLogic_VIA0 $T=183190 48080 0 0 $X=182940 $Y=47840
X2898 1 DigitalLDOLogic_VIA0 $T=183190 53520 0 0 $X=182940 $Y=53280
X2899 1 DigitalLDOLogic_VIA0 $T=183190 58960 0 0 $X=182940 $Y=58720
X2900 2 DigitalLDOLogic_VIA0 $T=185030 12720 0 0 $X=184780 $Y=12480
X2901 2 DigitalLDOLogic_VIA0 $T=185030 18160 0 0 $X=184780 $Y=17920
X2902 2 DigitalLDOLogic_VIA0 $T=185030 23600 0 0 $X=184780 $Y=23360
X2903 2 DigitalLDOLogic_VIA0 $T=185030 29040 0 0 $X=184780 $Y=28800
X2904 2 DigitalLDOLogic_VIA0 $T=185030 34480 0 0 $X=184780 $Y=34240
X2905 2 DigitalLDOLogic_VIA0 $T=185030 39920 0 0 $X=184780 $Y=39680
X2906 2 DigitalLDOLogic_VIA0 $T=185030 45360 0 0 $X=184780 $Y=45120
X2907 2 DigitalLDOLogic_VIA0 $T=185030 50800 0 0 $X=184780 $Y=50560
X2908 2 DigitalLDOLogic_VIA0 $T=185030 56240 0 0 $X=184780 $Y=56000
X2909 1 DigitalLDOLogic_VIA0 $T=185950 15440 0 0 $X=185700 $Y=15200
X2910 1 DigitalLDOLogic_VIA0 $T=185950 20880 0 0 $X=185700 $Y=20640
X2911 1 DigitalLDOLogic_VIA0 $T=185950 26320 0 0 $X=185700 $Y=26080
X2912 1 DigitalLDOLogic_VIA0 $T=185950 31760 0 0 $X=185700 $Y=31520
X2913 1 DigitalLDOLogic_VIA0 $T=185950 37200 0 0 $X=185700 $Y=36960
X2914 1 DigitalLDOLogic_VIA0 $T=185950 42640 0 0 $X=185700 $Y=42400
X2915 1 DigitalLDOLogic_VIA0 $T=185950 48080 0 0 $X=185700 $Y=47840
X2916 1 DigitalLDOLogic_VIA0 $T=185950 53520 0 0 $X=185700 $Y=53280
X2917 1 DigitalLDOLogic_VIA0 $T=185950 58960 0 0 $X=185700 $Y=58720
X2918 2 DigitalLDOLogic_VIA0 $T=187790 12720 0 0 $X=187540 $Y=12480
X2919 2 DigitalLDOLogic_VIA0 $T=187790 18160 0 0 $X=187540 $Y=17920
X2920 2 DigitalLDOLogic_VIA0 $T=187790 23600 0 0 $X=187540 $Y=23360
X2921 2 DigitalLDOLogic_VIA0 $T=187790 29040 0 0 $X=187540 $Y=28800
X2922 2 DigitalLDOLogic_VIA0 $T=187790 34480 0 0 $X=187540 $Y=34240
X2923 2 DigitalLDOLogic_VIA0 $T=187790 39920 0 0 $X=187540 $Y=39680
X2924 2 DigitalLDOLogic_VIA0 $T=187790 45360 0 0 $X=187540 $Y=45120
X2925 2 DigitalLDOLogic_VIA0 $T=187790 50800 0 0 $X=187540 $Y=50560
X2926 2 DigitalLDOLogic_VIA0 $T=187790 56240 0 0 $X=187540 $Y=56000
X2927 1 DigitalLDOLogic_VIA0 $T=188710 15440 0 0 $X=188460 $Y=15200
X2928 1 DigitalLDOLogic_VIA0 $T=188710 20880 0 0 $X=188460 $Y=20640
X2929 1 DigitalLDOLogic_VIA0 $T=188710 26320 0 0 $X=188460 $Y=26080
X2930 1 DigitalLDOLogic_VIA0 $T=188710 31760 0 0 $X=188460 $Y=31520
X2931 1 DigitalLDOLogic_VIA0 $T=188710 37200 0 0 $X=188460 $Y=36960
X2932 1 DigitalLDOLogic_VIA0 $T=188710 42640 0 0 $X=188460 $Y=42400
X2933 1 DigitalLDOLogic_VIA0 $T=188710 48080 0 0 $X=188460 $Y=47840
X2934 1 DigitalLDOLogic_VIA0 $T=188710 53520 0 0 $X=188460 $Y=53280
X2935 1 DigitalLDOLogic_VIA0 $T=188710 58960 0 0 $X=188460 $Y=58720
X2936 2 DigitalLDOLogic_VIA1 $T=11150 11700 0 0 $X=10900 $Y=11470
X2937 2 DigitalLDOLogic_VIA1 $T=11150 15780 0 0 $X=10900 $Y=15550
X2938 2 DigitalLDOLogic_VIA1 $T=11150 19860 0 0 $X=10900 $Y=19630
X2939 2 DigitalLDOLogic_VIA1 $T=11150 23940 0 0 $X=10900 $Y=23710
X2940 2 DigitalLDOLogic_VIA1 $T=11150 28020 0 0 $X=10900 $Y=27790
X2941 2 DigitalLDOLogic_VIA1 $T=11150 32100 0 0 $X=10900 $Y=31870
X2942 2 DigitalLDOLogic_VIA1 $T=11150 36180 0 0 $X=10900 $Y=35950
X2943 2 DigitalLDOLogic_VIA1 $T=11150 40260 0 0 $X=10900 $Y=40030
X2944 2 DigitalLDOLogic_VIA1 $T=11150 44340 0 0 $X=10900 $Y=44110
X2945 2 DigitalLDOLogic_VIA1 $T=11150 48420 0 0 $X=10900 $Y=48190
X2946 2 DigitalLDOLogic_VIA1 $T=11150 52500 0 0 $X=10900 $Y=52270
X2947 2 DigitalLDOLogic_VIA1 $T=11150 56580 0 0 $X=10900 $Y=56350
X2948 1 DigitalLDOLogic_VIA1 $T=12070 13060 0 0 $X=11820 $Y=12830
X2949 1 DigitalLDOLogic_VIA1 $T=12070 17140 0 0 $X=11820 $Y=16910
X2950 1 DigitalLDOLogic_VIA1 $T=12070 21220 0 0 $X=11820 $Y=20990
X2951 1 DigitalLDOLogic_VIA1 $T=12070 25300 0 0 $X=11820 $Y=25070
X2952 1 DigitalLDOLogic_VIA1 $T=12070 29380 0 0 $X=11820 $Y=29150
X2953 1 DigitalLDOLogic_VIA1 $T=12070 33460 0 0 $X=11820 $Y=33230
X2954 1 DigitalLDOLogic_VIA1 $T=12070 37540 0 0 $X=11820 $Y=37310
X2955 1 DigitalLDOLogic_VIA1 $T=12070 41620 0 0 $X=11820 $Y=41390
X2956 1 DigitalLDOLogic_VIA1 $T=12070 45700 0 0 $X=11820 $Y=45470
X2957 1 DigitalLDOLogic_VIA1 $T=12070 49780 0 0 $X=11820 $Y=49550
X2958 1 DigitalLDOLogic_VIA1 $T=12070 53860 0 0 $X=11820 $Y=53630
X2959 1 DigitalLDOLogic_VIA1 $T=12070 57940 0 0 $X=11820 $Y=57710
X2960 2 DigitalLDOLogic_VIA1 $T=13910 11700 0 0 $X=13660 $Y=11470
X2961 2 DigitalLDOLogic_VIA1 $T=13910 15780 0 0 $X=13660 $Y=15550
X2962 2 DigitalLDOLogic_VIA1 $T=13910 19860 0 0 $X=13660 $Y=19630
X2963 2 DigitalLDOLogic_VIA1 $T=13910 23940 0 0 $X=13660 $Y=23710
X2964 2 DigitalLDOLogic_VIA1 $T=13910 28020 0 0 $X=13660 $Y=27790
X2965 2 DigitalLDOLogic_VIA1 $T=13910 32100 0 0 $X=13660 $Y=31870
X2966 2 DigitalLDOLogic_VIA1 $T=13910 36180 0 0 $X=13660 $Y=35950
X2967 2 DigitalLDOLogic_VIA1 $T=13910 40260 0 0 $X=13660 $Y=40030
X2968 2 DigitalLDOLogic_VIA1 $T=13910 44340 0 0 $X=13660 $Y=44110
X2969 2 DigitalLDOLogic_VIA1 $T=13910 48420 0 0 $X=13660 $Y=48190
X2970 2 DigitalLDOLogic_VIA1 $T=13910 52500 0 0 $X=13660 $Y=52270
X2971 2 DigitalLDOLogic_VIA1 $T=13910 56580 0 0 $X=13660 $Y=56350
X2972 1 DigitalLDOLogic_VIA1 $T=14830 13060 0 0 $X=14580 $Y=12830
X2973 1 DigitalLDOLogic_VIA1 $T=14830 17140 0 0 $X=14580 $Y=16910
X2974 1 DigitalLDOLogic_VIA1 $T=14830 21220 0 0 $X=14580 $Y=20990
X2975 1 DigitalLDOLogic_VIA1 $T=14830 25300 0 0 $X=14580 $Y=25070
X2976 1 DigitalLDOLogic_VIA1 $T=14830 29380 0 0 $X=14580 $Y=29150
X2977 1 DigitalLDOLogic_VIA1 $T=14830 33460 0 0 $X=14580 $Y=33230
X2978 1 DigitalLDOLogic_VIA1 $T=14830 37540 0 0 $X=14580 $Y=37310
X2979 1 DigitalLDOLogic_VIA1 $T=14830 41620 0 0 $X=14580 $Y=41390
X2980 1 DigitalLDOLogic_VIA1 $T=14830 45700 0 0 $X=14580 $Y=45470
X2981 1 DigitalLDOLogic_VIA1 $T=14830 49780 0 0 $X=14580 $Y=49550
X2982 1 DigitalLDOLogic_VIA1 $T=14830 53860 0 0 $X=14580 $Y=53630
X2983 1 DigitalLDOLogic_VIA1 $T=14830 57940 0 0 $X=14580 $Y=57710
X2984 2 DigitalLDOLogic_VIA1 $T=16670 11700 0 0 $X=16420 $Y=11470
X2985 2 DigitalLDOLogic_VIA1 $T=16670 15780 0 0 $X=16420 $Y=15550
X2986 2 DigitalLDOLogic_VIA1 $T=16670 19860 0 0 $X=16420 $Y=19630
X2987 2 DigitalLDOLogic_VIA1 $T=16670 23940 0 0 $X=16420 $Y=23710
X2988 2 DigitalLDOLogic_VIA1 $T=16670 28020 0 0 $X=16420 $Y=27790
X2989 2 DigitalLDOLogic_VIA1 $T=16670 32100 0 0 $X=16420 $Y=31870
X2990 2 DigitalLDOLogic_VIA1 $T=16670 36180 0 0 $X=16420 $Y=35950
X2991 2 DigitalLDOLogic_VIA1 $T=16670 40260 0 0 $X=16420 $Y=40030
X2992 2 DigitalLDOLogic_VIA1 $T=16670 44340 0 0 $X=16420 $Y=44110
X2993 2 DigitalLDOLogic_VIA1 $T=16670 48420 0 0 $X=16420 $Y=48190
X2994 2 DigitalLDOLogic_VIA1 $T=16670 52500 0 0 $X=16420 $Y=52270
X2995 2 DigitalLDOLogic_VIA1 $T=16670 56580 0 0 $X=16420 $Y=56350
X2996 1 DigitalLDOLogic_VIA1 $T=17590 13060 0 0 $X=17340 $Y=12830
X2997 1 DigitalLDOLogic_VIA1 $T=17590 17140 0 0 $X=17340 $Y=16910
X2998 1 DigitalLDOLogic_VIA1 $T=17590 21220 0 0 $X=17340 $Y=20990
X2999 1 DigitalLDOLogic_VIA1 $T=17590 25300 0 0 $X=17340 $Y=25070
X3000 1 DigitalLDOLogic_VIA1 $T=17590 29380 0 0 $X=17340 $Y=29150
X3001 1 DigitalLDOLogic_VIA1 $T=17590 33460 0 0 $X=17340 $Y=33230
X3002 1 DigitalLDOLogic_VIA1 $T=17590 37540 0 0 $X=17340 $Y=37310
X3003 1 DigitalLDOLogic_VIA1 $T=17590 41620 0 0 $X=17340 $Y=41390
X3004 1 DigitalLDOLogic_VIA1 $T=17590 45700 0 0 $X=17340 $Y=45470
X3005 1 DigitalLDOLogic_VIA1 $T=17590 49780 0 0 $X=17340 $Y=49550
X3006 1 DigitalLDOLogic_VIA1 $T=17590 53860 0 0 $X=17340 $Y=53630
X3007 1 DigitalLDOLogic_VIA1 $T=17590 57940 0 0 $X=17340 $Y=57710
X3008 2 DigitalLDOLogic_VIA1 $T=19430 11700 0 0 $X=19180 $Y=11470
X3009 2 DigitalLDOLogic_VIA1 $T=19430 15780 0 0 $X=19180 $Y=15550
X3010 2 DigitalLDOLogic_VIA1 $T=19430 19860 0 0 $X=19180 $Y=19630
X3011 2 DigitalLDOLogic_VIA1 $T=19430 23940 0 0 $X=19180 $Y=23710
X3012 2 DigitalLDOLogic_VIA1 $T=19430 28020 0 0 $X=19180 $Y=27790
X3013 2 DigitalLDOLogic_VIA1 $T=19430 32100 0 0 $X=19180 $Y=31870
X3014 2 DigitalLDOLogic_VIA1 $T=19430 36180 0 0 $X=19180 $Y=35950
X3015 2 DigitalLDOLogic_VIA1 $T=19430 40260 0 0 $X=19180 $Y=40030
X3016 2 DigitalLDOLogic_VIA1 $T=19430 44340 0 0 $X=19180 $Y=44110
X3017 2 DigitalLDOLogic_VIA1 $T=19430 48420 0 0 $X=19180 $Y=48190
X3018 2 DigitalLDOLogic_VIA1 $T=19430 52500 0 0 $X=19180 $Y=52270
X3019 2 DigitalLDOLogic_VIA1 $T=19430 56580 0 0 $X=19180 $Y=56350
X3020 1 DigitalLDOLogic_VIA1 $T=20350 13060 0 0 $X=20100 $Y=12830
X3021 1 DigitalLDOLogic_VIA1 $T=20350 17140 0 0 $X=20100 $Y=16910
X3022 1 DigitalLDOLogic_VIA1 $T=20350 21220 0 0 $X=20100 $Y=20990
X3023 1 DigitalLDOLogic_VIA1 $T=20350 25300 0 0 $X=20100 $Y=25070
X3024 1 DigitalLDOLogic_VIA1 $T=20350 29380 0 0 $X=20100 $Y=29150
X3025 1 DigitalLDOLogic_VIA1 $T=20350 33460 0 0 $X=20100 $Y=33230
X3026 1 DigitalLDOLogic_VIA1 $T=20350 37540 0 0 $X=20100 $Y=37310
X3027 1 DigitalLDOLogic_VIA1 $T=20350 41620 0 0 $X=20100 $Y=41390
X3028 1 DigitalLDOLogic_VIA1 $T=20350 45700 0 0 $X=20100 $Y=45470
X3029 1 DigitalLDOLogic_VIA1 $T=20350 49780 0 0 $X=20100 $Y=49550
X3030 1 DigitalLDOLogic_VIA1 $T=20350 53860 0 0 $X=20100 $Y=53630
X3031 1 DigitalLDOLogic_VIA1 $T=20350 57940 0 0 $X=20100 $Y=57710
X3032 2 DigitalLDOLogic_VIA1 $T=22190 11700 0 0 $X=21940 $Y=11470
X3033 2 DigitalLDOLogic_VIA1 $T=22190 15780 0 0 $X=21940 $Y=15550
X3034 2 DigitalLDOLogic_VIA1 $T=22190 19860 0 0 $X=21940 $Y=19630
X3035 2 DigitalLDOLogic_VIA1 $T=22190 23940 0 0 $X=21940 $Y=23710
X3036 2 DigitalLDOLogic_VIA1 $T=22190 28020 0 0 $X=21940 $Y=27790
X3037 2 DigitalLDOLogic_VIA1 $T=22190 32100 0 0 $X=21940 $Y=31870
X3038 2 DigitalLDOLogic_VIA1 $T=22190 36180 0 0 $X=21940 $Y=35950
X3039 2 DigitalLDOLogic_VIA1 $T=22190 40260 0 0 $X=21940 $Y=40030
X3040 2 DigitalLDOLogic_VIA1 $T=22190 44340 0 0 $X=21940 $Y=44110
X3041 2 DigitalLDOLogic_VIA1 $T=22190 48420 0 0 $X=21940 $Y=48190
X3042 2 DigitalLDOLogic_VIA1 $T=22190 52500 0 0 $X=21940 $Y=52270
X3043 2 DigitalLDOLogic_VIA1 $T=22190 56580 0 0 $X=21940 $Y=56350
X3044 1 DigitalLDOLogic_VIA1 $T=23110 13060 0 0 $X=22860 $Y=12830
X3045 1 DigitalLDOLogic_VIA1 $T=23110 17140 0 0 $X=22860 $Y=16910
X3046 1 DigitalLDOLogic_VIA1 $T=23110 21220 0 0 $X=22860 $Y=20990
X3047 1 DigitalLDOLogic_VIA1 $T=23110 25300 0 0 $X=22860 $Y=25070
X3048 1 DigitalLDOLogic_VIA1 $T=23110 29380 0 0 $X=22860 $Y=29150
X3049 1 DigitalLDOLogic_VIA1 $T=23110 33460 0 0 $X=22860 $Y=33230
X3050 1 DigitalLDOLogic_VIA1 $T=23110 37540 0 0 $X=22860 $Y=37310
X3051 1 DigitalLDOLogic_VIA1 $T=23110 41620 0 0 $X=22860 $Y=41390
X3052 1 DigitalLDOLogic_VIA1 $T=23110 45700 0 0 $X=22860 $Y=45470
X3053 1 DigitalLDOLogic_VIA1 $T=23110 49780 0 0 $X=22860 $Y=49550
X3054 1 DigitalLDOLogic_VIA1 $T=23110 53860 0 0 $X=22860 $Y=53630
X3055 1 DigitalLDOLogic_VIA1 $T=23110 57940 0 0 $X=22860 $Y=57710
X3056 2 DigitalLDOLogic_VIA1 $T=24950 11700 0 0 $X=24700 $Y=11470
X3057 2 DigitalLDOLogic_VIA1 $T=24950 15780 0 0 $X=24700 $Y=15550
X3058 2 DigitalLDOLogic_VIA1 $T=24950 19860 0 0 $X=24700 $Y=19630
X3059 2 DigitalLDOLogic_VIA1 $T=24950 23940 0 0 $X=24700 $Y=23710
X3060 2 DigitalLDOLogic_VIA1 $T=24950 28020 0 0 $X=24700 $Y=27790
X3061 2 DigitalLDOLogic_VIA1 $T=24950 32100 0 0 $X=24700 $Y=31870
X3062 2 DigitalLDOLogic_VIA1 $T=24950 36180 0 0 $X=24700 $Y=35950
X3063 2 DigitalLDOLogic_VIA1 $T=24950 40260 0 0 $X=24700 $Y=40030
X3064 2 DigitalLDOLogic_VIA1 $T=24950 44340 0 0 $X=24700 $Y=44110
X3065 2 DigitalLDOLogic_VIA1 $T=24950 48420 0 0 $X=24700 $Y=48190
X3066 2 DigitalLDOLogic_VIA1 $T=24950 52500 0 0 $X=24700 $Y=52270
X3067 2 DigitalLDOLogic_VIA1 $T=24950 56580 0 0 $X=24700 $Y=56350
X3068 1 DigitalLDOLogic_VIA1 $T=25870 13060 0 0 $X=25620 $Y=12830
X3069 1 DigitalLDOLogic_VIA1 $T=25870 17140 0 0 $X=25620 $Y=16910
X3070 1 DigitalLDOLogic_VIA1 $T=25870 21220 0 0 $X=25620 $Y=20990
X3071 1 DigitalLDOLogic_VIA1 $T=25870 25300 0 0 $X=25620 $Y=25070
X3072 1 DigitalLDOLogic_VIA1 $T=25870 29380 0 0 $X=25620 $Y=29150
X3073 1 DigitalLDOLogic_VIA1 $T=25870 33460 0 0 $X=25620 $Y=33230
X3074 1 DigitalLDOLogic_VIA1 $T=25870 37540 0 0 $X=25620 $Y=37310
X3075 1 DigitalLDOLogic_VIA1 $T=25870 41620 0 0 $X=25620 $Y=41390
X3076 1 DigitalLDOLogic_VIA1 $T=25870 45700 0 0 $X=25620 $Y=45470
X3077 1 DigitalLDOLogic_VIA1 $T=25870 49780 0 0 $X=25620 $Y=49550
X3078 1 DigitalLDOLogic_VIA1 $T=25870 53860 0 0 $X=25620 $Y=53630
X3079 1 DigitalLDOLogic_VIA1 $T=25870 57940 0 0 $X=25620 $Y=57710
X3080 2 DigitalLDOLogic_VIA1 $T=27710 11700 0 0 $X=27460 $Y=11470
X3081 2 DigitalLDOLogic_VIA1 $T=27710 15780 0 0 $X=27460 $Y=15550
X3082 2 DigitalLDOLogic_VIA1 $T=27710 19860 0 0 $X=27460 $Y=19630
X3083 2 DigitalLDOLogic_VIA1 $T=27710 23940 0 0 $X=27460 $Y=23710
X3084 2 DigitalLDOLogic_VIA1 $T=27710 28020 0 0 $X=27460 $Y=27790
X3085 2 DigitalLDOLogic_VIA1 $T=27710 32100 0 0 $X=27460 $Y=31870
X3086 2 DigitalLDOLogic_VIA1 $T=27710 36180 0 0 $X=27460 $Y=35950
X3087 2 DigitalLDOLogic_VIA1 $T=27710 40260 0 0 $X=27460 $Y=40030
X3088 2 DigitalLDOLogic_VIA1 $T=27710 44340 0 0 $X=27460 $Y=44110
X3089 2 DigitalLDOLogic_VIA1 $T=27710 48420 0 0 $X=27460 $Y=48190
X3090 2 DigitalLDOLogic_VIA1 $T=27710 52500 0 0 $X=27460 $Y=52270
X3091 2 DigitalLDOLogic_VIA1 $T=27710 56580 0 0 $X=27460 $Y=56350
X3092 1 DigitalLDOLogic_VIA1 $T=28630 13060 0 0 $X=28380 $Y=12830
X3093 1 DigitalLDOLogic_VIA1 $T=28630 17140 0 0 $X=28380 $Y=16910
X3094 1 DigitalLDOLogic_VIA1 $T=28630 21220 0 0 $X=28380 $Y=20990
X3095 1 DigitalLDOLogic_VIA1 $T=28630 25300 0 0 $X=28380 $Y=25070
X3096 1 DigitalLDOLogic_VIA1 $T=28630 29380 0 0 $X=28380 $Y=29150
X3097 1 DigitalLDOLogic_VIA1 $T=28630 33460 0 0 $X=28380 $Y=33230
X3098 1 DigitalLDOLogic_VIA1 $T=28630 37540 0 0 $X=28380 $Y=37310
X3099 1 DigitalLDOLogic_VIA1 $T=28630 41620 0 0 $X=28380 $Y=41390
X3100 1 DigitalLDOLogic_VIA1 $T=28630 45700 0 0 $X=28380 $Y=45470
X3101 1 DigitalLDOLogic_VIA1 $T=28630 49780 0 0 $X=28380 $Y=49550
X3102 1 DigitalLDOLogic_VIA1 $T=28630 53860 0 0 $X=28380 $Y=53630
X3103 1 DigitalLDOLogic_VIA1 $T=28630 57940 0 0 $X=28380 $Y=57710
X3104 2 DigitalLDOLogic_VIA1 $T=30470 11700 0 0 $X=30220 $Y=11470
X3105 2 DigitalLDOLogic_VIA1 $T=30470 15780 0 0 $X=30220 $Y=15550
X3106 2 DigitalLDOLogic_VIA1 $T=30470 19860 0 0 $X=30220 $Y=19630
X3107 2 DigitalLDOLogic_VIA1 $T=30470 23940 0 0 $X=30220 $Y=23710
X3108 2 DigitalLDOLogic_VIA1 $T=30470 28020 0 0 $X=30220 $Y=27790
X3109 2 DigitalLDOLogic_VIA1 $T=30470 32100 0 0 $X=30220 $Y=31870
X3110 2 DigitalLDOLogic_VIA1 $T=30470 36180 0 0 $X=30220 $Y=35950
X3111 2 DigitalLDOLogic_VIA1 $T=30470 40260 0 0 $X=30220 $Y=40030
X3112 2 DigitalLDOLogic_VIA1 $T=30470 44340 0 0 $X=30220 $Y=44110
X3113 2 DigitalLDOLogic_VIA1 $T=30470 48420 0 0 $X=30220 $Y=48190
X3114 2 DigitalLDOLogic_VIA1 $T=30470 52500 0 0 $X=30220 $Y=52270
X3115 2 DigitalLDOLogic_VIA1 $T=30470 56580 0 0 $X=30220 $Y=56350
X3116 1 DigitalLDOLogic_VIA1 $T=31390 13060 0 0 $X=31140 $Y=12830
X3117 1 DigitalLDOLogic_VIA1 $T=31390 17140 0 0 $X=31140 $Y=16910
X3118 1 DigitalLDOLogic_VIA1 $T=31390 21220 0 0 $X=31140 $Y=20990
X3119 1 DigitalLDOLogic_VIA1 $T=31390 25300 0 0 $X=31140 $Y=25070
X3120 1 DigitalLDOLogic_VIA1 $T=31390 29380 0 0 $X=31140 $Y=29150
X3121 1 DigitalLDOLogic_VIA1 $T=31390 33460 0 0 $X=31140 $Y=33230
X3122 1 DigitalLDOLogic_VIA1 $T=31390 37540 0 0 $X=31140 $Y=37310
X3123 1 DigitalLDOLogic_VIA1 $T=31390 41620 0 0 $X=31140 $Y=41390
X3124 1 DigitalLDOLogic_VIA1 $T=31390 45700 0 0 $X=31140 $Y=45470
X3125 1 DigitalLDOLogic_VIA1 $T=31390 49780 0 0 $X=31140 $Y=49550
X3126 1 DigitalLDOLogic_VIA1 $T=31390 53860 0 0 $X=31140 $Y=53630
X3127 1 DigitalLDOLogic_VIA1 $T=31390 57940 0 0 $X=31140 $Y=57710
X3128 2 DigitalLDOLogic_VIA1 $T=33230 11700 0 0 $X=32980 $Y=11470
X3129 2 DigitalLDOLogic_VIA1 $T=33230 15780 0 0 $X=32980 $Y=15550
X3130 2 DigitalLDOLogic_VIA1 $T=33230 19860 0 0 $X=32980 $Y=19630
X3131 2 DigitalLDOLogic_VIA1 $T=33230 23940 0 0 $X=32980 $Y=23710
X3132 2 DigitalLDOLogic_VIA1 $T=33230 28020 0 0 $X=32980 $Y=27790
X3133 2 DigitalLDOLogic_VIA1 $T=33230 32100 0 0 $X=32980 $Y=31870
X3134 2 DigitalLDOLogic_VIA1 $T=33230 36180 0 0 $X=32980 $Y=35950
X3135 2 DigitalLDOLogic_VIA1 $T=33230 40260 0 0 $X=32980 $Y=40030
X3136 2 DigitalLDOLogic_VIA1 $T=33230 44340 0 0 $X=32980 $Y=44110
X3137 2 DigitalLDOLogic_VIA1 $T=33230 48420 0 0 $X=32980 $Y=48190
X3138 2 DigitalLDOLogic_VIA1 $T=33230 52500 0 0 $X=32980 $Y=52270
X3139 2 DigitalLDOLogic_VIA1 $T=33230 56580 0 0 $X=32980 $Y=56350
X3140 1 DigitalLDOLogic_VIA1 $T=34150 13060 0 0 $X=33900 $Y=12830
X3141 1 DigitalLDOLogic_VIA1 $T=34150 17140 0 0 $X=33900 $Y=16910
X3142 1 DigitalLDOLogic_VIA1 $T=34150 21220 0 0 $X=33900 $Y=20990
X3143 1 DigitalLDOLogic_VIA1 $T=34150 25300 0 0 $X=33900 $Y=25070
X3144 1 DigitalLDOLogic_VIA1 $T=34150 29380 0 0 $X=33900 $Y=29150
X3145 1 DigitalLDOLogic_VIA1 $T=34150 33460 0 0 $X=33900 $Y=33230
X3146 1 DigitalLDOLogic_VIA1 $T=34150 37540 0 0 $X=33900 $Y=37310
X3147 1 DigitalLDOLogic_VIA1 $T=34150 41620 0 0 $X=33900 $Y=41390
X3148 1 DigitalLDOLogic_VIA1 $T=34150 45700 0 0 $X=33900 $Y=45470
X3149 1 DigitalLDOLogic_VIA1 $T=34150 49780 0 0 $X=33900 $Y=49550
X3150 1 DigitalLDOLogic_VIA1 $T=34150 53860 0 0 $X=33900 $Y=53630
X3151 1 DigitalLDOLogic_VIA1 $T=34150 57940 0 0 $X=33900 $Y=57710
X3152 2 DigitalLDOLogic_VIA1 $T=35990 11700 0 0 $X=35740 $Y=11470
X3153 2 DigitalLDOLogic_VIA1 $T=35990 15780 0 0 $X=35740 $Y=15550
X3154 2 DigitalLDOLogic_VIA1 $T=35990 19860 0 0 $X=35740 $Y=19630
X3155 2 DigitalLDOLogic_VIA1 $T=35990 23940 0 0 $X=35740 $Y=23710
X3156 2 DigitalLDOLogic_VIA1 $T=35990 28020 0 0 $X=35740 $Y=27790
X3157 2 DigitalLDOLogic_VIA1 $T=35990 32100 0 0 $X=35740 $Y=31870
X3158 2 DigitalLDOLogic_VIA1 $T=35990 36180 0 0 $X=35740 $Y=35950
X3159 2 DigitalLDOLogic_VIA1 $T=35990 40260 0 0 $X=35740 $Y=40030
X3160 2 DigitalLDOLogic_VIA1 $T=35990 44340 0 0 $X=35740 $Y=44110
X3161 2 DigitalLDOLogic_VIA1 $T=35990 48420 0 0 $X=35740 $Y=48190
X3162 2 DigitalLDOLogic_VIA1 $T=35990 52500 0 0 $X=35740 $Y=52270
X3163 2 DigitalLDOLogic_VIA1 $T=35990 56580 0 0 $X=35740 $Y=56350
X3164 1 DigitalLDOLogic_VIA1 $T=36910 13060 0 0 $X=36660 $Y=12830
X3165 1 DigitalLDOLogic_VIA1 $T=36910 17140 0 0 $X=36660 $Y=16910
X3166 1 DigitalLDOLogic_VIA1 $T=36910 21220 0 0 $X=36660 $Y=20990
X3167 1 DigitalLDOLogic_VIA1 $T=36910 25300 0 0 $X=36660 $Y=25070
X3168 1 DigitalLDOLogic_VIA1 $T=36910 29380 0 0 $X=36660 $Y=29150
X3169 1 DigitalLDOLogic_VIA1 $T=36910 33460 0 0 $X=36660 $Y=33230
X3170 1 DigitalLDOLogic_VIA1 $T=36910 37540 0 0 $X=36660 $Y=37310
X3171 1 DigitalLDOLogic_VIA1 $T=36910 41620 0 0 $X=36660 $Y=41390
X3172 1 DigitalLDOLogic_VIA1 $T=36910 45700 0 0 $X=36660 $Y=45470
X3173 1 DigitalLDOLogic_VIA1 $T=36910 49780 0 0 $X=36660 $Y=49550
X3174 1 DigitalLDOLogic_VIA1 $T=36910 53860 0 0 $X=36660 $Y=53630
X3175 1 DigitalLDOLogic_VIA1 $T=36910 57940 0 0 $X=36660 $Y=57710
X3176 2 DigitalLDOLogic_VIA1 $T=38750 11700 0 0 $X=38500 $Y=11470
X3177 2 DigitalLDOLogic_VIA1 $T=38750 15780 0 0 $X=38500 $Y=15550
X3178 2 DigitalLDOLogic_VIA1 $T=38750 19860 0 0 $X=38500 $Y=19630
X3179 2 DigitalLDOLogic_VIA1 $T=38750 23940 0 0 $X=38500 $Y=23710
X3180 2 DigitalLDOLogic_VIA1 $T=38750 28020 0 0 $X=38500 $Y=27790
X3181 2 DigitalLDOLogic_VIA1 $T=38750 32100 0 0 $X=38500 $Y=31870
X3182 2 DigitalLDOLogic_VIA1 $T=38750 36180 0 0 $X=38500 $Y=35950
X3183 2 DigitalLDOLogic_VIA1 $T=38750 40260 0 0 $X=38500 $Y=40030
X3184 2 DigitalLDOLogic_VIA1 $T=38750 44340 0 0 $X=38500 $Y=44110
X3185 2 DigitalLDOLogic_VIA1 $T=38750 48420 0 0 $X=38500 $Y=48190
X3186 2 DigitalLDOLogic_VIA1 $T=38750 52500 0 0 $X=38500 $Y=52270
X3187 2 DigitalLDOLogic_VIA1 $T=38750 56580 0 0 $X=38500 $Y=56350
X3188 1 DigitalLDOLogic_VIA1 $T=39670 13060 0 0 $X=39420 $Y=12830
X3189 1 DigitalLDOLogic_VIA1 $T=39670 17140 0 0 $X=39420 $Y=16910
X3190 1 DigitalLDOLogic_VIA1 $T=39670 21220 0 0 $X=39420 $Y=20990
X3191 1 DigitalLDOLogic_VIA1 $T=39670 25300 0 0 $X=39420 $Y=25070
X3192 1 DigitalLDOLogic_VIA1 $T=39670 29380 0 0 $X=39420 $Y=29150
X3193 1 DigitalLDOLogic_VIA1 $T=39670 33460 0 0 $X=39420 $Y=33230
X3194 1 DigitalLDOLogic_VIA1 $T=39670 37540 0 0 $X=39420 $Y=37310
X3195 1 DigitalLDOLogic_VIA1 $T=39670 41620 0 0 $X=39420 $Y=41390
X3196 1 DigitalLDOLogic_VIA1 $T=39670 45700 0 0 $X=39420 $Y=45470
X3197 1 DigitalLDOLogic_VIA1 $T=39670 49780 0 0 $X=39420 $Y=49550
X3198 1 DigitalLDOLogic_VIA1 $T=39670 53860 0 0 $X=39420 $Y=53630
X3199 1 DigitalLDOLogic_VIA1 $T=39670 57940 0 0 $X=39420 $Y=57710
X3200 2 DigitalLDOLogic_VIA1 $T=41510 11700 0 0 $X=41260 $Y=11470
X3201 2 DigitalLDOLogic_VIA1 $T=41510 15780 0 0 $X=41260 $Y=15550
X3202 2 DigitalLDOLogic_VIA1 $T=41510 19860 0 0 $X=41260 $Y=19630
X3203 2 DigitalLDOLogic_VIA1 $T=41510 23940 0 0 $X=41260 $Y=23710
X3204 2 DigitalLDOLogic_VIA1 $T=41510 28020 0 0 $X=41260 $Y=27790
X3205 2 DigitalLDOLogic_VIA1 $T=41510 32100 0 0 $X=41260 $Y=31870
X3206 2 DigitalLDOLogic_VIA1 $T=41510 36180 0 0 $X=41260 $Y=35950
X3207 2 DigitalLDOLogic_VIA1 $T=41510 40260 0 0 $X=41260 $Y=40030
X3208 2 DigitalLDOLogic_VIA1 $T=41510 44340 0 0 $X=41260 $Y=44110
X3209 2 DigitalLDOLogic_VIA1 $T=41510 48420 0 0 $X=41260 $Y=48190
X3210 2 DigitalLDOLogic_VIA1 $T=41510 52500 0 0 $X=41260 $Y=52270
X3211 2 DigitalLDOLogic_VIA1 $T=41510 56580 0 0 $X=41260 $Y=56350
X3212 1 DigitalLDOLogic_VIA1 $T=42430 13060 0 0 $X=42180 $Y=12830
X3213 1 DigitalLDOLogic_VIA1 $T=42430 17140 0 0 $X=42180 $Y=16910
X3214 1 DigitalLDOLogic_VIA1 $T=42430 21220 0 0 $X=42180 $Y=20990
X3215 1 DigitalLDOLogic_VIA1 $T=42430 25300 0 0 $X=42180 $Y=25070
X3216 1 DigitalLDOLogic_VIA1 $T=42430 29380 0 0 $X=42180 $Y=29150
X3217 1 DigitalLDOLogic_VIA1 $T=42430 33460 0 0 $X=42180 $Y=33230
X3218 1 DigitalLDOLogic_VIA1 $T=42430 37540 0 0 $X=42180 $Y=37310
X3219 1 DigitalLDOLogic_VIA1 $T=42430 41620 0 0 $X=42180 $Y=41390
X3220 1 DigitalLDOLogic_VIA1 $T=42430 45700 0 0 $X=42180 $Y=45470
X3221 1 DigitalLDOLogic_VIA1 $T=42430 49780 0 0 $X=42180 $Y=49550
X3222 1 DigitalLDOLogic_VIA1 $T=42430 53860 0 0 $X=42180 $Y=53630
X3223 1 DigitalLDOLogic_VIA1 $T=42430 57940 0 0 $X=42180 $Y=57710
X3224 2 DigitalLDOLogic_VIA1 $T=44270 11700 0 0 $X=44020 $Y=11470
X3225 2 DigitalLDOLogic_VIA1 $T=44270 15780 0 0 $X=44020 $Y=15550
X3226 2 DigitalLDOLogic_VIA1 $T=44270 19860 0 0 $X=44020 $Y=19630
X3227 2 DigitalLDOLogic_VIA1 $T=44270 23940 0 0 $X=44020 $Y=23710
X3228 2 DigitalLDOLogic_VIA1 $T=44270 28020 0 0 $X=44020 $Y=27790
X3229 2 DigitalLDOLogic_VIA1 $T=44270 32100 0 0 $X=44020 $Y=31870
X3230 2 DigitalLDOLogic_VIA1 $T=44270 36180 0 0 $X=44020 $Y=35950
X3231 2 DigitalLDOLogic_VIA1 $T=44270 40260 0 0 $X=44020 $Y=40030
X3232 2 DigitalLDOLogic_VIA1 $T=44270 44340 0 0 $X=44020 $Y=44110
X3233 2 DigitalLDOLogic_VIA1 $T=44270 48420 0 0 $X=44020 $Y=48190
X3234 2 DigitalLDOLogic_VIA1 $T=44270 52500 0 0 $X=44020 $Y=52270
X3235 2 DigitalLDOLogic_VIA1 $T=44270 56580 0 0 $X=44020 $Y=56350
X3236 1 DigitalLDOLogic_VIA1 $T=45190 13060 0 0 $X=44940 $Y=12830
X3237 1 DigitalLDOLogic_VIA1 $T=45190 17140 0 0 $X=44940 $Y=16910
X3238 1 DigitalLDOLogic_VIA1 $T=45190 21220 0 0 $X=44940 $Y=20990
X3239 1 DigitalLDOLogic_VIA1 $T=45190 25300 0 0 $X=44940 $Y=25070
X3240 1 DigitalLDOLogic_VIA1 $T=45190 29380 0 0 $X=44940 $Y=29150
X3241 1 DigitalLDOLogic_VIA1 $T=45190 33460 0 0 $X=44940 $Y=33230
X3242 1 DigitalLDOLogic_VIA1 $T=45190 37540 0 0 $X=44940 $Y=37310
X3243 1 DigitalLDOLogic_VIA1 $T=45190 41620 0 0 $X=44940 $Y=41390
X3244 1 DigitalLDOLogic_VIA1 $T=45190 45700 0 0 $X=44940 $Y=45470
X3245 1 DigitalLDOLogic_VIA1 $T=45190 49780 0 0 $X=44940 $Y=49550
X3246 1 DigitalLDOLogic_VIA1 $T=45190 53860 0 0 $X=44940 $Y=53630
X3247 1 DigitalLDOLogic_VIA1 $T=45190 57940 0 0 $X=44940 $Y=57710
X3248 2 DigitalLDOLogic_VIA1 $T=47030 11700 0 0 $X=46780 $Y=11470
X3249 2 DigitalLDOLogic_VIA1 $T=47030 15780 0 0 $X=46780 $Y=15550
X3250 2 DigitalLDOLogic_VIA1 $T=47030 19860 0 0 $X=46780 $Y=19630
X3251 2 DigitalLDOLogic_VIA1 $T=47030 23940 0 0 $X=46780 $Y=23710
X3252 2 DigitalLDOLogic_VIA1 $T=47030 28020 0 0 $X=46780 $Y=27790
X3253 2 DigitalLDOLogic_VIA1 $T=47030 32100 0 0 $X=46780 $Y=31870
X3254 2 DigitalLDOLogic_VIA1 $T=47030 36180 0 0 $X=46780 $Y=35950
X3255 2 DigitalLDOLogic_VIA1 $T=47030 40260 0 0 $X=46780 $Y=40030
X3256 2 DigitalLDOLogic_VIA1 $T=47030 44340 0 0 $X=46780 $Y=44110
X3257 2 DigitalLDOLogic_VIA1 $T=47030 48420 0 0 $X=46780 $Y=48190
X3258 2 DigitalLDOLogic_VIA1 $T=47030 52500 0 0 $X=46780 $Y=52270
X3259 2 DigitalLDOLogic_VIA1 $T=47030 56580 0 0 $X=46780 $Y=56350
X3260 1 DigitalLDOLogic_VIA1 $T=47950 13060 0 0 $X=47700 $Y=12830
X3261 1 DigitalLDOLogic_VIA1 $T=47950 17140 0 0 $X=47700 $Y=16910
X3262 1 DigitalLDOLogic_VIA1 $T=47950 21220 0 0 $X=47700 $Y=20990
X3263 1 DigitalLDOLogic_VIA1 $T=47950 25300 0 0 $X=47700 $Y=25070
X3264 1 DigitalLDOLogic_VIA1 $T=47950 29380 0 0 $X=47700 $Y=29150
X3265 1 DigitalLDOLogic_VIA1 $T=47950 33460 0 0 $X=47700 $Y=33230
X3266 1 DigitalLDOLogic_VIA1 $T=47950 37540 0 0 $X=47700 $Y=37310
X3267 1 DigitalLDOLogic_VIA1 $T=47950 41620 0 0 $X=47700 $Y=41390
X3268 1 DigitalLDOLogic_VIA1 $T=47950 45700 0 0 $X=47700 $Y=45470
X3269 1 DigitalLDOLogic_VIA1 $T=47950 49780 0 0 $X=47700 $Y=49550
X3270 1 DigitalLDOLogic_VIA1 $T=47950 53860 0 0 $X=47700 $Y=53630
X3271 1 DigitalLDOLogic_VIA1 $T=47950 57940 0 0 $X=47700 $Y=57710
X3272 2 DigitalLDOLogic_VIA1 $T=49790 11700 0 0 $X=49540 $Y=11470
X3273 2 DigitalLDOLogic_VIA1 $T=49790 15780 0 0 $X=49540 $Y=15550
X3274 2 DigitalLDOLogic_VIA1 $T=49790 19860 0 0 $X=49540 $Y=19630
X3275 2 DigitalLDOLogic_VIA1 $T=49790 23940 0 0 $X=49540 $Y=23710
X3276 2 DigitalLDOLogic_VIA1 $T=49790 28020 0 0 $X=49540 $Y=27790
X3277 2 DigitalLDOLogic_VIA1 $T=49790 32100 0 0 $X=49540 $Y=31870
X3278 2 DigitalLDOLogic_VIA1 $T=49790 36180 0 0 $X=49540 $Y=35950
X3279 2 DigitalLDOLogic_VIA1 $T=49790 40260 0 0 $X=49540 $Y=40030
X3280 2 DigitalLDOLogic_VIA1 $T=49790 44340 0 0 $X=49540 $Y=44110
X3281 2 DigitalLDOLogic_VIA1 $T=49790 48420 0 0 $X=49540 $Y=48190
X3282 2 DigitalLDOLogic_VIA1 $T=49790 52500 0 0 $X=49540 $Y=52270
X3283 2 DigitalLDOLogic_VIA1 $T=49790 56580 0 0 $X=49540 $Y=56350
X3284 1 DigitalLDOLogic_VIA1 $T=50710 13060 0 0 $X=50460 $Y=12830
X3285 1 DigitalLDOLogic_VIA1 $T=50710 17140 0 0 $X=50460 $Y=16910
X3286 1 DigitalLDOLogic_VIA1 $T=50710 21220 0 0 $X=50460 $Y=20990
X3287 1 DigitalLDOLogic_VIA1 $T=50710 25300 0 0 $X=50460 $Y=25070
X3288 1 DigitalLDOLogic_VIA1 $T=50710 29380 0 0 $X=50460 $Y=29150
X3289 1 DigitalLDOLogic_VIA1 $T=50710 33460 0 0 $X=50460 $Y=33230
X3290 1 DigitalLDOLogic_VIA1 $T=50710 37540 0 0 $X=50460 $Y=37310
X3291 1 DigitalLDOLogic_VIA1 $T=50710 41620 0 0 $X=50460 $Y=41390
X3292 1 DigitalLDOLogic_VIA1 $T=50710 45700 0 0 $X=50460 $Y=45470
X3293 1 DigitalLDOLogic_VIA1 $T=50710 49780 0 0 $X=50460 $Y=49550
X3294 1 DigitalLDOLogic_VIA1 $T=50710 53860 0 0 $X=50460 $Y=53630
X3295 1 DigitalLDOLogic_VIA1 $T=50710 57940 0 0 $X=50460 $Y=57710
X3296 2 DigitalLDOLogic_VIA1 $T=52550 11700 0 0 $X=52300 $Y=11470
X3297 2 DigitalLDOLogic_VIA1 $T=52550 15780 0 0 $X=52300 $Y=15550
X3298 2 DigitalLDOLogic_VIA1 $T=52550 19860 0 0 $X=52300 $Y=19630
X3299 2 DigitalLDOLogic_VIA1 $T=52550 23940 0 0 $X=52300 $Y=23710
X3300 2 DigitalLDOLogic_VIA1 $T=52550 28020 0 0 $X=52300 $Y=27790
X3301 2 DigitalLDOLogic_VIA1 $T=52550 32100 0 0 $X=52300 $Y=31870
X3302 2 DigitalLDOLogic_VIA1 $T=52550 36180 0 0 $X=52300 $Y=35950
X3303 2 DigitalLDOLogic_VIA1 $T=52550 40260 0 0 $X=52300 $Y=40030
X3304 2 DigitalLDOLogic_VIA1 $T=52550 44340 0 0 $X=52300 $Y=44110
X3305 2 DigitalLDOLogic_VIA1 $T=52550 48420 0 0 $X=52300 $Y=48190
X3306 2 DigitalLDOLogic_VIA1 $T=52550 52500 0 0 $X=52300 $Y=52270
X3307 2 DigitalLDOLogic_VIA1 $T=52550 56580 0 0 $X=52300 $Y=56350
X3308 1 DigitalLDOLogic_VIA1 $T=53470 13060 0 0 $X=53220 $Y=12830
X3309 1 DigitalLDOLogic_VIA1 $T=53470 17140 0 0 $X=53220 $Y=16910
X3310 1 DigitalLDOLogic_VIA1 $T=53470 21220 0 0 $X=53220 $Y=20990
X3311 1 DigitalLDOLogic_VIA1 $T=53470 25300 0 0 $X=53220 $Y=25070
X3312 1 DigitalLDOLogic_VIA1 $T=53470 29380 0 0 $X=53220 $Y=29150
X3313 1 DigitalLDOLogic_VIA1 $T=53470 33460 0 0 $X=53220 $Y=33230
X3314 1 DigitalLDOLogic_VIA1 $T=53470 37540 0 0 $X=53220 $Y=37310
X3315 1 DigitalLDOLogic_VIA1 $T=53470 41620 0 0 $X=53220 $Y=41390
X3316 1 DigitalLDOLogic_VIA1 $T=53470 45700 0 0 $X=53220 $Y=45470
X3317 1 DigitalLDOLogic_VIA1 $T=53470 49780 0 0 $X=53220 $Y=49550
X3318 1 DigitalLDOLogic_VIA1 $T=53470 53860 0 0 $X=53220 $Y=53630
X3319 1 DigitalLDOLogic_VIA1 $T=53470 57940 0 0 $X=53220 $Y=57710
X3320 2 DigitalLDOLogic_VIA1 $T=55310 11700 0 0 $X=55060 $Y=11470
X3321 2 DigitalLDOLogic_VIA1 $T=55310 15780 0 0 $X=55060 $Y=15550
X3322 2 DigitalLDOLogic_VIA1 $T=55310 19860 0 0 $X=55060 $Y=19630
X3323 2 DigitalLDOLogic_VIA1 $T=55310 23940 0 0 $X=55060 $Y=23710
X3324 2 DigitalLDOLogic_VIA1 $T=55310 28020 0 0 $X=55060 $Y=27790
X3325 2 DigitalLDOLogic_VIA1 $T=55310 32100 0 0 $X=55060 $Y=31870
X3326 2 DigitalLDOLogic_VIA1 $T=55310 36180 0 0 $X=55060 $Y=35950
X3327 2 DigitalLDOLogic_VIA1 $T=55310 40260 0 0 $X=55060 $Y=40030
X3328 2 DigitalLDOLogic_VIA1 $T=55310 44340 0 0 $X=55060 $Y=44110
X3329 2 DigitalLDOLogic_VIA1 $T=55310 48420 0 0 $X=55060 $Y=48190
X3330 2 DigitalLDOLogic_VIA1 $T=55310 52500 0 0 $X=55060 $Y=52270
X3331 2 DigitalLDOLogic_VIA1 $T=55310 56580 0 0 $X=55060 $Y=56350
X3332 1 DigitalLDOLogic_VIA1 $T=56230 13060 0 0 $X=55980 $Y=12830
X3333 1 DigitalLDOLogic_VIA1 $T=56230 17140 0 0 $X=55980 $Y=16910
X3334 1 DigitalLDOLogic_VIA1 $T=56230 21220 0 0 $X=55980 $Y=20990
X3335 1 DigitalLDOLogic_VIA1 $T=56230 25300 0 0 $X=55980 $Y=25070
X3336 1 DigitalLDOLogic_VIA1 $T=56230 29380 0 0 $X=55980 $Y=29150
X3337 1 DigitalLDOLogic_VIA1 $T=56230 33460 0 0 $X=55980 $Y=33230
X3338 1 DigitalLDOLogic_VIA1 $T=56230 37540 0 0 $X=55980 $Y=37310
X3339 1 DigitalLDOLogic_VIA1 $T=56230 41620 0 0 $X=55980 $Y=41390
X3340 1 DigitalLDOLogic_VIA1 $T=56230 45700 0 0 $X=55980 $Y=45470
X3341 1 DigitalLDOLogic_VIA1 $T=56230 49780 0 0 $X=55980 $Y=49550
X3342 1 DigitalLDOLogic_VIA1 $T=56230 53860 0 0 $X=55980 $Y=53630
X3343 1 DigitalLDOLogic_VIA1 $T=56230 57940 0 0 $X=55980 $Y=57710
X3344 2 DigitalLDOLogic_VIA1 $T=58070 11700 0 0 $X=57820 $Y=11470
X3345 2 DigitalLDOLogic_VIA1 $T=58070 15780 0 0 $X=57820 $Y=15550
X3346 2 DigitalLDOLogic_VIA1 $T=58070 19860 0 0 $X=57820 $Y=19630
X3347 2 DigitalLDOLogic_VIA1 $T=58070 23940 0 0 $X=57820 $Y=23710
X3348 2 DigitalLDOLogic_VIA1 $T=58070 28020 0 0 $X=57820 $Y=27790
X3349 2 DigitalLDOLogic_VIA1 $T=58070 32100 0 0 $X=57820 $Y=31870
X3350 2 DigitalLDOLogic_VIA1 $T=58070 36180 0 0 $X=57820 $Y=35950
X3351 2 DigitalLDOLogic_VIA1 $T=58070 40260 0 0 $X=57820 $Y=40030
X3352 2 DigitalLDOLogic_VIA1 $T=58070 44340 0 0 $X=57820 $Y=44110
X3353 2 DigitalLDOLogic_VIA1 $T=58070 48420 0 0 $X=57820 $Y=48190
X3354 2 DigitalLDOLogic_VIA1 $T=58070 52500 0 0 $X=57820 $Y=52270
X3355 2 DigitalLDOLogic_VIA1 $T=58070 56580 0 0 $X=57820 $Y=56350
X3356 1 DigitalLDOLogic_VIA1 $T=58990 13060 0 0 $X=58740 $Y=12830
X3357 1 DigitalLDOLogic_VIA1 $T=58990 17140 0 0 $X=58740 $Y=16910
X3358 1 DigitalLDOLogic_VIA1 $T=58990 21220 0 0 $X=58740 $Y=20990
X3359 1 DigitalLDOLogic_VIA1 $T=58990 25300 0 0 $X=58740 $Y=25070
X3360 1 DigitalLDOLogic_VIA1 $T=58990 29380 0 0 $X=58740 $Y=29150
X3361 1 DigitalLDOLogic_VIA1 $T=58990 33460 0 0 $X=58740 $Y=33230
X3362 1 DigitalLDOLogic_VIA1 $T=58990 37540 0 0 $X=58740 $Y=37310
X3363 1 DigitalLDOLogic_VIA1 $T=58990 41620 0 0 $X=58740 $Y=41390
X3364 1 DigitalLDOLogic_VIA1 $T=58990 45700 0 0 $X=58740 $Y=45470
X3365 1 DigitalLDOLogic_VIA1 $T=58990 49780 0 0 $X=58740 $Y=49550
X3366 1 DigitalLDOLogic_VIA1 $T=58990 53860 0 0 $X=58740 $Y=53630
X3367 1 DigitalLDOLogic_VIA1 $T=58990 57940 0 0 $X=58740 $Y=57710
X3368 2 DigitalLDOLogic_VIA1 $T=60830 11700 0 0 $X=60580 $Y=11470
X3369 2 DigitalLDOLogic_VIA1 $T=60830 15780 0 0 $X=60580 $Y=15550
X3370 2 DigitalLDOLogic_VIA1 $T=60830 19860 0 0 $X=60580 $Y=19630
X3371 2 DigitalLDOLogic_VIA1 $T=60830 23940 0 0 $X=60580 $Y=23710
X3372 2 DigitalLDOLogic_VIA1 $T=60830 28020 0 0 $X=60580 $Y=27790
X3373 2 DigitalLDOLogic_VIA1 $T=60830 32100 0 0 $X=60580 $Y=31870
X3374 2 DigitalLDOLogic_VIA1 $T=60830 36180 0 0 $X=60580 $Y=35950
X3375 2 DigitalLDOLogic_VIA1 $T=60830 40260 0 0 $X=60580 $Y=40030
X3376 2 DigitalLDOLogic_VIA1 $T=60830 44340 0 0 $X=60580 $Y=44110
X3377 2 DigitalLDOLogic_VIA1 $T=60830 48420 0 0 $X=60580 $Y=48190
X3378 2 DigitalLDOLogic_VIA1 $T=60830 52500 0 0 $X=60580 $Y=52270
X3379 2 DigitalLDOLogic_VIA1 $T=60830 56580 0 0 $X=60580 $Y=56350
X3380 1 DigitalLDOLogic_VIA1 $T=61750 13060 0 0 $X=61500 $Y=12830
X3381 1 DigitalLDOLogic_VIA1 $T=61750 17140 0 0 $X=61500 $Y=16910
X3382 1 DigitalLDOLogic_VIA1 $T=61750 21220 0 0 $X=61500 $Y=20990
X3383 1 DigitalLDOLogic_VIA1 $T=61750 25300 0 0 $X=61500 $Y=25070
X3384 1 DigitalLDOLogic_VIA1 $T=61750 29380 0 0 $X=61500 $Y=29150
X3385 1 DigitalLDOLogic_VIA1 $T=61750 33460 0 0 $X=61500 $Y=33230
X3386 1 DigitalLDOLogic_VIA1 $T=61750 37540 0 0 $X=61500 $Y=37310
X3387 1 DigitalLDOLogic_VIA1 $T=61750 41620 0 0 $X=61500 $Y=41390
X3388 1 DigitalLDOLogic_VIA1 $T=61750 45700 0 0 $X=61500 $Y=45470
X3389 1 DigitalLDOLogic_VIA1 $T=61750 49780 0 0 $X=61500 $Y=49550
X3390 1 DigitalLDOLogic_VIA1 $T=61750 53860 0 0 $X=61500 $Y=53630
X3391 1 DigitalLDOLogic_VIA1 $T=61750 57940 0 0 $X=61500 $Y=57710
X3392 2 DigitalLDOLogic_VIA1 $T=63590 11700 0 0 $X=63340 $Y=11470
X3393 2 DigitalLDOLogic_VIA1 $T=63590 15780 0 0 $X=63340 $Y=15550
X3394 2 DigitalLDOLogic_VIA1 $T=63590 19860 0 0 $X=63340 $Y=19630
X3395 2 DigitalLDOLogic_VIA1 $T=63590 23940 0 0 $X=63340 $Y=23710
X3396 2 DigitalLDOLogic_VIA1 $T=63590 28020 0 0 $X=63340 $Y=27790
X3397 2 DigitalLDOLogic_VIA1 $T=63590 32100 0 0 $X=63340 $Y=31870
X3398 2 DigitalLDOLogic_VIA1 $T=63590 36180 0 0 $X=63340 $Y=35950
X3399 2 DigitalLDOLogic_VIA1 $T=63590 40260 0 0 $X=63340 $Y=40030
X3400 2 DigitalLDOLogic_VIA1 $T=63590 44340 0 0 $X=63340 $Y=44110
X3401 2 DigitalLDOLogic_VIA1 $T=63590 48420 0 0 $X=63340 $Y=48190
X3402 2 DigitalLDOLogic_VIA1 $T=63590 52500 0 0 $X=63340 $Y=52270
X3403 2 DigitalLDOLogic_VIA1 $T=63590 56580 0 0 $X=63340 $Y=56350
X3404 1 DigitalLDOLogic_VIA1 $T=64510 13060 0 0 $X=64260 $Y=12830
X3405 1 DigitalLDOLogic_VIA1 $T=64510 17140 0 0 $X=64260 $Y=16910
X3406 1 DigitalLDOLogic_VIA1 $T=64510 21220 0 0 $X=64260 $Y=20990
X3407 1 DigitalLDOLogic_VIA1 $T=64510 25300 0 0 $X=64260 $Y=25070
X3408 1 DigitalLDOLogic_VIA1 $T=64510 29380 0 0 $X=64260 $Y=29150
X3409 1 DigitalLDOLogic_VIA1 $T=64510 33460 0 0 $X=64260 $Y=33230
X3410 1 DigitalLDOLogic_VIA1 $T=64510 37540 0 0 $X=64260 $Y=37310
X3411 1 DigitalLDOLogic_VIA1 $T=64510 41620 0 0 $X=64260 $Y=41390
X3412 1 DigitalLDOLogic_VIA1 $T=64510 45700 0 0 $X=64260 $Y=45470
X3413 1 DigitalLDOLogic_VIA1 $T=64510 49780 0 0 $X=64260 $Y=49550
X3414 1 DigitalLDOLogic_VIA1 $T=64510 53860 0 0 $X=64260 $Y=53630
X3415 1 DigitalLDOLogic_VIA1 $T=64510 57940 0 0 $X=64260 $Y=57710
X3416 2 DigitalLDOLogic_VIA1 $T=66350 11700 0 0 $X=66100 $Y=11470
X3417 2 DigitalLDOLogic_VIA1 $T=66350 15780 0 0 $X=66100 $Y=15550
X3418 2 DigitalLDOLogic_VIA1 $T=66350 19860 0 0 $X=66100 $Y=19630
X3419 2 DigitalLDOLogic_VIA1 $T=66350 23940 0 0 $X=66100 $Y=23710
X3420 2 DigitalLDOLogic_VIA1 $T=66350 28020 0 0 $X=66100 $Y=27790
X3421 2 DigitalLDOLogic_VIA1 $T=66350 32100 0 0 $X=66100 $Y=31870
X3422 2 DigitalLDOLogic_VIA1 $T=66350 36180 0 0 $X=66100 $Y=35950
X3423 2 DigitalLDOLogic_VIA1 $T=66350 40260 0 0 $X=66100 $Y=40030
X3424 2 DigitalLDOLogic_VIA1 $T=66350 44340 0 0 $X=66100 $Y=44110
X3425 2 DigitalLDOLogic_VIA1 $T=66350 48420 0 0 $X=66100 $Y=48190
X3426 2 DigitalLDOLogic_VIA1 $T=66350 52500 0 0 $X=66100 $Y=52270
X3427 2 DigitalLDOLogic_VIA1 $T=66350 56580 0 0 $X=66100 $Y=56350
X3428 1 DigitalLDOLogic_VIA1 $T=67270 13060 0 0 $X=67020 $Y=12830
X3429 1 DigitalLDOLogic_VIA1 $T=67270 17140 0 0 $X=67020 $Y=16910
X3430 1 DigitalLDOLogic_VIA1 $T=67270 21220 0 0 $X=67020 $Y=20990
X3431 1 DigitalLDOLogic_VIA1 $T=67270 25300 0 0 $X=67020 $Y=25070
X3432 1 DigitalLDOLogic_VIA1 $T=67270 29380 0 0 $X=67020 $Y=29150
X3433 1 DigitalLDOLogic_VIA1 $T=67270 33460 0 0 $X=67020 $Y=33230
X3434 1 DigitalLDOLogic_VIA1 $T=67270 37540 0 0 $X=67020 $Y=37310
X3435 1 DigitalLDOLogic_VIA1 $T=67270 41620 0 0 $X=67020 $Y=41390
X3436 1 DigitalLDOLogic_VIA1 $T=67270 45700 0 0 $X=67020 $Y=45470
X3437 1 DigitalLDOLogic_VIA1 $T=67270 49780 0 0 $X=67020 $Y=49550
X3438 1 DigitalLDOLogic_VIA1 $T=67270 53860 0 0 $X=67020 $Y=53630
X3439 1 DigitalLDOLogic_VIA1 $T=67270 57940 0 0 $X=67020 $Y=57710
X3440 2 DigitalLDOLogic_VIA1 $T=69110 11700 0 0 $X=68860 $Y=11470
X3441 2 DigitalLDOLogic_VIA1 $T=69110 15780 0 0 $X=68860 $Y=15550
X3442 2 DigitalLDOLogic_VIA1 $T=69110 19860 0 0 $X=68860 $Y=19630
X3443 2 DigitalLDOLogic_VIA1 $T=69110 23940 0 0 $X=68860 $Y=23710
X3444 2 DigitalLDOLogic_VIA1 $T=69110 28020 0 0 $X=68860 $Y=27790
X3445 2 DigitalLDOLogic_VIA1 $T=69110 32100 0 0 $X=68860 $Y=31870
X3446 2 DigitalLDOLogic_VIA1 $T=69110 36180 0 0 $X=68860 $Y=35950
X3447 2 DigitalLDOLogic_VIA1 $T=69110 40260 0 0 $X=68860 $Y=40030
X3448 2 DigitalLDOLogic_VIA1 $T=69110 44340 0 0 $X=68860 $Y=44110
X3449 2 DigitalLDOLogic_VIA1 $T=69110 48420 0 0 $X=68860 $Y=48190
X3450 2 DigitalLDOLogic_VIA1 $T=69110 52500 0 0 $X=68860 $Y=52270
X3451 2 DigitalLDOLogic_VIA1 $T=69110 56580 0 0 $X=68860 $Y=56350
X3452 1 DigitalLDOLogic_VIA1 $T=70030 13060 0 0 $X=69780 $Y=12830
X3453 1 DigitalLDOLogic_VIA1 $T=70030 17140 0 0 $X=69780 $Y=16910
X3454 1 DigitalLDOLogic_VIA1 $T=70030 21220 0 0 $X=69780 $Y=20990
X3455 1 DigitalLDOLogic_VIA1 $T=70030 25300 0 0 $X=69780 $Y=25070
X3456 1 DigitalLDOLogic_VIA1 $T=70030 29380 0 0 $X=69780 $Y=29150
X3457 1 DigitalLDOLogic_VIA1 $T=70030 33460 0 0 $X=69780 $Y=33230
X3458 1 DigitalLDOLogic_VIA1 $T=70030 37540 0 0 $X=69780 $Y=37310
X3459 1 DigitalLDOLogic_VIA1 $T=70030 41620 0 0 $X=69780 $Y=41390
X3460 1 DigitalLDOLogic_VIA1 $T=70030 45700 0 0 $X=69780 $Y=45470
X3461 1 DigitalLDOLogic_VIA1 $T=70030 49780 0 0 $X=69780 $Y=49550
X3462 1 DigitalLDOLogic_VIA1 $T=70030 53860 0 0 $X=69780 $Y=53630
X3463 1 DigitalLDOLogic_VIA1 $T=70030 57940 0 0 $X=69780 $Y=57710
X3464 2 DigitalLDOLogic_VIA1 $T=71870 11700 0 0 $X=71620 $Y=11470
X3465 2 DigitalLDOLogic_VIA1 $T=71870 15780 0 0 $X=71620 $Y=15550
X3466 2 DigitalLDOLogic_VIA1 $T=71870 19860 0 0 $X=71620 $Y=19630
X3467 2 DigitalLDOLogic_VIA1 $T=71870 23940 0 0 $X=71620 $Y=23710
X3468 2 DigitalLDOLogic_VIA1 $T=71870 28020 0 0 $X=71620 $Y=27790
X3469 2 DigitalLDOLogic_VIA1 $T=71870 32100 0 0 $X=71620 $Y=31870
X3470 2 DigitalLDOLogic_VIA1 $T=71870 36180 0 0 $X=71620 $Y=35950
X3471 2 DigitalLDOLogic_VIA1 $T=71870 40260 0 0 $X=71620 $Y=40030
X3472 2 DigitalLDOLogic_VIA1 $T=71870 44340 0 0 $X=71620 $Y=44110
X3473 2 DigitalLDOLogic_VIA1 $T=71870 48420 0 0 $X=71620 $Y=48190
X3474 2 DigitalLDOLogic_VIA1 $T=71870 52500 0 0 $X=71620 $Y=52270
X3475 2 DigitalLDOLogic_VIA1 $T=71870 56580 0 0 $X=71620 $Y=56350
X3476 1 DigitalLDOLogic_VIA1 $T=72790 13060 0 0 $X=72540 $Y=12830
X3477 1 DigitalLDOLogic_VIA1 $T=72790 17140 0 0 $X=72540 $Y=16910
X3478 1 DigitalLDOLogic_VIA1 $T=72790 21220 0 0 $X=72540 $Y=20990
X3479 1 DigitalLDOLogic_VIA1 $T=72790 25300 0 0 $X=72540 $Y=25070
X3480 1 DigitalLDOLogic_VIA1 $T=72790 29380 0 0 $X=72540 $Y=29150
X3481 1 DigitalLDOLogic_VIA1 $T=72790 33460 0 0 $X=72540 $Y=33230
X3482 1 DigitalLDOLogic_VIA1 $T=72790 37540 0 0 $X=72540 $Y=37310
X3483 1 DigitalLDOLogic_VIA1 $T=72790 41620 0 0 $X=72540 $Y=41390
X3484 1 DigitalLDOLogic_VIA1 $T=72790 45700 0 0 $X=72540 $Y=45470
X3485 1 DigitalLDOLogic_VIA1 $T=72790 49780 0 0 $X=72540 $Y=49550
X3486 1 DigitalLDOLogic_VIA1 $T=72790 53860 0 0 $X=72540 $Y=53630
X3487 1 DigitalLDOLogic_VIA1 $T=72790 57940 0 0 $X=72540 $Y=57710
X3488 2 DigitalLDOLogic_VIA1 $T=74630 11700 0 0 $X=74380 $Y=11470
X3489 2 DigitalLDOLogic_VIA1 $T=74630 15780 0 0 $X=74380 $Y=15550
X3490 2 DigitalLDOLogic_VIA1 $T=74630 19860 0 0 $X=74380 $Y=19630
X3491 2 DigitalLDOLogic_VIA1 $T=74630 23940 0 0 $X=74380 $Y=23710
X3492 2 DigitalLDOLogic_VIA1 $T=74630 28020 0 0 $X=74380 $Y=27790
X3493 2 DigitalLDOLogic_VIA1 $T=74630 32100 0 0 $X=74380 $Y=31870
X3494 2 DigitalLDOLogic_VIA1 $T=74630 36180 0 0 $X=74380 $Y=35950
X3495 2 DigitalLDOLogic_VIA1 $T=74630 40260 0 0 $X=74380 $Y=40030
X3496 2 DigitalLDOLogic_VIA1 $T=74630 44340 0 0 $X=74380 $Y=44110
X3497 2 DigitalLDOLogic_VIA1 $T=74630 48420 0 0 $X=74380 $Y=48190
X3498 2 DigitalLDOLogic_VIA1 $T=74630 52500 0 0 $X=74380 $Y=52270
X3499 2 DigitalLDOLogic_VIA1 $T=74630 56580 0 0 $X=74380 $Y=56350
X3500 1 DigitalLDOLogic_VIA1 $T=75550 13060 0 0 $X=75300 $Y=12830
X3501 1 DigitalLDOLogic_VIA1 $T=75550 17140 0 0 $X=75300 $Y=16910
X3502 1 DigitalLDOLogic_VIA1 $T=75550 21220 0 0 $X=75300 $Y=20990
X3503 1 DigitalLDOLogic_VIA1 $T=75550 25300 0 0 $X=75300 $Y=25070
X3504 1 DigitalLDOLogic_VIA1 $T=75550 29380 0 0 $X=75300 $Y=29150
X3505 1 DigitalLDOLogic_VIA1 $T=75550 33460 0 0 $X=75300 $Y=33230
X3506 1 DigitalLDOLogic_VIA1 $T=75550 37540 0 0 $X=75300 $Y=37310
X3507 1 DigitalLDOLogic_VIA1 $T=75550 41620 0 0 $X=75300 $Y=41390
X3508 1 DigitalLDOLogic_VIA1 $T=75550 45700 0 0 $X=75300 $Y=45470
X3509 1 DigitalLDOLogic_VIA1 $T=75550 49780 0 0 $X=75300 $Y=49550
X3510 1 DigitalLDOLogic_VIA1 $T=75550 53860 0 0 $X=75300 $Y=53630
X3511 1 DigitalLDOLogic_VIA1 $T=75550 57940 0 0 $X=75300 $Y=57710
X3512 2 DigitalLDOLogic_VIA1 $T=77390 11700 0 0 $X=77140 $Y=11470
X3513 2 DigitalLDOLogic_VIA1 $T=77390 15780 0 0 $X=77140 $Y=15550
X3514 2 DigitalLDOLogic_VIA1 $T=77390 19860 0 0 $X=77140 $Y=19630
X3515 2 DigitalLDOLogic_VIA1 $T=77390 23940 0 0 $X=77140 $Y=23710
X3516 2 DigitalLDOLogic_VIA1 $T=77390 28020 0 0 $X=77140 $Y=27790
X3517 2 DigitalLDOLogic_VIA1 $T=77390 32100 0 0 $X=77140 $Y=31870
X3518 2 DigitalLDOLogic_VIA1 $T=77390 36180 0 0 $X=77140 $Y=35950
X3519 2 DigitalLDOLogic_VIA1 $T=77390 40260 0 0 $X=77140 $Y=40030
X3520 2 DigitalLDOLogic_VIA1 $T=77390 44340 0 0 $X=77140 $Y=44110
X3521 2 DigitalLDOLogic_VIA1 $T=77390 48420 0 0 $X=77140 $Y=48190
X3522 2 DigitalLDOLogic_VIA1 $T=77390 52500 0 0 $X=77140 $Y=52270
X3523 2 DigitalLDOLogic_VIA1 $T=77390 56580 0 0 $X=77140 $Y=56350
X3524 1 DigitalLDOLogic_VIA1 $T=78310 13060 0 0 $X=78060 $Y=12830
X3525 1 DigitalLDOLogic_VIA1 $T=78310 17140 0 0 $X=78060 $Y=16910
X3526 1 DigitalLDOLogic_VIA1 $T=78310 21220 0 0 $X=78060 $Y=20990
X3527 1 DigitalLDOLogic_VIA1 $T=78310 25300 0 0 $X=78060 $Y=25070
X3528 1 DigitalLDOLogic_VIA1 $T=78310 29380 0 0 $X=78060 $Y=29150
X3529 1 DigitalLDOLogic_VIA1 $T=78310 33460 0 0 $X=78060 $Y=33230
X3530 1 DigitalLDOLogic_VIA1 $T=78310 37540 0 0 $X=78060 $Y=37310
X3531 1 DigitalLDOLogic_VIA1 $T=78310 41620 0 0 $X=78060 $Y=41390
X3532 1 DigitalLDOLogic_VIA1 $T=78310 45700 0 0 $X=78060 $Y=45470
X3533 1 DigitalLDOLogic_VIA1 $T=78310 49780 0 0 $X=78060 $Y=49550
X3534 1 DigitalLDOLogic_VIA1 $T=78310 53860 0 0 $X=78060 $Y=53630
X3535 1 DigitalLDOLogic_VIA1 $T=78310 57940 0 0 $X=78060 $Y=57710
X3536 2 DigitalLDOLogic_VIA1 $T=80150 11700 0 0 $X=79900 $Y=11470
X3537 2 DigitalLDOLogic_VIA1 $T=80150 15780 0 0 $X=79900 $Y=15550
X3538 2 DigitalLDOLogic_VIA1 $T=80150 19860 0 0 $X=79900 $Y=19630
X3539 2 DigitalLDOLogic_VIA1 $T=80150 23940 0 0 $X=79900 $Y=23710
X3540 2 DigitalLDOLogic_VIA1 $T=80150 28020 0 0 $X=79900 $Y=27790
X3541 2 DigitalLDOLogic_VIA1 $T=80150 32100 0 0 $X=79900 $Y=31870
X3542 2 DigitalLDOLogic_VIA1 $T=80150 36180 0 0 $X=79900 $Y=35950
X3543 2 DigitalLDOLogic_VIA1 $T=80150 40260 0 0 $X=79900 $Y=40030
X3544 2 DigitalLDOLogic_VIA1 $T=80150 44340 0 0 $X=79900 $Y=44110
X3545 2 DigitalLDOLogic_VIA1 $T=80150 48420 0 0 $X=79900 $Y=48190
X3546 2 DigitalLDOLogic_VIA1 $T=80150 52500 0 0 $X=79900 $Y=52270
X3547 2 DigitalLDOLogic_VIA1 $T=80150 56580 0 0 $X=79900 $Y=56350
X3548 1 DigitalLDOLogic_VIA1 $T=81070 13060 0 0 $X=80820 $Y=12830
X3549 1 DigitalLDOLogic_VIA1 $T=81070 17140 0 0 $X=80820 $Y=16910
X3550 1 DigitalLDOLogic_VIA1 $T=81070 21220 0 0 $X=80820 $Y=20990
X3551 1 DigitalLDOLogic_VIA1 $T=81070 25300 0 0 $X=80820 $Y=25070
X3552 1 DigitalLDOLogic_VIA1 $T=81070 29380 0 0 $X=80820 $Y=29150
X3553 1 DigitalLDOLogic_VIA1 $T=81070 33460 0 0 $X=80820 $Y=33230
X3554 1 DigitalLDOLogic_VIA1 $T=81070 37540 0 0 $X=80820 $Y=37310
X3555 1 DigitalLDOLogic_VIA1 $T=81070 41620 0 0 $X=80820 $Y=41390
X3556 1 DigitalLDOLogic_VIA1 $T=81070 45700 0 0 $X=80820 $Y=45470
X3557 1 DigitalLDOLogic_VIA1 $T=81070 49780 0 0 $X=80820 $Y=49550
X3558 1 DigitalLDOLogic_VIA1 $T=81070 53860 0 0 $X=80820 $Y=53630
X3559 1 DigitalLDOLogic_VIA1 $T=81070 57940 0 0 $X=80820 $Y=57710
X3560 2 DigitalLDOLogic_VIA1 $T=82910 11700 0 0 $X=82660 $Y=11470
X3561 2 DigitalLDOLogic_VIA1 $T=82910 15780 0 0 $X=82660 $Y=15550
X3562 2 DigitalLDOLogic_VIA1 $T=82910 19860 0 0 $X=82660 $Y=19630
X3563 2 DigitalLDOLogic_VIA1 $T=82910 23940 0 0 $X=82660 $Y=23710
X3564 2 DigitalLDOLogic_VIA1 $T=82910 28020 0 0 $X=82660 $Y=27790
X3565 2 DigitalLDOLogic_VIA1 $T=82910 32100 0 0 $X=82660 $Y=31870
X3566 2 DigitalLDOLogic_VIA1 $T=82910 36180 0 0 $X=82660 $Y=35950
X3567 2 DigitalLDOLogic_VIA1 $T=82910 40260 0 0 $X=82660 $Y=40030
X3568 2 DigitalLDOLogic_VIA1 $T=82910 44340 0 0 $X=82660 $Y=44110
X3569 2 DigitalLDOLogic_VIA1 $T=82910 48420 0 0 $X=82660 $Y=48190
X3570 2 DigitalLDOLogic_VIA1 $T=82910 52500 0 0 $X=82660 $Y=52270
X3571 2 DigitalLDOLogic_VIA1 $T=82910 56580 0 0 $X=82660 $Y=56350
X3572 1 DigitalLDOLogic_VIA1 $T=83830 13060 0 0 $X=83580 $Y=12830
X3573 1 DigitalLDOLogic_VIA1 $T=83830 17140 0 0 $X=83580 $Y=16910
X3574 1 DigitalLDOLogic_VIA1 $T=83830 21220 0 0 $X=83580 $Y=20990
X3575 1 DigitalLDOLogic_VIA1 $T=83830 25300 0 0 $X=83580 $Y=25070
X3576 1 DigitalLDOLogic_VIA1 $T=83830 29380 0 0 $X=83580 $Y=29150
X3577 1 DigitalLDOLogic_VIA1 $T=83830 33460 0 0 $X=83580 $Y=33230
X3578 1 DigitalLDOLogic_VIA1 $T=83830 37540 0 0 $X=83580 $Y=37310
X3579 1 DigitalLDOLogic_VIA1 $T=83830 41620 0 0 $X=83580 $Y=41390
X3580 1 DigitalLDOLogic_VIA1 $T=83830 45700 0 0 $X=83580 $Y=45470
X3581 1 DigitalLDOLogic_VIA1 $T=83830 49780 0 0 $X=83580 $Y=49550
X3582 1 DigitalLDOLogic_VIA1 $T=83830 53860 0 0 $X=83580 $Y=53630
X3583 1 DigitalLDOLogic_VIA1 $T=83830 57940 0 0 $X=83580 $Y=57710
X3584 2 DigitalLDOLogic_VIA1 $T=85670 11700 0 0 $X=85420 $Y=11470
X3585 2 DigitalLDOLogic_VIA1 $T=85670 15780 0 0 $X=85420 $Y=15550
X3586 2 DigitalLDOLogic_VIA1 $T=85670 19860 0 0 $X=85420 $Y=19630
X3587 2 DigitalLDOLogic_VIA1 $T=85670 23940 0 0 $X=85420 $Y=23710
X3588 2 DigitalLDOLogic_VIA1 $T=85670 28020 0 0 $X=85420 $Y=27790
X3589 2 DigitalLDOLogic_VIA1 $T=85670 32100 0 0 $X=85420 $Y=31870
X3590 2 DigitalLDOLogic_VIA1 $T=85670 36180 0 0 $X=85420 $Y=35950
X3591 2 DigitalLDOLogic_VIA1 $T=85670 40260 0 0 $X=85420 $Y=40030
X3592 2 DigitalLDOLogic_VIA1 $T=85670 44340 0 0 $X=85420 $Y=44110
X3593 2 DigitalLDOLogic_VIA1 $T=85670 48420 0 0 $X=85420 $Y=48190
X3594 2 DigitalLDOLogic_VIA1 $T=85670 52500 0 0 $X=85420 $Y=52270
X3595 2 DigitalLDOLogic_VIA1 $T=85670 56580 0 0 $X=85420 $Y=56350
X3596 1 DigitalLDOLogic_VIA1 $T=86590 13060 0 0 $X=86340 $Y=12830
X3597 1 DigitalLDOLogic_VIA1 $T=86590 17140 0 0 $X=86340 $Y=16910
X3598 1 DigitalLDOLogic_VIA1 $T=86590 21220 0 0 $X=86340 $Y=20990
X3599 1 DigitalLDOLogic_VIA1 $T=86590 25300 0 0 $X=86340 $Y=25070
X3600 1 DigitalLDOLogic_VIA1 $T=86590 29380 0 0 $X=86340 $Y=29150
X3601 1 DigitalLDOLogic_VIA1 $T=86590 33460 0 0 $X=86340 $Y=33230
X3602 1 DigitalLDOLogic_VIA1 $T=86590 37540 0 0 $X=86340 $Y=37310
X3603 1 DigitalLDOLogic_VIA1 $T=86590 41620 0 0 $X=86340 $Y=41390
X3604 1 DigitalLDOLogic_VIA1 $T=86590 45700 0 0 $X=86340 $Y=45470
X3605 1 DigitalLDOLogic_VIA1 $T=86590 49780 0 0 $X=86340 $Y=49550
X3606 1 DigitalLDOLogic_VIA1 $T=86590 53860 0 0 $X=86340 $Y=53630
X3607 1 DigitalLDOLogic_VIA1 $T=86590 57940 0 0 $X=86340 $Y=57710
X3608 2 DigitalLDOLogic_VIA1 $T=88430 11700 0 0 $X=88180 $Y=11470
X3609 2 DigitalLDOLogic_VIA1 $T=88430 15780 0 0 $X=88180 $Y=15550
X3610 2 DigitalLDOLogic_VIA1 $T=88430 19860 0 0 $X=88180 $Y=19630
X3611 2 DigitalLDOLogic_VIA1 $T=88430 23940 0 0 $X=88180 $Y=23710
X3612 2 DigitalLDOLogic_VIA1 $T=88430 28020 0 0 $X=88180 $Y=27790
X3613 2 DigitalLDOLogic_VIA1 $T=88430 32100 0 0 $X=88180 $Y=31870
X3614 2 DigitalLDOLogic_VIA1 $T=88430 36180 0 0 $X=88180 $Y=35950
X3615 2 DigitalLDOLogic_VIA1 $T=88430 40260 0 0 $X=88180 $Y=40030
X3616 2 DigitalLDOLogic_VIA1 $T=88430 44340 0 0 $X=88180 $Y=44110
X3617 2 DigitalLDOLogic_VIA1 $T=88430 48420 0 0 $X=88180 $Y=48190
X3618 2 DigitalLDOLogic_VIA1 $T=88430 52500 0 0 $X=88180 $Y=52270
X3619 2 DigitalLDOLogic_VIA1 $T=88430 56580 0 0 $X=88180 $Y=56350
X3620 1 DigitalLDOLogic_VIA1 $T=89350 13060 0 0 $X=89100 $Y=12830
X3621 1 DigitalLDOLogic_VIA1 $T=89350 17140 0 0 $X=89100 $Y=16910
X3622 1 DigitalLDOLogic_VIA1 $T=89350 21220 0 0 $X=89100 $Y=20990
X3623 1 DigitalLDOLogic_VIA1 $T=89350 25300 0 0 $X=89100 $Y=25070
X3624 1 DigitalLDOLogic_VIA1 $T=89350 29380 0 0 $X=89100 $Y=29150
X3625 1 DigitalLDOLogic_VIA1 $T=89350 33460 0 0 $X=89100 $Y=33230
X3626 1 DigitalLDOLogic_VIA1 $T=89350 37540 0 0 $X=89100 $Y=37310
X3627 1 DigitalLDOLogic_VIA1 $T=89350 41620 0 0 $X=89100 $Y=41390
X3628 1 DigitalLDOLogic_VIA1 $T=89350 45700 0 0 $X=89100 $Y=45470
X3629 1 DigitalLDOLogic_VIA1 $T=89350 49780 0 0 $X=89100 $Y=49550
X3630 1 DigitalLDOLogic_VIA1 $T=89350 53860 0 0 $X=89100 $Y=53630
X3631 1 DigitalLDOLogic_VIA1 $T=89350 57940 0 0 $X=89100 $Y=57710
X3632 2 DigitalLDOLogic_VIA1 $T=91190 11700 0 0 $X=90940 $Y=11470
X3633 2 DigitalLDOLogic_VIA1 $T=91190 15780 0 0 $X=90940 $Y=15550
X3634 2 DigitalLDOLogic_VIA1 $T=91190 19860 0 0 $X=90940 $Y=19630
X3635 2 DigitalLDOLogic_VIA1 $T=91190 23940 0 0 $X=90940 $Y=23710
X3636 2 DigitalLDOLogic_VIA1 $T=91190 28020 0 0 $X=90940 $Y=27790
X3637 2 DigitalLDOLogic_VIA1 $T=91190 32100 0 0 $X=90940 $Y=31870
X3638 2 DigitalLDOLogic_VIA1 $T=91190 36180 0 0 $X=90940 $Y=35950
X3639 2 DigitalLDOLogic_VIA1 $T=91190 40260 0 0 $X=90940 $Y=40030
X3640 2 DigitalLDOLogic_VIA1 $T=91190 44340 0 0 $X=90940 $Y=44110
X3641 2 DigitalLDOLogic_VIA1 $T=91190 48420 0 0 $X=90940 $Y=48190
X3642 2 DigitalLDOLogic_VIA1 $T=91190 52500 0 0 $X=90940 $Y=52270
X3643 2 DigitalLDOLogic_VIA1 $T=91190 56580 0 0 $X=90940 $Y=56350
X3644 1 DigitalLDOLogic_VIA1 $T=92110 13060 0 0 $X=91860 $Y=12830
X3645 1 DigitalLDOLogic_VIA1 $T=92110 17140 0 0 $X=91860 $Y=16910
X3646 1 DigitalLDOLogic_VIA1 $T=92110 21220 0 0 $X=91860 $Y=20990
X3647 1 DigitalLDOLogic_VIA1 $T=92110 25300 0 0 $X=91860 $Y=25070
X3648 1 DigitalLDOLogic_VIA1 $T=92110 29380 0 0 $X=91860 $Y=29150
X3649 1 DigitalLDOLogic_VIA1 $T=92110 33460 0 0 $X=91860 $Y=33230
X3650 1 DigitalLDOLogic_VIA1 $T=92110 37540 0 0 $X=91860 $Y=37310
X3651 1 DigitalLDOLogic_VIA1 $T=92110 41620 0 0 $X=91860 $Y=41390
X3652 1 DigitalLDOLogic_VIA1 $T=92110 45700 0 0 $X=91860 $Y=45470
X3653 1 DigitalLDOLogic_VIA1 $T=92110 49780 0 0 $X=91860 $Y=49550
X3654 1 DigitalLDOLogic_VIA1 $T=92110 53860 0 0 $X=91860 $Y=53630
X3655 1 DigitalLDOLogic_VIA1 $T=92110 57940 0 0 $X=91860 $Y=57710
X3656 2 DigitalLDOLogic_VIA1 $T=93950 11700 0 0 $X=93700 $Y=11470
X3657 2 DigitalLDOLogic_VIA1 $T=93950 15780 0 0 $X=93700 $Y=15550
X3658 2 DigitalLDOLogic_VIA1 $T=93950 19860 0 0 $X=93700 $Y=19630
X3659 2 DigitalLDOLogic_VIA1 $T=93950 23940 0 0 $X=93700 $Y=23710
X3660 2 DigitalLDOLogic_VIA1 $T=93950 28020 0 0 $X=93700 $Y=27790
X3661 2 DigitalLDOLogic_VIA1 $T=93950 32100 0 0 $X=93700 $Y=31870
X3662 2 DigitalLDOLogic_VIA1 $T=93950 36180 0 0 $X=93700 $Y=35950
X3663 2 DigitalLDOLogic_VIA1 $T=93950 40260 0 0 $X=93700 $Y=40030
X3664 2 DigitalLDOLogic_VIA1 $T=93950 44340 0 0 $X=93700 $Y=44110
X3665 2 DigitalLDOLogic_VIA1 $T=93950 48420 0 0 $X=93700 $Y=48190
X3666 2 DigitalLDOLogic_VIA1 $T=93950 52500 0 0 $X=93700 $Y=52270
X3667 2 DigitalLDOLogic_VIA1 $T=93950 56580 0 0 $X=93700 $Y=56350
X3668 1 DigitalLDOLogic_VIA1 $T=94870 13060 0 0 $X=94620 $Y=12830
X3669 1 DigitalLDOLogic_VIA1 $T=94870 17140 0 0 $X=94620 $Y=16910
X3670 1 DigitalLDOLogic_VIA1 $T=94870 21220 0 0 $X=94620 $Y=20990
X3671 1 DigitalLDOLogic_VIA1 $T=94870 25300 0 0 $X=94620 $Y=25070
X3672 1 DigitalLDOLogic_VIA1 $T=94870 29380 0 0 $X=94620 $Y=29150
X3673 1 DigitalLDOLogic_VIA1 $T=94870 33460 0 0 $X=94620 $Y=33230
X3674 1 DigitalLDOLogic_VIA1 $T=94870 37540 0 0 $X=94620 $Y=37310
X3675 1 DigitalLDOLogic_VIA1 $T=94870 41620 0 0 $X=94620 $Y=41390
X3676 1 DigitalLDOLogic_VIA1 $T=94870 45700 0 0 $X=94620 $Y=45470
X3677 1 DigitalLDOLogic_VIA1 $T=94870 49780 0 0 $X=94620 $Y=49550
X3678 1 DigitalLDOLogic_VIA1 $T=94870 53860 0 0 $X=94620 $Y=53630
X3679 1 DigitalLDOLogic_VIA1 $T=94870 57940 0 0 $X=94620 $Y=57710
X3680 2 DigitalLDOLogic_VIA1 $T=96710 11700 0 0 $X=96460 $Y=11470
X3681 2 DigitalLDOLogic_VIA1 $T=96710 15780 0 0 $X=96460 $Y=15550
X3682 2 DigitalLDOLogic_VIA1 $T=96710 19860 0 0 $X=96460 $Y=19630
X3683 2 DigitalLDOLogic_VIA1 $T=96710 23940 0 0 $X=96460 $Y=23710
X3684 2 DigitalLDOLogic_VIA1 $T=96710 28020 0 0 $X=96460 $Y=27790
X3685 2 DigitalLDOLogic_VIA1 $T=96710 32100 0 0 $X=96460 $Y=31870
X3686 2 DigitalLDOLogic_VIA1 $T=96710 36180 0 0 $X=96460 $Y=35950
X3687 2 DigitalLDOLogic_VIA1 $T=96710 40260 0 0 $X=96460 $Y=40030
X3688 2 DigitalLDOLogic_VIA1 $T=96710 44340 0 0 $X=96460 $Y=44110
X3689 2 DigitalLDOLogic_VIA1 $T=96710 48420 0 0 $X=96460 $Y=48190
X3690 2 DigitalLDOLogic_VIA1 $T=96710 52500 0 0 $X=96460 $Y=52270
X3691 2 DigitalLDOLogic_VIA1 $T=96710 56580 0 0 $X=96460 $Y=56350
X3692 1 DigitalLDOLogic_VIA1 $T=97630 13060 0 0 $X=97380 $Y=12830
X3693 1 DigitalLDOLogic_VIA1 $T=97630 17140 0 0 $X=97380 $Y=16910
X3694 1 DigitalLDOLogic_VIA1 $T=97630 21220 0 0 $X=97380 $Y=20990
X3695 1 DigitalLDOLogic_VIA1 $T=97630 25300 0 0 $X=97380 $Y=25070
X3696 1 DigitalLDOLogic_VIA1 $T=97630 29380 0 0 $X=97380 $Y=29150
X3697 1 DigitalLDOLogic_VIA1 $T=97630 33460 0 0 $X=97380 $Y=33230
X3698 1 DigitalLDOLogic_VIA1 $T=97630 37540 0 0 $X=97380 $Y=37310
X3699 1 DigitalLDOLogic_VIA1 $T=97630 41620 0 0 $X=97380 $Y=41390
X3700 1 DigitalLDOLogic_VIA1 $T=97630 45700 0 0 $X=97380 $Y=45470
X3701 1 DigitalLDOLogic_VIA1 $T=97630 49780 0 0 $X=97380 $Y=49550
X3702 1 DigitalLDOLogic_VIA1 $T=97630 53860 0 0 $X=97380 $Y=53630
X3703 1 DigitalLDOLogic_VIA1 $T=97630 57940 0 0 $X=97380 $Y=57710
X3704 2 DigitalLDOLogic_VIA1 $T=99470 11700 0 0 $X=99220 $Y=11470
X3705 2 DigitalLDOLogic_VIA1 $T=99470 15780 0 0 $X=99220 $Y=15550
X3706 2 DigitalLDOLogic_VIA1 $T=99470 19860 0 0 $X=99220 $Y=19630
X3707 2 DigitalLDOLogic_VIA1 $T=99470 23940 0 0 $X=99220 $Y=23710
X3708 2 DigitalLDOLogic_VIA1 $T=99470 28020 0 0 $X=99220 $Y=27790
X3709 2 DigitalLDOLogic_VIA1 $T=99470 32100 0 0 $X=99220 $Y=31870
X3710 2 DigitalLDOLogic_VIA1 $T=99470 36180 0 0 $X=99220 $Y=35950
X3711 2 DigitalLDOLogic_VIA1 $T=99470 40260 0 0 $X=99220 $Y=40030
X3712 2 DigitalLDOLogic_VIA1 $T=99470 44340 0 0 $X=99220 $Y=44110
X3713 2 DigitalLDOLogic_VIA1 $T=99470 48420 0 0 $X=99220 $Y=48190
X3714 2 DigitalLDOLogic_VIA1 $T=99470 52500 0 0 $X=99220 $Y=52270
X3715 2 DigitalLDOLogic_VIA1 $T=99470 56580 0 0 $X=99220 $Y=56350
X3716 1 DigitalLDOLogic_VIA1 $T=100390 13060 0 0 $X=100140 $Y=12830
X3717 1 DigitalLDOLogic_VIA1 $T=100390 17140 0 0 $X=100140 $Y=16910
X3718 1 DigitalLDOLogic_VIA1 $T=100390 21220 0 0 $X=100140 $Y=20990
X3719 1 DigitalLDOLogic_VIA1 $T=100390 25300 0 0 $X=100140 $Y=25070
X3720 1 DigitalLDOLogic_VIA1 $T=100390 29380 0 0 $X=100140 $Y=29150
X3721 1 DigitalLDOLogic_VIA1 $T=100390 33460 0 0 $X=100140 $Y=33230
X3722 1 DigitalLDOLogic_VIA1 $T=100390 37540 0 0 $X=100140 $Y=37310
X3723 1 DigitalLDOLogic_VIA1 $T=100390 41620 0 0 $X=100140 $Y=41390
X3724 1 DigitalLDOLogic_VIA1 $T=100390 45700 0 0 $X=100140 $Y=45470
X3725 1 DigitalLDOLogic_VIA1 $T=100390 49780 0 0 $X=100140 $Y=49550
X3726 1 DigitalLDOLogic_VIA1 $T=100390 53860 0 0 $X=100140 $Y=53630
X3727 1 DigitalLDOLogic_VIA1 $T=100390 57940 0 0 $X=100140 $Y=57710
X3728 2 DigitalLDOLogic_VIA1 $T=102230 11700 0 0 $X=101980 $Y=11470
X3729 2 DigitalLDOLogic_VIA1 $T=102230 15780 0 0 $X=101980 $Y=15550
X3730 2 DigitalLDOLogic_VIA1 $T=102230 19860 0 0 $X=101980 $Y=19630
X3731 2 DigitalLDOLogic_VIA1 $T=102230 23940 0 0 $X=101980 $Y=23710
X3732 2 DigitalLDOLogic_VIA1 $T=102230 28020 0 0 $X=101980 $Y=27790
X3733 2 DigitalLDOLogic_VIA1 $T=102230 32100 0 0 $X=101980 $Y=31870
X3734 2 DigitalLDOLogic_VIA1 $T=102230 36180 0 0 $X=101980 $Y=35950
X3735 2 DigitalLDOLogic_VIA1 $T=102230 40260 0 0 $X=101980 $Y=40030
X3736 2 DigitalLDOLogic_VIA1 $T=102230 44340 0 0 $X=101980 $Y=44110
X3737 2 DigitalLDOLogic_VIA1 $T=102230 48420 0 0 $X=101980 $Y=48190
X3738 2 DigitalLDOLogic_VIA1 $T=102230 52500 0 0 $X=101980 $Y=52270
X3739 2 DigitalLDOLogic_VIA1 $T=102230 56580 0 0 $X=101980 $Y=56350
X3740 1 DigitalLDOLogic_VIA1 $T=103150 13060 0 0 $X=102900 $Y=12830
X3741 1 DigitalLDOLogic_VIA1 $T=103150 17140 0 0 $X=102900 $Y=16910
X3742 1 DigitalLDOLogic_VIA1 $T=103150 21220 0 0 $X=102900 $Y=20990
X3743 1 DigitalLDOLogic_VIA1 $T=103150 25300 0 0 $X=102900 $Y=25070
X3744 1 DigitalLDOLogic_VIA1 $T=103150 29380 0 0 $X=102900 $Y=29150
X3745 1 DigitalLDOLogic_VIA1 $T=103150 33460 0 0 $X=102900 $Y=33230
X3746 1 DigitalLDOLogic_VIA1 $T=103150 37540 0 0 $X=102900 $Y=37310
X3747 1 DigitalLDOLogic_VIA1 $T=103150 41620 0 0 $X=102900 $Y=41390
X3748 1 DigitalLDOLogic_VIA1 $T=103150 45700 0 0 $X=102900 $Y=45470
X3749 1 DigitalLDOLogic_VIA1 $T=103150 49780 0 0 $X=102900 $Y=49550
X3750 1 DigitalLDOLogic_VIA1 $T=103150 53860 0 0 $X=102900 $Y=53630
X3751 1 DigitalLDOLogic_VIA1 $T=103150 57940 0 0 $X=102900 $Y=57710
X3752 2 DigitalLDOLogic_VIA1 $T=104990 11700 0 0 $X=104740 $Y=11470
X3753 2 DigitalLDOLogic_VIA1 $T=104990 15780 0 0 $X=104740 $Y=15550
X3754 2 DigitalLDOLogic_VIA1 $T=104990 19860 0 0 $X=104740 $Y=19630
X3755 2 DigitalLDOLogic_VIA1 $T=104990 23940 0 0 $X=104740 $Y=23710
X3756 2 DigitalLDOLogic_VIA1 $T=104990 28020 0 0 $X=104740 $Y=27790
X3757 2 DigitalLDOLogic_VIA1 $T=104990 32100 0 0 $X=104740 $Y=31870
X3758 2 DigitalLDOLogic_VIA1 $T=104990 36180 0 0 $X=104740 $Y=35950
X3759 2 DigitalLDOLogic_VIA1 $T=104990 40260 0 0 $X=104740 $Y=40030
X3760 2 DigitalLDOLogic_VIA1 $T=104990 44340 0 0 $X=104740 $Y=44110
X3761 2 DigitalLDOLogic_VIA1 $T=104990 48420 0 0 $X=104740 $Y=48190
X3762 2 DigitalLDOLogic_VIA1 $T=104990 52500 0 0 $X=104740 $Y=52270
X3763 2 DigitalLDOLogic_VIA1 $T=104990 56580 0 0 $X=104740 $Y=56350
X3764 1 DigitalLDOLogic_VIA1 $T=105910 13060 0 0 $X=105660 $Y=12830
X3765 1 DigitalLDOLogic_VIA1 $T=105910 17140 0 0 $X=105660 $Y=16910
X3766 1 DigitalLDOLogic_VIA1 $T=105910 21220 0 0 $X=105660 $Y=20990
X3767 1 DigitalLDOLogic_VIA1 $T=105910 25300 0 0 $X=105660 $Y=25070
X3768 1 DigitalLDOLogic_VIA1 $T=105910 29380 0 0 $X=105660 $Y=29150
X3769 1 DigitalLDOLogic_VIA1 $T=105910 33460 0 0 $X=105660 $Y=33230
X3770 1 DigitalLDOLogic_VIA1 $T=105910 37540 0 0 $X=105660 $Y=37310
X3771 1 DigitalLDOLogic_VIA1 $T=105910 41620 0 0 $X=105660 $Y=41390
X3772 1 DigitalLDOLogic_VIA1 $T=105910 45700 0 0 $X=105660 $Y=45470
X3773 1 DigitalLDOLogic_VIA1 $T=105910 49780 0 0 $X=105660 $Y=49550
X3774 1 DigitalLDOLogic_VIA1 $T=105910 53860 0 0 $X=105660 $Y=53630
X3775 1 DigitalLDOLogic_VIA1 $T=105910 57940 0 0 $X=105660 $Y=57710
X3776 2 DigitalLDOLogic_VIA1 $T=107750 11700 0 0 $X=107500 $Y=11470
X3777 2 DigitalLDOLogic_VIA1 $T=107750 15780 0 0 $X=107500 $Y=15550
X3778 2 DigitalLDOLogic_VIA1 $T=107750 19860 0 0 $X=107500 $Y=19630
X3779 2 DigitalLDOLogic_VIA1 $T=107750 23940 0 0 $X=107500 $Y=23710
X3780 2 DigitalLDOLogic_VIA1 $T=107750 28020 0 0 $X=107500 $Y=27790
X3781 2 DigitalLDOLogic_VIA1 $T=107750 32100 0 0 $X=107500 $Y=31870
X3782 2 DigitalLDOLogic_VIA1 $T=107750 36180 0 0 $X=107500 $Y=35950
X3783 2 DigitalLDOLogic_VIA1 $T=107750 40260 0 0 $X=107500 $Y=40030
X3784 2 DigitalLDOLogic_VIA1 $T=107750 44340 0 0 $X=107500 $Y=44110
X3785 2 DigitalLDOLogic_VIA1 $T=107750 48420 0 0 $X=107500 $Y=48190
X3786 2 DigitalLDOLogic_VIA1 $T=107750 52500 0 0 $X=107500 $Y=52270
X3787 2 DigitalLDOLogic_VIA1 $T=107750 56580 0 0 $X=107500 $Y=56350
X3788 1 DigitalLDOLogic_VIA1 $T=108670 13060 0 0 $X=108420 $Y=12830
X3789 1 DigitalLDOLogic_VIA1 $T=108670 17140 0 0 $X=108420 $Y=16910
X3790 1 DigitalLDOLogic_VIA1 $T=108670 21220 0 0 $X=108420 $Y=20990
X3791 1 DigitalLDOLogic_VIA1 $T=108670 25300 0 0 $X=108420 $Y=25070
X3792 1 DigitalLDOLogic_VIA1 $T=108670 29380 0 0 $X=108420 $Y=29150
X3793 1 DigitalLDOLogic_VIA1 $T=108670 33460 0 0 $X=108420 $Y=33230
X3794 1 DigitalLDOLogic_VIA1 $T=108670 37540 0 0 $X=108420 $Y=37310
X3795 1 DigitalLDOLogic_VIA1 $T=108670 41620 0 0 $X=108420 $Y=41390
X3796 1 DigitalLDOLogic_VIA1 $T=108670 45700 0 0 $X=108420 $Y=45470
X3797 1 DigitalLDOLogic_VIA1 $T=108670 49780 0 0 $X=108420 $Y=49550
X3798 1 DigitalLDOLogic_VIA1 $T=108670 53860 0 0 $X=108420 $Y=53630
X3799 1 DigitalLDOLogic_VIA1 $T=108670 57940 0 0 $X=108420 $Y=57710
X3800 2 DigitalLDOLogic_VIA1 $T=110510 11700 0 0 $X=110260 $Y=11470
X3801 2 DigitalLDOLogic_VIA1 $T=110510 15780 0 0 $X=110260 $Y=15550
X3802 2 DigitalLDOLogic_VIA1 $T=110510 19860 0 0 $X=110260 $Y=19630
X3803 2 DigitalLDOLogic_VIA1 $T=110510 23940 0 0 $X=110260 $Y=23710
X3804 2 DigitalLDOLogic_VIA1 $T=110510 28020 0 0 $X=110260 $Y=27790
X3805 2 DigitalLDOLogic_VIA1 $T=110510 32100 0 0 $X=110260 $Y=31870
X3806 2 DigitalLDOLogic_VIA1 $T=110510 36180 0 0 $X=110260 $Y=35950
X3807 2 DigitalLDOLogic_VIA1 $T=110510 40260 0 0 $X=110260 $Y=40030
X3808 2 DigitalLDOLogic_VIA1 $T=110510 44340 0 0 $X=110260 $Y=44110
X3809 2 DigitalLDOLogic_VIA1 $T=110510 48420 0 0 $X=110260 $Y=48190
X3810 2 DigitalLDOLogic_VIA1 $T=110510 52500 0 0 $X=110260 $Y=52270
X3811 2 DigitalLDOLogic_VIA1 $T=110510 56580 0 0 $X=110260 $Y=56350
X3812 1 DigitalLDOLogic_VIA1 $T=111430 13060 0 0 $X=111180 $Y=12830
X3813 1 DigitalLDOLogic_VIA1 $T=111430 17140 0 0 $X=111180 $Y=16910
X3814 1 DigitalLDOLogic_VIA1 $T=111430 21220 0 0 $X=111180 $Y=20990
X3815 1 DigitalLDOLogic_VIA1 $T=111430 25300 0 0 $X=111180 $Y=25070
X3816 1 DigitalLDOLogic_VIA1 $T=111430 29380 0 0 $X=111180 $Y=29150
X3817 1 DigitalLDOLogic_VIA1 $T=111430 33460 0 0 $X=111180 $Y=33230
X3818 1 DigitalLDOLogic_VIA1 $T=111430 37540 0 0 $X=111180 $Y=37310
X3819 1 DigitalLDOLogic_VIA1 $T=111430 41620 0 0 $X=111180 $Y=41390
X3820 1 DigitalLDOLogic_VIA1 $T=111430 45700 0 0 $X=111180 $Y=45470
X3821 1 DigitalLDOLogic_VIA1 $T=111430 49780 0 0 $X=111180 $Y=49550
X3822 1 DigitalLDOLogic_VIA1 $T=111430 53860 0 0 $X=111180 $Y=53630
X3823 1 DigitalLDOLogic_VIA1 $T=111430 57940 0 0 $X=111180 $Y=57710
X3824 2 DigitalLDOLogic_VIA1 $T=113270 11700 0 0 $X=113020 $Y=11470
X3825 2 DigitalLDOLogic_VIA1 $T=113270 15780 0 0 $X=113020 $Y=15550
X3826 2 DigitalLDOLogic_VIA1 $T=113270 19860 0 0 $X=113020 $Y=19630
X3827 2 DigitalLDOLogic_VIA1 $T=113270 23940 0 0 $X=113020 $Y=23710
X3828 2 DigitalLDOLogic_VIA1 $T=113270 28020 0 0 $X=113020 $Y=27790
X3829 2 DigitalLDOLogic_VIA1 $T=113270 32100 0 0 $X=113020 $Y=31870
X3830 2 DigitalLDOLogic_VIA1 $T=113270 36180 0 0 $X=113020 $Y=35950
X3831 2 DigitalLDOLogic_VIA1 $T=113270 40260 0 0 $X=113020 $Y=40030
X3832 2 DigitalLDOLogic_VIA1 $T=113270 44340 0 0 $X=113020 $Y=44110
X3833 2 DigitalLDOLogic_VIA1 $T=113270 48420 0 0 $X=113020 $Y=48190
X3834 2 DigitalLDOLogic_VIA1 $T=113270 52500 0 0 $X=113020 $Y=52270
X3835 2 DigitalLDOLogic_VIA1 $T=113270 56580 0 0 $X=113020 $Y=56350
X3836 1 DigitalLDOLogic_VIA1 $T=114190 13060 0 0 $X=113940 $Y=12830
X3837 1 DigitalLDOLogic_VIA1 $T=114190 17140 0 0 $X=113940 $Y=16910
X3838 1 DigitalLDOLogic_VIA1 $T=114190 21220 0 0 $X=113940 $Y=20990
X3839 1 DigitalLDOLogic_VIA1 $T=114190 25300 0 0 $X=113940 $Y=25070
X3840 1 DigitalLDOLogic_VIA1 $T=114190 29380 0 0 $X=113940 $Y=29150
X3841 1 DigitalLDOLogic_VIA1 $T=114190 33460 0 0 $X=113940 $Y=33230
X3842 1 DigitalLDOLogic_VIA1 $T=114190 37540 0 0 $X=113940 $Y=37310
X3843 1 DigitalLDOLogic_VIA1 $T=114190 41620 0 0 $X=113940 $Y=41390
X3844 1 DigitalLDOLogic_VIA1 $T=114190 45700 0 0 $X=113940 $Y=45470
X3845 1 DigitalLDOLogic_VIA1 $T=114190 49780 0 0 $X=113940 $Y=49550
X3846 1 DigitalLDOLogic_VIA1 $T=114190 53860 0 0 $X=113940 $Y=53630
X3847 1 DigitalLDOLogic_VIA1 $T=114190 57940 0 0 $X=113940 $Y=57710
X3848 2 DigitalLDOLogic_VIA1 $T=116030 11700 0 0 $X=115780 $Y=11470
X3849 2 DigitalLDOLogic_VIA1 $T=116030 15780 0 0 $X=115780 $Y=15550
X3850 2 DigitalLDOLogic_VIA1 $T=116030 19860 0 0 $X=115780 $Y=19630
X3851 2 DigitalLDOLogic_VIA1 $T=116030 23940 0 0 $X=115780 $Y=23710
X3852 2 DigitalLDOLogic_VIA1 $T=116030 28020 0 0 $X=115780 $Y=27790
X3853 2 DigitalLDOLogic_VIA1 $T=116030 32100 0 0 $X=115780 $Y=31870
X3854 2 DigitalLDOLogic_VIA1 $T=116030 36180 0 0 $X=115780 $Y=35950
X3855 2 DigitalLDOLogic_VIA1 $T=116030 40260 0 0 $X=115780 $Y=40030
X3856 2 DigitalLDOLogic_VIA1 $T=116030 44340 0 0 $X=115780 $Y=44110
X3857 2 DigitalLDOLogic_VIA1 $T=116030 48420 0 0 $X=115780 $Y=48190
X3858 2 DigitalLDOLogic_VIA1 $T=116030 52500 0 0 $X=115780 $Y=52270
X3859 2 DigitalLDOLogic_VIA1 $T=116030 56580 0 0 $X=115780 $Y=56350
X3860 1 DigitalLDOLogic_VIA1 $T=116950 13060 0 0 $X=116700 $Y=12830
X3861 1 DigitalLDOLogic_VIA1 $T=116950 17140 0 0 $X=116700 $Y=16910
X3862 1 DigitalLDOLogic_VIA1 $T=116950 21220 0 0 $X=116700 $Y=20990
X3863 1 DigitalLDOLogic_VIA1 $T=116950 25300 0 0 $X=116700 $Y=25070
X3864 1 DigitalLDOLogic_VIA1 $T=116950 29380 0 0 $X=116700 $Y=29150
X3865 1 DigitalLDOLogic_VIA1 $T=116950 33460 0 0 $X=116700 $Y=33230
X3866 1 DigitalLDOLogic_VIA1 $T=116950 37540 0 0 $X=116700 $Y=37310
X3867 1 DigitalLDOLogic_VIA1 $T=116950 41620 0 0 $X=116700 $Y=41390
X3868 1 DigitalLDOLogic_VIA1 $T=116950 45700 0 0 $X=116700 $Y=45470
X3869 1 DigitalLDOLogic_VIA1 $T=116950 49780 0 0 $X=116700 $Y=49550
X3870 1 DigitalLDOLogic_VIA1 $T=116950 53860 0 0 $X=116700 $Y=53630
X3871 1 DigitalLDOLogic_VIA1 $T=116950 57940 0 0 $X=116700 $Y=57710
X3872 2 DigitalLDOLogic_VIA1 $T=118790 11700 0 0 $X=118540 $Y=11470
X3873 2 DigitalLDOLogic_VIA1 $T=118790 15780 0 0 $X=118540 $Y=15550
X3874 2 DigitalLDOLogic_VIA1 $T=118790 19860 0 0 $X=118540 $Y=19630
X3875 2 DigitalLDOLogic_VIA1 $T=118790 23940 0 0 $X=118540 $Y=23710
X3876 2 DigitalLDOLogic_VIA1 $T=118790 28020 0 0 $X=118540 $Y=27790
X3877 2 DigitalLDOLogic_VIA1 $T=118790 32100 0 0 $X=118540 $Y=31870
X3878 2 DigitalLDOLogic_VIA1 $T=118790 36180 0 0 $X=118540 $Y=35950
X3879 2 DigitalLDOLogic_VIA1 $T=118790 40260 0 0 $X=118540 $Y=40030
X3880 2 DigitalLDOLogic_VIA1 $T=118790 44340 0 0 $X=118540 $Y=44110
X3881 2 DigitalLDOLogic_VIA1 $T=118790 48420 0 0 $X=118540 $Y=48190
X3882 2 DigitalLDOLogic_VIA1 $T=118790 52500 0 0 $X=118540 $Y=52270
X3883 2 DigitalLDOLogic_VIA1 $T=118790 56580 0 0 $X=118540 $Y=56350
X3884 1 DigitalLDOLogic_VIA1 $T=119710 13060 0 0 $X=119460 $Y=12830
X3885 1 DigitalLDOLogic_VIA1 $T=119710 17140 0 0 $X=119460 $Y=16910
X3886 1 DigitalLDOLogic_VIA1 $T=119710 21220 0 0 $X=119460 $Y=20990
X3887 1 DigitalLDOLogic_VIA1 $T=119710 25300 0 0 $X=119460 $Y=25070
X3888 1 DigitalLDOLogic_VIA1 $T=119710 29380 0 0 $X=119460 $Y=29150
X3889 1 DigitalLDOLogic_VIA1 $T=119710 33460 0 0 $X=119460 $Y=33230
X3890 1 DigitalLDOLogic_VIA1 $T=119710 37540 0 0 $X=119460 $Y=37310
X3891 1 DigitalLDOLogic_VIA1 $T=119710 41620 0 0 $X=119460 $Y=41390
X3892 1 DigitalLDOLogic_VIA1 $T=119710 45700 0 0 $X=119460 $Y=45470
X3893 1 DigitalLDOLogic_VIA1 $T=119710 49780 0 0 $X=119460 $Y=49550
X3894 1 DigitalLDOLogic_VIA1 $T=119710 53860 0 0 $X=119460 $Y=53630
X3895 1 DigitalLDOLogic_VIA1 $T=119710 57940 0 0 $X=119460 $Y=57710
X3896 2 DigitalLDOLogic_VIA1 $T=121550 11700 0 0 $X=121300 $Y=11470
X3897 2 DigitalLDOLogic_VIA1 $T=121550 15780 0 0 $X=121300 $Y=15550
X3898 2 DigitalLDOLogic_VIA1 $T=121550 19860 0 0 $X=121300 $Y=19630
X3899 2 DigitalLDOLogic_VIA1 $T=121550 23940 0 0 $X=121300 $Y=23710
X3900 2 DigitalLDOLogic_VIA1 $T=121550 28020 0 0 $X=121300 $Y=27790
X3901 2 DigitalLDOLogic_VIA1 $T=121550 32100 0 0 $X=121300 $Y=31870
X3902 2 DigitalLDOLogic_VIA1 $T=121550 36180 0 0 $X=121300 $Y=35950
X3903 2 DigitalLDOLogic_VIA1 $T=121550 40260 0 0 $X=121300 $Y=40030
X3904 2 DigitalLDOLogic_VIA1 $T=121550 44340 0 0 $X=121300 $Y=44110
X3905 2 DigitalLDOLogic_VIA1 $T=121550 48420 0 0 $X=121300 $Y=48190
X3906 2 DigitalLDOLogic_VIA1 $T=121550 52500 0 0 $X=121300 $Y=52270
X3907 2 DigitalLDOLogic_VIA1 $T=121550 56580 0 0 $X=121300 $Y=56350
X3908 1 DigitalLDOLogic_VIA1 $T=122470 13060 0 0 $X=122220 $Y=12830
X3909 1 DigitalLDOLogic_VIA1 $T=122470 17140 0 0 $X=122220 $Y=16910
X3910 1 DigitalLDOLogic_VIA1 $T=122470 21220 0 0 $X=122220 $Y=20990
X3911 1 DigitalLDOLogic_VIA1 $T=122470 25300 0 0 $X=122220 $Y=25070
X3912 1 DigitalLDOLogic_VIA1 $T=122470 29380 0 0 $X=122220 $Y=29150
X3913 1 DigitalLDOLogic_VIA1 $T=122470 33460 0 0 $X=122220 $Y=33230
X3914 1 DigitalLDOLogic_VIA1 $T=122470 37540 0 0 $X=122220 $Y=37310
X3915 1 DigitalLDOLogic_VIA1 $T=122470 41620 0 0 $X=122220 $Y=41390
X3916 1 DigitalLDOLogic_VIA1 $T=122470 45700 0 0 $X=122220 $Y=45470
X3917 1 DigitalLDOLogic_VIA1 $T=122470 49780 0 0 $X=122220 $Y=49550
X3918 1 DigitalLDOLogic_VIA1 $T=122470 53860 0 0 $X=122220 $Y=53630
X3919 1 DigitalLDOLogic_VIA1 $T=122470 57940 0 0 $X=122220 $Y=57710
X3920 2 DigitalLDOLogic_VIA1 $T=124310 11700 0 0 $X=124060 $Y=11470
X3921 2 DigitalLDOLogic_VIA1 $T=124310 15780 0 0 $X=124060 $Y=15550
X3922 2 DigitalLDOLogic_VIA1 $T=124310 19860 0 0 $X=124060 $Y=19630
X3923 2 DigitalLDOLogic_VIA1 $T=124310 23940 0 0 $X=124060 $Y=23710
X3924 2 DigitalLDOLogic_VIA1 $T=124310 28020 0 0 $X=124060 $Y=27790
X3925 2 DigitalLDOLogic_VIA1 $T=124310 32100 0 0 $X=124060 $Y=31870
X3926 2 DigitalLDOLogic_VIA1 $T=124310 36180 0 0 $X=124060 $Y=35950
X3927 2 DigitalLDOLogic_VIA1 $T=124310 40260 0 0 $X=124060 $Y=40030
X3928 2 DigitalLDOLogic_VIA1 $T=124310 44340 0 0 $X=124060 $Y=44110
X3929 2 DigitalLDOLogic_VIA1 $T=124310 48420 0 0 $X=124060 $Y=48190
X3930 2 DigitalLDOLogic_VIA1 $T=124310 52500 0 0 $X=124060 $Y=52270
X3931 2 DigitalLDOLogic_VIA1 $T=124310 56580 0 0 $X=124060 $Y=56350
X3932 1 DigitalLDOLogic_VIA1 $T=125230 13060 0 0 $X=124980 $Y=12830
X3933 1 DigitalLDOLogic_VIA1 $T=125230 17140 0 0 $X=124980 $Y=16910
X3934 1 DigitalLDOLogic_VIA1 $T=125230 21220 0 0 $X=124980 $Y=20990
X3935 1 DigitalLDOLogic_VIA1 $T=125230 25300 0 0 $X=124980 $Y=25070
X3936 1 DigitalLDOLogic_VIA1 $T=125230 29380 0 0 $X=124980 $Y=29150
X3937 1 DigitalLDOLogic_VIA1 $T=125230 33460 0 0 $X=124980 $Y=33230
X3938 1 DigitalLDOLogic_VIA1 $T=125230 37540 0 0 $X=124980 $Y=37310
X3939 1 DigitalLDOLogic_VIA1 $T=125230 41620 0 0 $X=124980 $Y=41390
X3940 1 DigitalLDOLogic_VIA1 $T=125230 45700 0 0 $X=124980 $Y=45470
X3941 1 DigitalLDOLogic_VIA1 $T=125230 49780 0 0 $X=124980 $Y=49550
X3942 1 DigitalLDOLogic_VIA1 $T=125230 53860 0 0 $X=124980 $Y=53630
X3943 1 DigitalLDOLogic_VIA1 $T=125230 57940 0 0 $X=124980 $Y=57710
X3944 2 DigitalLDOLogic_VIA1 $T=127070 11700 0 0 $X=126820 $Y=11470
X3945 2 DigitalLDOLogic_VIA1 $T=127070 15780 0 0 $X=126820 $Y=15550
X3946 2 DigitalLDOLogic_VIA1 $T=127070 19860 0 0 $X=126820 $Y=19630
X3947 2 DigitalLDOLogic_VIA1 $T=127070 23940 0 0 $X=126820 $Y=23710
X3948 2 DigitalLDOLogic_VIA1 $T=127070 28020 0 0 $X=126820 $Y=27790
X3949 2 DigitalLDOLogic_VIA1 $T=127070 32100 0 0 $X=126820 $Y=31870
X3950 2 DigitalLDOLogic_VIA1 $T=127070 36180 0 0 $X=126820 $Y=35950
X3951 2 DigitalLDOLogic_VIA1 $T=127070 40260 0 0 $X=126820 $Y=40030
X3952 2 DigitalLDOLogic_VIA1 $T=127070 44340 0 0 $X=126820 $Y=44110
X3953 2 DigitalLDOLogic_VIA1 $T=127070 48420 0 0 $X=126820 $Y=48190
X3954 2 DigitalLDOLogic_VIA1 $T=127070 52500 0 0 $X=126820 $Y=52270
X3955 2 DigitalLDOLogic_VIA1 $T=127070 56580 0 0 $X=126820 $Y=56350
X3956 1 DigitalLDOLogic_VIA1 $T=127990 13060 0 0 $X=127740 $Y=12830
X3957 1 DigitalLDOLogic_VIA1 $T=127990 17140 0 0 $X=127740 $Y=16910
X3958 1 DigitalLDOLogic_VIA1 $T=127990 21220 0 0 $X=127740 $Y=20990
X3959 1 DigitalLDOLogic_VIA1 $T=127990 25300 0 0 $X=127740 $Y=25070
X3960 1 DigitalLDOLogic_VIA1 $T=127990 29380 0 0 $X=127740 $Y=29150
X3961 1 DigitalLDOLogic_VIA1 $T=127990 33460 0 0 $X=127740 $Y=33230
X3962 1 DigitalLDOLogic_VIA1 $T=127990 37540 0 0 $X=127740 $Y=37310
X3963 1 DigitalLDOLogic_VIA1 $T=127990 41620 0 0 $X=127740 $Y=41390
X3964 1 DigitalLDOLogic_VIA1 $T=127990 45700 0 0 $X=127740 $Y=45470
X3965 1 DigitalLDOLogic_VIA1 $T=127990 49780 0 0 $X=127740 $Y=49550
X3966 1 DigitalLDOLogic_VIA1 $T=127990 53860 0 0 $X=127740 $Y=53630
X3967 1 DigitalLDOLogic_VIA1 $T=127990 57940 0 0 $X=127740 $Y=57710
X3968 2 DigitalLDOLogic_VIA1 $T=129830 11700 0 0 $X=129580 $Y=11470
X3969 2 DigitalLDOLogic_VIA1 $T=129830 15780 0 0 $X=129580 $Y=15550
X3970 2 DigitalLDOLogic_VIA1 $T=129830 19860 0 0 $X=129580 $Y=19630
X3971 2 DigitalLDOLogic_VIA1 $T=129830 23940 0 0 $X=129580 $Y=23710
X3972 2 DigitalLDOLogic_VIA1 $T=129830 28020 0 0 $X=129580 $Y=27790
X3973 2 DigitalLDOLogic_VIA1 $T=129830 32100 0 0 $X=129580 $Y=31870
X3974 2 DigitalLDOLogic_VIA1 $T=129830 36180 0 0 $X=129580 $Y=35950
X3975 2 DigitalLDOLogic_VIA1 $T=129830 40260 0 0 $X=129580 $Y=40030
X3976 2 DigitalLDOLogic_VIA1 $T=129830 44340 0 0 $X=129580 $Y=44110
X3977 2 DigitalLDOLogic_VIA1 $T=129830 48420 0 0 $X=129580 $Y=48190
X3978 2 DigitalLDOLogic_VIA1 $T=129830 52500 0 0 $X=129580 $Y=52270
X3979 2 DigitalLDOLogic_VIA1 $T=129830 56580 0 0 $X=129580 $Y=56350
X3980 1 DigitalLDOLogic_VIA1 $T=130750 13060 0 0 $X=130500 $Y=12830
X3981 1 DigitalLDOLogic_VIA1 $T=130750 17140 0 0 $X=130500 $Y=16910
X3982 1 DigitalLDOLogic_VIA1 $T=130750 21220 0 0 $X=130500 $Y=20990
X3983 1 DigitalLDOLogic_VIA1 $T=130750 25300 0 0 $X=130500 $Y=25070
X3984 1 DigitalLDOLogic_VIA1 $T=130750 29380 0 0 $X=130500 $Y=29150
X3985 1 DigitalLDOLogic_VIA1 $T=130750 33460 0 0 $X=130500 $Y=33230
X3986 1 DigitalLDOLogic_VIA1 $T=130750 37540 0 0 $X=130500 $Y=37310
X3987 1 DigitalLDOLogic_VIA1 $T=130750 41620 0 0 $X=130500 $Y=41390
X3988 1 DigitalLDOLogic_VIA1 $T=130750 45700 0 0 $X=130500 $Y=45470
X3989 1 DigitalLDOLogic_VIA1 $T=130750 49780 0 0 $X=130500 $Y=49550
X3990 1 DigitalLDOLogic_VIA1 $T=130750 53860 0 0 $X=130500 $Y=53630
X3991 1 DigitalLDOLogic_VIA1 $T=130750 57940 0 0 $X=130500 $Y=57710
X3992 2 DigitalLDOLogic_VIA1 $T=132590 11700 0 0 $X=132340 $Y=11470
X3993 2 DigitalLDOLogic_VIA1 $T=132590 15780 0 0 $X=132340 $Y=15550
X3994 2 DigitalLDOLogic_VIA1 $T=132590 19860 0 0 $X=132340 $Y=19630
X3995 2 DigitalLDOLogic_VIA1 $T=132590 23940 0 0 $X=132340 $Y=23710
X3996 2 DigitalLDOLogic_VIA1 $T=132590 28020 0 0 $X=132340 $Y=27790
X3997 2 DigitalLDOLogic_VIA1 $T=132590 32100 0 0 $X=132340 $Y=31870
X3998 2 DigitalLDOLogic_VIA1 $T=132590 36180 0 0 $X=132340 $Y=35950
X3999 2 DigitalLDOLogic_VIA1 $T=132590 40260 0 0 $X=132340 $Y=40030
X4000 2 DigitalLDOLogic_VIA1 $T=132590 44340 0 0 $X=132340 $Y=44110
X4001 2 DigitalLDOLogic_VIA1 $T=132590 48420 0 0 $X=132340 $Y=48190
X4002 2 DigitalLDOLogic_VIA1 $T=132590 52500 0 0 $X=132340 $Y=52270
X4003 2 DigitalLDOLogic_VIA1 $T=132590 56580 0 0 $X=132340 $Y=56350
X4004 1 DigitalLDOLogic_VIA1 $T=133510 13060 0 0 $X=133260 $Y=12830
X4005 1 DigitalLDOLogic_VIA1 $T=133510 17140 0 0 $X=133260 $Y=16910
X4006 1 DigitalLDOLogic_VIA1 $T=133510 21220 0 0 $X=133260 $Y=20990
X4007 1 DigitalLDOLogic_VIA1 $T=133510 25300 0 0 $X=133260 $Y=25070
X4008 1 DigitalLDOLogic_VIA1 $T=133510 29380 0 0 $X=133260 $Y=29150
X4009 1 DigitalLDOLogic_VIA1 $T=133510 33460 0 0 $X=133260 $Y=33230
X4010 1 DigitalLDOLogic_VIA1 $T=133510 37540 0 0 $X=133260 $Y=37310
X4011 1 DigitalLDOLogic_VIA1 $T=133510 41620 0 0 $X=133260 $Y=41390
X4012 1 DigitalLDOLogic_VIA1 $T=133510 45700 0 0 $X=133260 $Y=45470
X4013 1 DigitalLDOLogic_VIA1 $T=133510 49780 0 0 $X=133260 $Y=49550
X4014 1 DigitalLDOLogic_VIA1 $T=133510 53860 0 0 $X=133260 $Y=53630
X4015 1 DigitalLDOLogic_VIA1 $T=133510 57940 0 0 $X=133260 $Y=57710
X4016 2 DigitalLDOLogic_VIA1 $T=135350 11700 0 0 $X=135100 $Y=11470
X4017 2 DigitalLDOLogic_VIA1 $T=135350 15780 0 0 $X=135100 $Y=15550
X4018 2 DigitalLDOLogic_VIA1 $T=135350 19860 0 0 $X=135100 $Y=19630
X4019 2 DigitalLDOLogic_VIA1 $T=135350 23940 0 0 $X=135100 $Y=23710
X4020 2 DigitalLDOLogic_VIA1 $T=135350 28020 0 0 $X=135100 $Y=27790
X4021 2 DigitalLDOLogic_VIA1 $T=135350 32100 0 0 $X=135100 $Y=31870
X4022 2 DigitalLDOLogic_VIA1 $T=135350 36180 0 0 $X=135100 $Y=35950
X4023 2 DigitalLDOLogic_VIA1 $T=135350 40260 0 0 $X=135100 $Y=40030
X4024 2 DigitalLDOLogic_VIA1 $T=135350 44340 0 0 $X=135100 $Y=44110
X4025 2 DigitalLDOLogic_VIA1 $T=135350 48420 0 0 $X=135100 $Y=48190
X4026 2 DigitalLDOLogic_VIA1 $T=135350 52500 0 0 $X=135100 $Y=52270
X4027 2 DigitalLDOLogic_VIA1 $T=135350 56580 0 0 $X=135100 $Y=56350
X4028 1 DigitalLDOLogic_VIA1 $T=136270 13060 0 0 $X=136020 $Y=12830
X4029 1 DigitalLDOLogic_VIA1 $T=136270 17140 0 0 $X=136020 $Y=16910
X4030 1 DigitalLDOLogic_VIA1 $T=136270 21220 0 0 $X=136020 $Y=20990
X4031 1 DigitalLDOLogic_VIA1 $T=136270 25300 0 0 $X=136020 $Y=25070
X4032 1 DigitalLDOLogic_VIA1 $T=136270 29380 0 0 $X=136020 $Y=29150
X4033 1 DigitalLDOLogic_VIA1 $T=136270 33460 0 0 $X=136020 $Y=33230
X4034 1 DigitalLDOLogic_VIA1 $T=136270 37540 0 0 $X=136020 $Y=37310
X4035 1 DigitalLDOLogic_VIA1 $T=136270 41620 0 0 $X=136020 $Y=41390
X4036 1 DigitalLDOLogic_VIA1 $T=136270 45700 0 0 $X=136020 $Y=45470
X4037 1 DigitalLDOLogic_VIA1 $T=136270 49780 0 0 $X=136020 $Y=49550
X4038 1 DigitalLDOLogic_VIA1 $T=136270 53860 0 0 $X=136020 $Y=53630
X4039 1 DigitalLDOLogic_VIA1 $T=136270 57940 0 0 $X=136020 $Y=57710
X4040 2 DigitalLDOLogic_VIA1 $T=138110 11700 0 0 $X=137860 $Y=11470
X4041 2 DigitalLDOLogic_VIA1 $T=138110 15780 0 0 $X=137860 $Y=15550
X4042 2 DigitalLDOLogic_VIA1 $T=138110 19860 0 0 $X=137860 $Y=19630
X4043 2 DigitalLDOLogic_VIA1 $T=138110 23940 0 0 $X=137860 $Y=23710
X4044 2 DigitalLDOLogic_VIA1 $T=138110 28020 0 0 $X=137860 $Y=27790
X4045 2 DigitalLDOLogic_VIA1 $T=138110 32100 0 0 $X=137860 $Y=31870
X4046 2 DigitalLDOLogic_VIA1 $T=138110 36180 0 0 $X=137860 $Y=35950
X4047 2 DigitalLDOLogic_VIA1 $T=138110 40260 0 0 $X=137860 $Y=40030
X4048 2 DigitalLDOLogic_VIA1 $T=138110 44340 0 0 $X=137860 $Y=44110
X4049 2 DigitalLDOLogic_VIA1 $T=138110 48420 0 0 $X=137860 $Y=48190
X4050 2 DigitalLDOLogic_VIA1 $T=138110 52500 0 0 $X=137860 $Y=52270
X4051 2 DigitalLDOLogic_VIA1 $T=138110 56580 0 0 $X=137860 $Y=56350
X4052 1 DigitalLDOLogic_VIA1 $T=139030 13060 0 0 $X=138780 $Y=12830
X4053 1 DigitalLDOLogic_VIA1 $T=139030 17140 0 0 $X=138780 $Y=16910
X4054 1 DigitalLDOLogic_VIA1 $T=139030 21220 0 0 $X=138780 $Y=20990
X4055 1 DigitalLDOLogic_VIA1 $T=139030 25300 0 0 $X=138780 $Y=25070
X4056 1 DigitalLDOLogic_VIA1 $T=139030 29380 0 0 $X=138780 $Y=29150
X4057 1 DigitalLDOLogic_VIA1 $T=139030 33460 0 0 $X=138780 $Y=33230
X4058 1 DigitalLDOLogic_VIA1 $T=139030 37540 0 0 $X=138780 $Y=37310
X4059 1 DigitalLDOLogic_VIA1 $T=139030 41620 0 0 $X=138780 $Y=41390
X4060 1 DigitalLDOLogic_VIA1 $T=139030 45700 0 0 $X=138780 $Y=45470
X4061 1 DigitalLDOLogic_VIA1 $T=139030 49780 0 0 $X=138780 $Y=49550
X4062 1 DigitalLDOLogic_VIA1 $T=139030 53860 0 0 $X=138780 $Y=53630
X4063 1 DigitalLDOLogic_VIA1 $T=139030 57940 0 0 $X=138780 $Y=57710
X4064 2 DigitalLDOLogic_VIA1 $T=140870 11700 0 0 $X=140620 $Y=11470
X4065 2 DigitalLDOLogic_VIA1 $T=140870 15780 0 0 $X=140620 $Y=15550
X4066 2 DigitalLDOLogic_VIA1 $T=140870 19860 0 0 $X=140620 $Y=19630
X4067 2 DigitalLDOLogic_VIA1 $T=140870 23940 0 0 $X=140620 $Y=23710
X4068 2 DigitalLDOLogic_VIA1 $T=140870 28020 0 0 $X=140620 $Y=27790
X4069 2 DigitalLDOLogic_VIA1 $T=140870 32100 0 0 $X=140620 $Y=31870
X4070 2 DigitalLDOLogic_VIA1 $T=140870 36180 0 0 $X=140620 $Y=35950
X4071 2 DigitalLDOLogic_VIA1 $T=140870 40260 0 0 $X=140620 $Y=40030
X4072 2 DigitalLDOLogic_VIA1 $T=140870 44340 0 0 $X=140620 $Y=44110
X4073 2 DigitalLDOLogic_VIA1 $T=140870 48420 0 0 $X=140620 $Y=48190
X4074 2 DigitalLDOLogic_VIA1 $T=140870 52500 0 0 $X=140620 $Y=52270
X4075 2 DigitalLDOLogic_VIA1 $T=140870 56580 0 0 $X=140620 $Y=56350
X4076 1 DigitalLDOLogic_VIA1 $T=141790 13060 0 0 $X=141540 $Y=12830
X4077 1 DigitalLDOLogic_VIA1 $T=141790 17140 0 0 $X=141540 $Y=16910
X4078 1 DigitalLDOLogic_VIA1 $T=141790 21220 0 0 $X=141540 $Y=20990
X4079 1 DigitalLDOLogic_VIA1 $T=141790 25300 0 0 $X=141540 $Y=25070
X4080 1 DigitalLDOLogic_VIA1 $T=141790 29380 0 0 $X=141540 $Y=29150
X4081 1 DigitalLDOLogic_VIA1 $T=141790 33460 0 0 $X=141540 $Y=33230
X4082 1 DigitalLDOLogic_VIA1 $T=141790 37540 0 0 $X=141540 $Y=37310
X4083 1 DigitalLDOLogic_VIA1 $T=141790 41620 0 0 $X=141540 $Y=41390
X4084 1 DigitalLDOLogic_VIA1 $T=141790 45700 0 0 $X=141540 $Y=45470
X4085 1 DigitalLDOLogic_VIA1 $T=141790 49780 0 0 $X=141540 $Y=49550
X4086 1 DigitalLDOLogic_VIA1 $T=141790 53860 0 0 $X=141540 $Y=53630
X4087 1 DigitalLDOLogic_VIA1 $T=141790 57940 0 0 $X=141540 $Y=57710
X4088 2 DigitalLDOLogic_VIA1 $T=143630 11700 0 0 $X=143380 $Y=11470
X4089 2 DigitalLDOLogic_VIA1 $T=143630 15780 0 0 $X=143380 $Y=15550
X4090 2 DigitalLDOLogic_VIA1 $T=143630 19860 0 0 $X=143380 $Y=19630
X4091 2 DigitalLDOLogic_VIA1 $T=143630 23940 0 0 $X=143380 $Y=23710
X4092 2 DigitalLDOLogic_VIA1 $T=143630 28020 0 0 $X=143380 $Y=27790
X4093 2 DigitalLDOLogic_VIA1 $T=143630 32100 0 0 $X=143380 $Y=31870
X4094 2 DigitalLDOLogic_VIA1 $T=143630 36180 0 0 $X=143380 $Y=35950
X4095 2 DigitalLDOLogic_VIA1 $T=143630 40260 0 0 $X=143380 $Y=40030
X4096 2 DigitalLDOLogic_VIA1 $T=143630 44340 0 0 $X=143380 $Y=44110
X4097 2 DigitalLDOLogic_VIA1 $T=143630 48420 0 0 $X=143380 $Y=48190
X4098 2 DigitalLDOLogic_VIA1 $T=143630 52500 0 0 $X=143380 $Y=52270
X4099 2 DigitalLDOLogic_VIA1 $T=143630 56580 0 0 $X=143380 $Y=56350
X4100 1 DigitalLDOLogic_VIA1 $T=144550 13060 0 0 $X=144300 $Y=12830
X4101 1 DigitalLDOLogic_VIA1 $T=144550 17140 0 0 $X=144300 $Y=16910
X4102 1 DigitalLDOLogic_VIA1 $T=144550 21220 0 0 $X=144300 $Y=20990
X4103 1 DigitalLDOLogic_VIA1 $T=144550 25300 0 0 $X=144300 $Y=25070
X4104 1 DigitalLDOLogic_VIA1 $T=144550 29380 0 0 $X=144300 $Y=29150
X4105 1 DigitalLDOLogic_VIA1 $T=144550 33460 0 0 $X=144300 $Y=33230
X4106 1 DigitalLDOLogic_VIA1 $T=144550 37540 0 0 $X=144300 $Y=37310
X4107 1 DigitalLDOLogic_VIA1 $T=144550 41620 0 0 $X=144300 $Y=41390
X4108 1 DigitalLDOLogic_VIA1 $T=144550 45700 0 0 $X=144300 $Y=45470
X4109 1 DigitalLDOLogic_VIA1 $T=144550 49780 0 0 $X=144300 $Y=49550
X4110 1 DigitalLDOLogic_VIA1 $T=144550 53860 0 0 $X=144300 $Y=53630
X4111 1 DigitalLDOLogic_VIA1 $T=144550 57940 0 0 $X=144300 $Y=57710
X4112 2 DigitalLDOLogic_VIA1 $T=146390 11700 0 0 $X=146140 $Y=11470
X4113 2 DigitalLDOLogic_VIA1 $T=146390 15780 0 0 $X=146140 $Y=15550
X4114 2 DigitalLDOLogic_VIA1 $T=146390 19860 0 0 $X=146140 $Y=19630
X4115 2 DigitalLDOLogic_VIA1 $T=146390 23940 0 0 $X=146140 $Y=23710
X4116 2 DigitalLDOLogic_VIA1 $T=146390 28020 0 0 $X=146140 $Y=27790
X4117 2 DigitalLDOLogic_VIA1 $T=146390 32100 0 0 $X=146140 $Y=31870
X4118 2 DigitalLDOLogic_VIA1 $T=146390 36180 0 0 $X=146140 $Y=35950
X4119 2 DigitalLDOLogic_VIA1 $T=146390 40260 0 0 $X=146140 $Y=40030
X4120 2 DigitalLDOLogic_VIA1 $T=146390 44340 0 0 $X=146140 $Y=44110
X4121 2 DigitalLDOLogic_VIA1 $T=146390 48420 0 0 $X=146140 $Y=48190
X4122 2 DigitalLDOLogic_VIA1 $T=146390 52500 0 0 $X=146140 $Y=52270
X4123 2 DigitalLDOLogic_VIA1 $T=146390 56580 0 0 $X=146140 $Y=56350
X4124 1 DigitalLDOLogic_VIA1 $T=147310 13060 0 0 $X=147060 $Y=12830
X4125 1 DigitalLDOLogic_VIA1 $T=147310 17140 0 0 $X=147060 $Y=16910
X4126 1 DigitalLDOLogic_VIA1 $T=147310 21220 0 0 $X=147060 $Y=20990
X4127 1 DigitalLDOLogic_VIA1 $T=147310 25300 0 0 $X=147060 $Y=25070
X4128 1 DigitalLDOLogic_VIA1 $T=147310 29380 0 0 $X=147060 $Y=29150
X4129 1 DigitalLDOLogic_VIA1 $T=147310 33460 0 0 $X=147060 $Y=33230
X4130 1 DigitalLDOLogic_VIA1 $T=147310 37540 0 0 $X=147060 $Y=37310
X4131 1 DigitalLDOLogic_VIA1 $T=147310 41620 0 0 $X=147060 $Y=41390
X4132 1 DigitalLDOLogic_VIA1 $T=147310 45700 0 0 $X=147060 $Y=45470
X4133 1 DigitalLDOLogic_VIA1 $T=147310 49780 0 0 $X=147060 $Y=49550
X4134 1 DigitalLDOLogic_VIA1 $T=147310 53860 0 0 $X=147060 $Y=53630
X4135 1 DigitalLDOLogic_VIA1 $T=147310 57940 0 0 $X=147060 $Y=57710
X4136 2 DigitalLDOLogic_VIA1 $T=149150 11700 0 0 $X=148900 $Y=11470
X4137 2 DigitalLDOLogic_VIA1 $T=149150 15780 0 0 $X=148900 $Y=15550
X4138 2 DigitalLDOLogic_VIA1 $T=149150 19860 0 0 $X=148900 $Y=19630
X4139 2 DigitalLDOLogic_VIA1 $T=149150 23940 0 0 $X=148900 $Y=23710
X4140 2 DigitalLDOLogic_VIA1 $T=149150 28020 0 0 $X=148900 $Y=27790
X4141 2 DigitalLDOLogic_VIA1 $T=149150 32100 0 0 $X=148900 $Y=31870
X4142 2 DigitalLDOLogic_VIA1 $T=149150 36180 0 0 $X=148900 $Y=35950
X4143 2 DigitalLDOLogic_VIA1 $T=149150 40260 0 0 $X=148900 $Y=40030
X4144 2 DigitalLDOLogic_VIA1 $T=149150 44340 0 0 $X=148900 $Y=44110
X4145 2 DigitalLDOLogic_VIA1 $T=149150 48420 0 0 $X=148900 $Y=48190
X4146 2 DigitalLDOLogic_VIA1 $T=149150 52500 0 0 $X=148900 $Y=52270
X4147 2 DigitalLDOLogic_VIA1 $T=149150 56580 0 0 $X=148900 $Y=56350
X4148 1 DigitalLDOLogic_VIA1 $T=150070 13060 0 0 $X=149820 $Y=12830
X4149 1 DigitalLDOLogic_VIA1 $T=150070 17140 0 0 $X=149820 $Y=16910
X4150 1 DigitalLDOLogic_VIA1 $T=150070 21220 0 0 $X=149820 $Y=20990
X4151 1 DigitalLDOLogic_VIA1 $T=150070 25300 0 0 $X=149820 $Y=25070
X4152 1 DigitalLDOLogic_VIA1 $T=150070 29380 0 0 $X=149820 $Y=29150
X4153 1 DigitalLDOLogic_VIA1 $T=150070 33460 0 0 $X=149820 $Y=33230
X4154 1 DigitalLDOLogic_VIA1 $T=150070 37540 0 0 $X=149820 $Y=37310
X4155 1 DigitalLDOLogic_VIA1 $T=150070 41620 0 0 $X=149820 $Y=41390
X4156 1 DigitalLDOLogic_VIA1 $T=150070 45700 0 0 $X=149820 $Y=45470
X4157 1 DigitalLDOLogic_VIA1 $T=150070 49780 0 0 $X=149820 $Y=49550
X4158 1 DigitalLDOLogic_VIA1 $T=150070 53860 0 0 $X=149820 $Y=53630
X4159 1 DigitalLDOLogic_VIA1 $T=150070 57940 0 0 $X=149820 $Y=57710
X4160 2 DigitalLDOLogic_VIA1 $T=151910 11700 0 0 $X=151660 $Y=11470
X4161 2 DigitalLDOLogic_VIA1 $T=151910 15780 0 0 $X=151660 $Y=15550
X4162 2 DigitalLDOLogic_VIA1 $T=151910 19860 0 0 $X=151660 $Y=19630
X4163 2 DigitalLDOLogic_VIA1 $T=151910 23940 0 0 $X=151660 $Y=23710
X4164 2 DigitalLDOLogic_VIA1 $T=151910 28020 0 0 $X=151660 $Y=27790
X4165 2 DigitalLDOLogic_VIA1 $T=151910 32100 0 0 $X=151660 $Y=31870
X4166 2 DigitalLDOLogic_VIA1 $T=151910 36180 0 0 $X=151660 $Y=35950
X4167 2 DigitalLDOLogic_VIA1 $T=151910 40260 0 0 $X=151660 $Y=40030
X4168 2 DigitalLDOLogic_VIA1 $T=151910 44340 0 0 $X=151660 $Y=44110
X4169 2 DigitalLDOLogic_VIA1 $T=151910 48420 0 0 $X=151660 $Y=48190
X4170 2 DigitalLDOLogic_VIA1 $T=151910 52500 0 0 $X=151660 $Y=52270
X4171 2 DigitalLDOLogic_VIA1 $T=151910 56580 0 0 $X=151660 $Y=56350
X4172 1 DigitalLDOLogic_VIA1 $T=152830 13060 0 0 $X=152580 $Y=12830
X4173 1 DigitalLDOLogic_VIA1 $T=152830 17140 0 0 $X=152580 $Y=16910
X4174 1 DigitalLDOLogic_VIA1 $T=152830 21220 0 0 $X=152580 $Y=20990
X4175 1 DigitalLDOLogic_VIA1 $T=152830 25300 0 0 $X=152580 $Y=25070
X4176 1 DigitalLDOLogic_VIA1 $T=152830 29380 0 0 $X=152580 $Y=29150
X4177 1 DigitalLDOLogic_VIA1 $T=152830 33460 0 0 $X=152580 $Y=33230
X4178 1 DigitalLDOLogic_VIA1 $T=152830 37540 0 0 $X=152580 $Y=37310
X4179 1 DigitalLDOLogic_VIA1 $T=152830 41620 0 0 $X=152580 $Y=41390
X4180 1 DigitalLDOLogic_VIA1 $T=152830 45700 0 0 $X=152580 $Y=45470
X4181 1 DigitalLDOLogic_VIA1 $T=152830 49780 0 0 $X=152580 $Y=49550
X4182 1 DigitalLDOLogic_VIA1 $T=152830 53860 0 0 $X=152580 $Y=53630
X4183 1 DigitalLDOLogic_VIA1 $T=152830 57940 0 0 $X=152580 $Y=57710
X4184 2 DigitalLDOLogic_VIA1 $T=154670 11700 0 0 $X=154420 $Y=11470
X4185 2 DigitalLDOLogic_VIA1 $T=154670 15780 0 0 $X=154420 $Y=15550
X4186 2 DigitalLDOLogic_VIA1 $T=154670 19860 0 0 $X=154420 $Y=19630
X4187 2 DigitalLDOLogic_VIA1 $T=154670 23940 0 0 $X=154420 $Y=23710
X4188 2 DigitalLDOLogic_VIA1 $T=154670 28020 0 0 $X=154420 $Y=27790
X4189 2 DigitalLDOLogic_VIA1 $T=154670 32100 0 0 $X=154420 $Y=31870
X4190 2 DigitalLDOLogic_VIA1 $T=154670 36180 0 0 $X=154420 $Y=35950
X4191 2 DigitalLDOLogic_VIA1 $T=154670 40260 0 0 $X=154420 $Y=40030
X4192 2 DigitalLDOLogic_VIA1 $T=154670 44340 0 0 $X=154420 $Y=44110
X4193 2 DigitalLDOLogic_VIA1 $T=154670 48420 0 0 $X=154420 $Y=48190
X4194 2 DigitalLDOLogic_VIA1 $T=154670 52500 0 0 $X=154420 $Y=52270
X4195 2 DigitalLDOLogic_VIA1 $T=154670 56580 0 0 $X=154420 $Y=56350
X4196 1 DigitalLDOLogic_VIA1 $T=155590 13060 0 0 $X=155340 $Y=12830
X4197 1 DigitalLDOLogic_VIA1 $T=155590 17140 0 0 $X=155340 $Y=16910
X4198 1 DigitalLDOLogic_VIA1 $T=155590 21220 0 0 $X=155340 $Y=20990
X4199 1 DigitalLDOLogic_VIA1 $T=155590 25300 0 0 $X=155340 $Y=25070
X4200 1 DigitalLDOLogic_VIA1 $T=155590 29380 0 0 $X=155340 $Y=29150
X4201 1 DigitalLDOLogic_VIA1 $T=155590 33460 0 0 $X=155340 $Y=33230
X4202 1 DigitalLDOLogic_VIA1 $T=155590 37540 0 0 $X=155340 $Y=37310
X4203 1 DigitalLDOLogic_VIA1 $T=155590 41620 0 0 $X=155340 $Y=41390
X4204 1 DigitalLDOLogic_VIA1 $T=155590 45700 0 0 $X=155340 $Y=45470
X4205 1 DigitalLDOLogic_VIA1 $T=155590 49780 0 0 $X=155340 $Y=49550
X4206 1 DigitalLDOLogic_VIA1 $T=155590 53860 0 0 $X=155340 $Y=53630
X4207 1 DigitalLDOLogic_VIA1 $T=155590 57940 0 0 $X=155340 $Y=57710
X4208 2 DigitalLDOLogic_VIA1 $T=157430 11700 0 0 $X=157180 $Y=11470
X4209 2 DigitalLDOLogic_VIA1 $T=157430 15780 0 0 $X=157180 $Y=15550
X4210 2 DigitalLDOLogic_VIA1 $T=157430 19860 0 0 $X=157180 $Y=19630
X4211 2 DigitalLDOLogic_VIA1 $T=157430 23940 0 0 $X=157180 $Y=23710
X4212 2 DigitalLDOLogic_VIA1 $T=157430 28020 0 0 $X=157180 $Y=27790
X4213 2 DigitalLDOLogic_VIA1 $T=157430 32100 0 0 $X=157180 $Y=31870
X4214 2 DigitalLDOLogic_VIA1 $T=157430 36180 0 0 $X=157180 $Y=35950
X4215 2 DigitalLDOLogic_VIA1 $T=157430 40260 0 0 $X=157180 $Y=40030
X4216 2 DigitalLDOLogic_VIA1 $T=157430 44340 0 0 $X=157180 $Y=44110
X4217 2 DigitalLDOLogic_VIA1 $T=157430 48420 0 0 $X=157180 $Y=48190
X4218 2 DigitalLDOLogic_VIA1 $T=157430 52500 0 0 $X=157180 $Y=52270
X4219 2 DigitalLDOLogic_VIA1 $T=157430 56580 0 0 $X=157180 $Y=56350
X4220 1 DigitalLDOLogic_VIA1 $T=158350 13060 0 0 $X=158100 $Y=12830
X4221 1 DigitalLDOLogic_VIA1 $T=158350 17140 0 0 $X=158100 $Y=16910
X4222 1 DigitalLDOLogic_VIA1 $T=158350 21220 0 0 $X=158100 $Y=20990
X4223 1 DigitalLDOLogic_VIA1 $T=158350 25300 0 0 $X=158100 $Y=25070
X4224 1 DigitalLDOLogic_VIA1 $T=158350 29380 0 0 $X=158100 $Y=29150
X4225 1 DigitalLDOLogic_VIA1 $T=158350 33460 0 0 $X=158100 $Y=33230
X4226 1 DigitalLDOLogic_VIA1 $T=158350 37540 0 0 $X=158100 $Y=37310
X4227 1 DigitalLDOLogic_VIA1 $T=158350 41620 0 0 $X=158100 $Y=41390
X4228 1 DigitalLDOLogic_VIA1 $T=158350 45700 0 0 $X=158100 $Y=45470
X4229 1 DigitalLDOLogic_VIA1 $T=158350 49780 0 0 $X=158100 $Y=49550
X4230 1 DigitalLDOLogic_VIA1 $T=158350 53860 0 0 $X=158100 $Y=53630
X4231 1 DigitalLDOLogic_VIA1 $T=158350 57940 0 0 $X=158100 $Y=57710
X4232 2 DigitalLDOLogic_VIA1 $T=160190 11700 0 0 $X=159940 $Y=11470
X4233 2 DigitalLDOLogic_VIA1 $T=160190 15780 0 0 $X=159940 $Y=15550
X4234 2 DigitalLDOLogic_VIA1 $T=160190 19860 0 0 $X=159940 $Y=19630
X4235 2 DigitalLDOLogic_VIA1 $T=160190 23940 0 0 $X=159940 $Y=23710
X4236 2 DigitalLDOLogic_VIA1 $T=160190 28020 0 0 $X=159940 $Y=27790
X4237 2 DigitalLDOLogic_VIA1 $T=160190 32100 0 0 $X=159940 $Y=31870
X4238 2 DigitalLDOLogic_VIA1 $T=160190 36180 0 0 $X=159940 $Y=35950
X4239 2 DigitalLDOLogic_VIA1 $T=160190 40260 0 0 $X=159940 $Y=40030
X4240 2 DigitalLDOLogic_VIA1 $T=160190 44340 0 0 $X=159940 $Y=44110
X4241 2 DigitalLDOLogic_VIA1 $T=160190 48420 0 0 $X=159940 $Y=48190
X4242 2 DigitalLDOLogic_VIA1 $T=160190 52500 0 0 $X=159940 $Y=52270
X4243 2 DigitalLDOLogic_VIA1 $T=160190 56580 0 0 $X=159940 $Y=56350
X4244 1 DigitalLDOLogic_VIA1 $T=161110 13060 0 0 $X=160860 $Y=12830
X4245 1 DigitalLDOLogic_VIA1 $T=161110 17140 0 0 $X=160860 $Y=16910
X4246 1 DigitalLDOLogic_VIA1 $T=161110 21220 0 0 $X=160860 $Y=20990
X4247 1 DigitalLDOLogic_VIA1 $T=161110 25300 0 0 $X=160860 $Y=25070
X4248 1 DigitalLDOLogic_VIA1 $T=161110 29380 0 0 $X=160860 $Y=29150
X4249 1 DigitalLDOLogic_VIA1 $T=161110 33460 0 0 $X=160860 $Y=33230
X4250 1 DigitalLDOLogic_VIA1 $T=161110 37540 0 0 $X=160860 $Y=37310
X4251 1 DigitalLDOLogic_VIA1 $T=161110 41620 0 0 $X=160860 $Y=41390
X4252 1 DigitalLDOLogic_VIA1 $T=161110 45700 0 0 $X=160860 $Y=45470
X4253 1 DigitalLDOLogic_VIA1 $T=161110 49780 0 0 $X=160860 $Y=49550
X4254 1 DigitalLDOLogic_VIA1 $T=161110 53860 0 0 $X=160860 $Y=53630
X4255 1 DigitalLDOLogic_VIA1 $T=161110 57940 0 0 $X=160860 $Y=57710
X4256 2 DigitalLDOLogic_VIA1 $T=162950 11700 0 0 $X=162700 $Y=11470
X4257 2 DigitalLDOLogic_VIA1 $T=162950 15780 0 0 $X=162700 $Y=15550
X4258 2 DigitalLDOLogic_VIA1 $T=162950 19860 0 0 $X=162700 $Y=19630
X4259 2 DigitalLDOLogic_VIA1 $T=162950 23940 0 0 $X=162700 $Y=23710
X4260 2 DigitalLDOLogic_VIA1 $T=162950 28020 0 0 $X=162700 $Y=27790
X4261 2 DigitalLDOLogic_VIA1 $T=162950 32100 0 0 $X=162700 $Y=31870
X4262 2 DigitalLDOLogic_VIA1 $T=162950 36180 0 0 $X=162700 $Y=35950
X4263 2 DigitalLDOLogic_VIA1 $T=162950 40260 0 0 $X=162700 $Y=40030
X4264 2 DigitalLDOLogic_VIA1 $T=162950 44340 0 0 $X=162700 $Y=44110
X4265 2 DigitalLDOLogic_VIA1 $T=162950 48420 0 0 $X=162700 $Y=48190
X4266 2 DigitalLDOLogic_VIA1 $T=162950 52500 0 0 $X=162700 $Y=52270
X4267 2 DigitalLDOLogic_VIA1 $T=162950 56580 0 0 $X=162700 $Y=56350
X4268 1 DigitalLDOLogic_VIA1 $T=163870 13060 0 0 $X=163620 $Y=12830
X4269 1 DigitalLDOLogic_VIA1 $T=163870 17140 0 0 $X=163620 $Y=16910
X4270 1 DigitalLDOLogic_VIA1 $T=163870 21220 0 0 $X=163620 $Y=20990
X4271 1 DigitalLDOLogic_VIA1 $T=163870 25300 0 0 $X=163620 $Y=25070
X4272 1 DigitalLDOLogic_VIA1 $T=163870 29380 0 0 $X=163620 $Y=29150
X4273 1 DigitalLDOLogic_VIA1 $T=163870 33460 0 0 $X=163620 $Y=33230
X4274 1 DigitalLDOLogic_VIA1 $T=163870 37540 0 0 $X=163620 $Y=37310
X4275 1 DigitalLDOLogic_VIA1 $T=163870 41620 0 0 $X=163620 $Y=41390
X4276 1 DigitalLDOLogic_VIA1 $T=163870 45700 0 0 $X=163620 $Y=45470
X4277 1 DigitalLDOLogic_VIA1 $T=163870 49780 0 0 $X=163620 $Y=49550
X4278 1 DigitalLDOLogic_VIA1 $T=163870 53860 0 0 $X=163620 $Y=53630
X4279 1 DigitalLDOLogic_VIA1 $T=163870 57940 0 0 $X=163620 $Y=57710
X4280 2 DigitalLDOLogic_VIA1 $T=165710 11700 0 0 $X=165460 $Y=11470
X4281 2 DigitalLDOLogic_VIA1 $T=165710 15780 0 0 $X=165460 $Y=15550
X4282 2 DigitalLDOLogic_VIA1 $T=165710 19860 0 0 $X=165460 $Y=19630
X4283 2 DigitalLDOLogic_VIA1 $T=165710 23940 0 0 $X=165460 $Y=23710
X4284 2 DigitalLDOLogic_VIA1 $T=165710 28020 0 0 $X=165460 $Y=27790
X4285 2 DigitalLDOLogic_VIA1 $T=165710 32100 0 0 $X=165460 $Y=31870
X4286 2 DigitalLDOLogic_VIA1 $T=165710 36180 0 0 $X=165460 $Y=35950
X4287 2 DigitalLDOLogic_VIA1 $T=165710 40260 0 0 $X=165460 $Y=40030
X4288 2 DigitalLDOLogic_VIA1 $T=165710 44340 0 0 $X=165460 $Y=44110
X4289 2 DigitalLDOLogic_VIA1 $T=165710 48420 0 0 $X=165460 $Y=48190
X4290 2 DigitalLDOLogic_VIA1 $T=165710 52500 0 0 $X=165460 $Y=52270
X4291 2 DigitalLDOLogic_VIA1 $T=165710 56580 0 0 $X=165460 $Y=56350
X4292 1 DigitalLDOLogic_VIA1 $T=166630 13060 0 0 $X=166380 $Y=12830
X4293 1 DigitalLDOLogic_VIA1 $T=166630 17140 0 0 $X=166380 $Y=16910
X4294 1 DigitalLDOLogic_VIA1 $T=166630 21220 0 0 $X=166380 $Y=20990
X4295 1 DigitalLDOLogic_VIA1 $T=166630 25300 0 0 $X=166380 $Y=25070
X4296 1 DigitalLDOLogic_VIA1 $T=166630 29380 0 0 $X=166380 $Y=29150
X4297 1 DigitalLDOLogic_VIA1 $T=166630 33460 0 0 $X=166380 $Y=33230
X4298 1 DigitalLDOLogic_VIA1 $T=166630 37540 0 0 $X=166380 $Y=37310
X4299 1 DigitalLDOLogic_VIA1 $T=166630 41620 0 0 $X=166380 $Y=41390
X4300 1 DigitalLDOLogic_VIA1 $T=166630 45700 0 0 $X=166380 $Y=45470
X4301 1 DigitalLDOLogic_VIA1 $T=166630 49780 0 0 $X=166380 $Y=49550
X4302 1 DigitalLDOLogic_VIA1 $T=166630 53860 0 0 $X=166380 $Y=53630
X4303 1 DigitalLDOLogic_VIA1 $T=166630 57940 0 0 $X=166380 $Y=57710
X4304 2 DigitalLDOLogic_VIA1 $T=168470 11700 0 0 $X=168220 $Y=11470
X4305 2 DigitalLDOLogic_VIA1 $T=168470 15780 0 0 $X=168220 $Y=15550
X4306 2 DigitalLDOLogic_VIA1 $T=168470 19860 0 0 $X=168220 $Y=19630
X4307 2 DigitalLDOLogic_VIA1 $T=168470 23940 0 0 $X=168220 $Y=23710
X4308 2 DigitalLDOLogic_VIA1 $T=168470 28020 0 0 $X=168220 $Y=27790
X4309 2 DigitalLDOLogic_VIA1 $T=168470 32100 0 0 $X=168220 $Y=31870
X4310 2 DigitalLDOLogic_VIA1 $T=168470 36180 0 0 $X=168220 $Y=35950
X4311 2 DigitalLDOLogic_VIA1 $T=168470 40260 0 0 $X=168220 $Y=40030
X4312 2 DigitalLDOLogic_VIA1 $T=168470 44340 0 0 $X=168220 $Y=44110
X4313 2 DigitalLDOLogic_VIA1 $T=168470 48420 0 0 $X=168220 $Y=48190
X4314 2 DigitalLDOLogic_VIA1 $T=168470 52500 0 0 $X=168220 $Y=52270
X4315 2 DigitalLDOLogic_VIA1 $T=168470 56580 0 0 $X=168220 $Y=56350
X4316 1 DigitalLDOLogic_VIA1 $T=169390 13060 0 0 $X=169140 $Y=12830
X4317 1 DigitalLDOLogic_VIA1 $T=169390 17140 0 0 $X=169140 $Y=16910
X4318 1 DigitalLDOLogic_VIA1 $T=169390 21220 0 0 $X=169140 $Y=20990
X4319 1 DigitalLDOLogic_VIA1 $T=169390 25300 0 0 $X=169140 $Y=25070
X4320 1 DigitalLDOLogic_VIA1 $T=169390 29380 0 0 $X=169140 $Y=29150
X4321 1 DigitalLDOLogic_VIA1 $T=169390 33460 0 0 $X=169140 $Y=33230
X4322 1 DigitalLDOLogic_VIA1 $T=169390 37540 0 0 $X=169140 $Y=37310
X4323 1 DigitalLDOLogic_VIA1 $T=169390 41620 0 0 $X=169140 $Y=41390
X4324 1 DigitalLDOLogic_VIA1 $T=169390 45700 0 0 $X=169140 $Y=45470
X4325 1 DigitalLDOLogic_VIA1 $T=169390 49780 0 0 $X=169140 $Y=49550
X4326 1 DigitalLDOLogic_VIA1 $T=169390 53860 0 0 $X=169140 $Y=53630
X4327 1 DigitalLDOLogic_VIA1 $T=169390 57940 0 0 $X=169140 $Y=57710
X4328 2 DigitalLDOLogic_VIA1 $T=171230 11700 0 0 $X=170980 $Y=11470
X4329 2 DigitalLDOLogic_VIA1 $T=171230 15780 0 0 $X=170980 $Y=15550
X4330 2 DigitalLDOLogic_VIA1 $T=171230 19860 0 0 $X=170980 $Y=19630
X4331 2 DigitalLDOLogic_VIA1 $T=171230 23940 0 0 $X=170980 $Y=23710
X4332 2 DigitalLDOLogic_VIA1 $T=171230 28020 0 0 $X=170980 $Y=27790
X4333 2 DigitalLDOLogic_VIA1 $T=171230 32100 0 0 $X=170980 $Y=31870
X4334 2 DigitalLDOLogic_VIA1 $T=171230 36180 0 0 $X=170980 $Y=35950
X4335 2 DigitalLDOLogic_VIA1 $T=171230 40260 0 0 $X=170980 $Y=40030
X4336 2 DigitalLDOLogic_VIA1 $T=171230 44340 0 0 $X=170980 $Y=44110
X4337 2 DigitalLDOLogic_VIA1 $T=171230 48420 0 0 $X=170980 $Y=48190
X4338 2 DigitalLDOLogic_VIA1 $T=171230 52500 0 0 $X=170980 $Y=52270
X4339 2 DigitalLDOLogic_VIA1 $T=171230 56580 0 0 $X=170980 $Y=56350
X4340 1 DigitalLDOLogic_VIA1 $T=172150 13060 0 0 $X=171900 $Y=12830
X4341 1 DigitalLDOLogic_VIA1 $T=172150 17140 0 0 $X=171900 $Y=16910
X4342 1 DigitalLDOLogic_VIA1 $T=172150 21220 0 0 $X=171900 $Y=20990
X4343 1 DigitalLDOLogic_VIA1 $T=172150 25300 0 0 $X=171900 $Y=25070
X4344 1 DigitalLDOLogic_VIA1 $T=172150 29380 0 0 $X=171900 $Y=29150
X4345 1 DigitalLDOLogic_VIA1 $T=172150 33460 0 0 $X=171900 $Y=33230
X4346 1 DigitalLDOLogic_VIA1 $T=172150 37540 0 0 $X=171900 $Y=37310
X4347 1 DigitalLDOLogic_VIA1 $T=172150 41620 0 0 $X=171900 $Y=41390
X4348 1 DigitalLDOLogic_VIA1 $T=172150 45700 0 0 $X=171900 $Y=45470
X4349 1 DigitalLDOLogic_VIA1 $T=172150 49780 0 0 $X=171900 $Y=49550
X4350 1 DigitalLDOLogic_VIA1 $T=172150 53860 0 0 $X=171900 $Y=53630
X4351 1 DigitalLDOLogic_VIA1 $T=172150 57940 0 0 $X=171900 $Y=57710
X4352 2 DigitalLDOLogic_VIA1 $T=173990 11700 0 0 $X=173740 $Y=11470
X4353 2 DigitalLDOLogic_VIA1 $T=173990 15780 0 0 $X=173740 $Y=15550
X4354 2 DigitalLDOLogic_VIA1 $T=173990 19860 0 0 $X=173740 $Y=19630
X4355 2 DigitalLDOLogic_VIA1 $T=173990 23940 0 0 $X=173740 $Y=23710
X4356 2 DigitalLDOLogic_VIA1 $T=173990 28020 0 0 $X=173740 $Y=27790
X4357 2 DigitalLDOLogic_VIA1 $T=173990 32100 0 0 $X=173740 $Y=31870
X4358 2 DigitalLDOLogic_VIA1 $T=173990 36180 0 0 $X=173740 $Y=35950
X4359 2 DigitalLDOLogic_VIA1 $T=173990 40260 0 0 $X=173740 $Y=40030
X4360 2 DigitalLDOLogic_VIA1 $T=173990 44340 0 0 $X=173740 $Y=44110
X4361 2 DigitalLDOLogic_VIA1 $T=173990 48420 0 0 $X=173740 $Y=48190
X4362 2 DigitalLDOLogic_VIA1 $T=173990 52500 0 0 $X=173740 $Y=52270
X4363 2 DigitalLDOLogic_VIA1 $T=173990 56580 0 0 $X=173740 $Y=56350
X4364 1 DigitalLDOLogic_VIA1 $T=174910 13060 0 0 $X=174660 $Y=12830
X4365 1 DigitalLDOLogic_VIA1 $T=174910 17140 0 0 $X=174660 $Y=16910
X4366 1 DigitalLDOLogic_VIA1 $T=174910 21220 0 0 $X=174660 $Y=20990
X4367 1 DigitalLDOLogic_VIA1 $T=174910 25300 0 0 $X=174660 $Y=25070
X4368 1 DigitalLDOLogic_VIA1 $T=174910 29380 0 0 $X=174660 $Y=29150
X4369 1 DigitalLDOLogic_VIA1 $T=174910 33460 0 0 $X=174660 $Y=33230
X4370 1 DigitalLDOLogic_VIA1 $T=174910 37540 0 0 $X=174660 $Y=37310
X4371 1 DigitalLDOLogic_VIA1 $T=174910 41620 0 0 $X=174660 $Y=41390
X4372 1 DigitalLDOLogic_VIA1 $T=174910 45700 0 0 $X=174660 $Y=45470
X4373 1 DigitalLDOLogic_VIA1 $T=174910 49780 0 0 $X=174660 $Y=49550
X4374 1 DigitalLDOLogic_VIA1 $T=174910 53860 0 0 $X=174660 $Y=53630
X4375 1 DigitalLDOLogic_VIA1 $T=174910 57940 0 0 $X=174660 $Y=57710
X4376 2 DigitalLDOLogic_VIA1 $T=176750 11700 0 0 $X=176500 $Y=11470
X4377 2 DigitalLDOLogic_VIA1 $T=176750 15780 0 0 $X=176500 $Y=15550
X4378 2 DigitalLDOLogic_VIA1 $T=176750 19860 0 0 $X=176500 $Y=19630
X4379 2 DigitalLDOLogic_VIA1 $T=176750 23940 0 0 $X=176500 $Y=23710
X4380 2 DigitalLDOLogic_VIA1 $T=176750 28020 0 0 $X=176500 $Y=27790
X4381 2 DigitalLDOLogic_VIA1 $T=176750 32100 0 0 $X=176500 $Y=31870
X4382 2 DigitalLDOLogic_VIA1 $T=176750 36180 0 0 $X=176500 $Y=35950
X4383 2 DigitalLDOLogic_VIA1 $T=176750 40260 0 0 $X=176500 $Y=40030
X4384 2 DigitalLDOLogic_VIA1 $T=176750 44340 0 0 $X=176500 $Y=44110
X4385 2 DigitalLDOLogic_VIA1 $T=176750 48420 0 0 $X=176500 $Y=48190
X4386 2 DigitalLDOLogic_VIA1 $T=176750 52500 0 0 $X=176500 $Y=52270
X4387 2 DigitalLDOLogic_VIA1 $T=176750 56580 0 0 $X=176500 $Y=56350
X4388 1 DigitalLDOLogic_VIA1 $T=177670 13060 0 0 $X=177420 $Y=12830
X4389 1 DigitalLDOLogic_VIA1 $T=177670 17140 0 0 $X=177420 $Y=16910
X4390 1 DigitalLDOLogic_VIA1 $T=177670 21220 0 0 $X=177420 $Y=20990
X4391 1 DigitalLDOLogic_VIA1 $T=177670 25300 0 0 $X=177420 $Y=25070
X4392 1 DigitalLDOLogic_VIA1 $T=177670 29380 0 0 $X=177420 $Y=29150
X4393 1 DigitalLDOLogic_VIA1 $T=177670 33460 0 0 $X=177420 $Y=33230
X4394 1 DigitalLDOLogic_VIA1 $T=177670 37540 0 0 $X=177420 $Y=37310
X4395 1 DigitalLDOLogic_VIA1 $T=177670 41620 0 0 $X=177420 $Y=41390
X4396 1 DigitalLDOLogic_VIA1 $T=177670 45700 0 0 $X=177420 $Y=45470
X4397 1 DigitalLDOLogic_VIA1 $T=177670 49780 0 0 $X=177420 $Y=49550
X4398 1 DigitalLDOLogic_VIA1 $T=177670 53860 0 0 $X=177420 $Y=53630
X4399 1 DigitalLDOLogic_VIA1 $T=177670 57940 0 0 $X=177420 $Y=57710
X4400 2 DigitalLDOLogic_VIA1 $T=179510 11700 0 0 $X=179260 $Y=11470
X4401 2 DigitalLDOLogic_VIA1 $T=179510 15780 0 0 $X=179260 $Y=15550
X4402 2 DigitalLDOLogic_VIA1 $T=179510 19860 0 0 $X=179260 $Y=19630
X4403 2 DigitalLDOLogic_VIA1 $T=179510 23940 0 0 $X=179260 $Y=23710
X4404 2 DigitalLDOLogic_VIA1 $T=179510 28020 0 0 $X=179260 $Y=27790
X4405 2 DigitalLDOLogic_VIA1 $T=179510 32100 0 0 $X=179260 $Y=31870
X4406 2 DigitalLDOLogic_VIA1 $T=179510 36180 0 0 $X=179260 $Y=35950
X4407 2 DigitalLDOLogic_VIA1 $T=179510 40260 0 0 $X=179260 $Y=40030
X4408 2 DigitalLDOLogic_VIA1 $T=179510 44340 0 0 $X=179260 $Y=44110
X4409 2 DigitalLDOLogic_VIA1 $T=179510 48420 0 0 $X=179260 $Y=48190
X4410 2 DigitalLDOLogic_VIA1 $T=179510 52500 0 0 $X=179260 $Y=52270
X4411 2 DigitalLDOLogic_VIA1 $T=179510 56580 0 0 $X=179260 $Y=56350
X4412 1 DigitalLDOLogic_VIA1 $T=180430 13060 0 0 $X=180180 $Y=12830
X4413 1 DigitalLDOLogic_VIA1 $T=180430 17140 0 0 $X=180180 $Y=16910
X4414 1 DigitalLDOLogic_VIA1 $T=180430 21220 0 0 $X=180180 $Y=20990
X4415 1 DigitalLDOLogic_VIA1 $T=180430 25300 0 0 $X=180180 $Y=25070
X4416 1 DigitalLDOLogic_VIA1 $T=180430 29380 0 0 $X=180180 $Y=29150
X4417 1 DigitalLDOLogic_VIA1 $T=180430 33460 0 0 $X=180180 $Y=33230
X4418 1 DigitalLDOLogic_VIA1 $T=180430 37540 0 0 $X=180180 $Y=37310
X4419 1 DigitalLDOLogic_VIA1 $T=180430 41620 0 0 $X=180180 $Y=41390
X4420 1 DigitalLDOLogic_VIA1 $T=180430 45700 0 0 $X=180180 $Y=45470
X4421 1 DigitalLDOLogic_VIA1 $T=180430 49780 0 0 $X=180180 $Y=49550
X4422 1 DigitalLDOLogic_VIA1 $T=180430 53860 0 0 $X=180180 $Y=53630
X4423 1 DigitalLDOLogic_VIA1 $T=180430 57940 0 0 $X=180180 $Y=57710
X4424 2 DigitalLDOLogic_VIA1 $T=182270 11700 0 0 $X=182020 $Y=11470
X4425 2 DigitalLDOLogic_VIA1 $T=182270 15780 0 0 $X=182020 $Y=15550
X4426 2 DigitalLDOLogic_VIA1 $T=182270 19860 0 0 $X=182020 $Y=19630
X4427 2 DigitalLDOLogic_VIA1 $T=182270 23940 0 0 $X=182020 $Y=23710
X4428 2 DigitalLDOLogic_VIA1 $T=182270 28020 0 0 $X=182020 $Y=27790
X4429 2 DigitalLDOLogic_VIA1 $T=182270 32100 0 0 $X=182020 $Y=31870
X4430 2 DigitalLDOLogic_VIA1 $T=182270 36180 0 0 $X=182020 $Y=35950
X4431 2 DigitalLDOLogic_VIA1 $T=182270 40260 0 0 $X=182020 $Y=40030
X4432 2 DigitalLDOLogic_VIA1 $T=182270 44340 0 0 $X=182020 $Y=44110
X4433 2 DigitalLDOLogic_VIA1 $T=182270 48420 0 0 $X=182020 $Y=48190
X4434 2 DigitalLDOLogic_VIA1 $T=182270 52500 0 0 $X=182020 $Y=52270
X4435 2 DigitalLDOLogic_VIA1 $T=182270 56580 0 0 $X=182020 $Y=56350
X4436 1 DigitalLDOLogic_VIA1 $T=183190 13060 0 0 $X=182940 $Y=12830
X4437 1 DigitalLDOLogic_VIA1 $T=183190 17140 0 0 $X=182940 $Y=16910
X4438 1 DigitalLDOLogic_VIA1 $T=183190 21220 0 0 $X=182940 $Y=20990
X4439 1 DigitalLDOLogic_VIA1 $T=183190 25300 0 0 $X=182940 $Y=25070
X4440 1 DigitalLDOLogic_VIA1 $T=183190 29380 0 0 $X=182940 $Y=29150
X4441 1 DigitalLDOLogic_VIA1 $T=183190 33460 0 0 $X=182940 $Y=33230
X4442 1 DigitalLDOLogic_VIA1 $T=183190 37540 0 0 $X=182940 $Y=37310
X4443 1 DigitalLDOLogic_VIA1 $T=183190 41620 0 0 $X=182940 $Y=41390
X4444 1 DigitalLDOLogic_VIA1 $T=183190 45700 0 0 $X=182940 $Y=45470
X4445 1 DigitalLDOLogic_VIA1 $T=183190 49780 0 0 $X=182940 $Y=49550
X4446 1 DigitalLDOLogic_VIA1 $T=183190 53860 0 0 $X=182940 $Y=53630
X4447 1 DigitalLDOLogic_VIA1 $T=183190 57940 0 0 $X=182940 $Y=57710
X4448 2 DigitalLDOLogic_VIA1 $T=185030 11700 0 0 $X=184780 $Y=11470
X4449 2 DigitalLDOLogic_VIA1 $T=185030 15780 0 0 $X=184780 $Y=15550
X4450 2 DigitalLDOLogic_VIA1 $T=185030 19860 0 0 $X=184780 $Y=19630
X4451 2 DigitalLDOLogic_VIA1 $T=185030 23940 0 0 $X=184780 $Y=23710
X4452 2 DigitalLDOLogic_VIA1 $T=185030 28020 0 0 $X=184780 $Y=27790
X4453 2 DigitalLDOLogic_VIA1 $T=185030 32100 0 0 $X=184780 $Y=31870
X4454 2 DigitalLDOLogic_VIA1 $T=185030 36180 0 0 $X=184780 $Y=35950
X4455 2 DigitalLDOLogic_VIA1 $T=185030 40260 0 0 $X=184780 $Y=40030
X4456 2 DigitalLDOLogic_VIA1 $T=185030 44340 0 0 $X=184780 $Y=44110
X4457 2 DigitalLDOLogic_VIA1 $T=185030 48420 0 0 $X=184780 $Y=48190
X4458 2 DigitalLDOLogic_VIA1 $T=185030 52500 0 0 $X=184780 $Y=52270
X4459 2 DigitalLDOLogic_VIA1 $T=185030 56580 0 0 $X=184780 $Y=56350
X4460 1 DigitalLDOLogic_VIA1 $T=185950 13060 0 0 $X=185700 $Y=12830
X4461 1 DigitalLDOLogic_VIA1 $T=185950 17140 0 0 $X=185700 $Y=16910
X4462 1 DigitalLDOLogic_VIA1 $T=185950 21220 0 0 $X=185700 $Y=20990
X4463 1 DigitalLDOLogic_VIA1 $T=185950 25300 0 0 $X=185700 $Y=25070
X4464 1 DigitalLDOLogic_VIA1 $T=185950 29380 0 0 $X=185700 $Y=29150
X4465 1 DigitalLDOLogic_VIA1 $T=185950 33460 0 0 $X=185700 $Y=33230
X4466 1 DigitalLDOLogic_VIA1 $T=185950 37540 0 0 $X=185700 $Y=37310
X4467 1 DigitalLDOLogic_VIA1 $T=185950 41620 0 0 $X=185700 $Y=41390
X4468 1 DigitalLDOLogic_VIA1 $T=185950 45700 0 0 $X=185700 $Y=45470
X4469 1 DigitalLDOLogic_VIA1 $T=185950 49780 0 0 $X=185700 $Y=49550
X4470 1 DigitalLDOLogic_VIA1 $T=185950 53860 0 0 $X=185700 $Y=53630
X4471 1 DigitalLDOLogic_VIA1 $T=185950 57940 0 0 $X=185700 $Y=57710
X4472 2 DigitalLDOLogic_VIA1 $T=187790 11700 0 0 $X=187540 $Y=11470
X4473 2 DigitalLDOLogic_VIA1 $T=187790 15780 0 0 $X=187540 $Y=15550
X4474 2 DigitalLDOLogic_VIA1 $T=187790 19860 0 0 $X=187540 $Y=19630
X4475 2 DigitalLDOLogic_VIA1 $T=187790 23940 0 0 $X=187540 $Y=23710
X4476 2 DigitalLDOLogic_VIA1 $T=187790 28020 0 0 $X=187540 $Y=27790
X4477 2 DigitalLDOLogic_VIA1 $T=187790 32100 0 0 $X=187540 $Y=31870
X4478 2 DigitalLDOLogic_VIA1 $T=187790 36180 0 0 $X=187540 $Y=35950
X4479 2 DigitalLDOLogic_VIA1 $T=187790 40260 0 0 $X=187540 $Y=40030
X4480 2 DigitalLDOLogic_VIA1 $T=187790 44340 0 0 $X=187540 $Y=44110
X4481 2 DigitalLDOLogic_VIA1 $T=187790 48420 0 0 $X=187540 $Y=48190
X4482 2 DigitalLDOLogic_VIA1 $T=187790 52500 0 0 $X=187540 $Y=52270
X4483 2 DigitalLDOLogic_VIA1 $T=187790 56580 0 0 $X=187540 $Y=56350
X4484 1 DigitalLDOLogic_VIA1 $T=188710 13060 0 0 $X=188460 $Y=12830
X4485 1 DigitalLDOLogic_VIA1 $T=188710 17140 0 0 $X=188460 $Y=16910
X4486 1 DigitalLDOLogic_VIA1 $T=188710 21220 0 0 $X=188460 $Y=20990
X4487 1 DigitalLDOLogic_VIA1 $T=188710 25300 0 0 $X=188460 $Y=25070
X4488 1 DigitalLDOLogic_VIA1 $T=188710 29380 0 0 $X=188460 $Y=29150
X4489 1 DigitalLDOLogic_VIA1 $T=188710 33460 0 0 $X=188460 $Y=33230
X4490 1 DigitalLDOLogic_VIA1 $T=188710 37540 0 0 $X=188460 $Y=37310
X4491 1 DigitalLDOLogic_VIA1 $T=188710 41620 0 0 $X=188460 $Y=41390
X4492 1 DigitalLDOLogic_VIA1 $T=188710 45700 0 0 $X=188460 $Y=45470
X4493 1 DigitalLDOLogic_VIA1 $T=188710 49780 0 0 $X=188460 $Y=49550
X4494 1 DigitalLDOLogic_VIA1 $T=188710 53860 0 0 $X=188460 $Y=53630
X4495 1 DigitalLDOLogic_VIA1 $T=188710 57940 0 0 $X=188460 $Y=57710
X4496 2 DigitalLDOLogic_VIA2 $T=12300 11700 0 0 $X=11830 $Y=11470
X4497 2 DigitalLDOLogic_VIA2 $T=12300 15780 0 0 $X=11830 $Y=15550
X4498 2 DigitalLDOLogic_VIA2 $T=12300 19860 0 0 $X=11830 $Y=19630
X4499 2 DigitalLDOLogic_VIA2 $T=12300 23940 0 0 $X=11830 $Y=23710
X4500 2 DigitalLDOLogic_VIA2 $T=12300 28020 0 0 $X=11830 $Y=27790
X4501 2 DigitalLDOLogic_VIA2 $T=12300 32100 0 0 $X=11830 $Y=31870
X4502 2 DigitalLDOLogic_VIA2 $T=12300 36180 0 0 $X=11830 $Y=35950
X4503 2 DigitalLDOLogic_VIA2 $T=12300 40260 0 0 $X=11830 $Y=40030
X4504 2 DigitalLDOLogic_VIA2 $T=12300 44340 0 0 $X=11830 $Y=44110
X4505 2 DigitalLDOLogic_VIA2 $T=12300 48420 0 0 $X=11830 $Y=48190
X4506 2 DigitalLDOLogic_VIA2 $T=12300 52500 0 0 $X=11830 $Y=52270
X4507 2 DigitalLDOLogic_VIA2 $T=12300 56580 0 0 $X=11830 $Y=56350
X4508 1 DigitalLDOLogic_VIA2 $T=14140 13060 0 0 $X=13670 $Y=12830
X4509 1 DigitalLDOLogic_VIA2 $T=14140 17140 0 0 $X=13670 $Y=16910
X4510 1 DigitalLDOLogic_VIA2 $T=14140 21220 0 0 $X=13670 $Y=20990
X4511 1 DigitalLDOLogic_VIA2 $T=14140 25300 0 0 $X=13670 $Y=25070
X4512 1 DigitalLDOLogic_VIA2 $T=14140 29380 0 0 $X=13670 $Y=29150
X4513 1 DigitalLDOLogic_VIA2 $T=14140 33460 0 0 $X=13670 $Y=33230
X4514 1 DigitalLDOLogic_VIA2 $T=14140 37540 0 0 $X=13670 $Y=37310
X4515 1 DigitalLDOLogic_VIA2 $T=14140 41620 0 0 $X=13670 $Y=41390
X4516 1 DigitalLDOLogic_VIA2 $T=14140 45700 0 0 $X=13670 $Y=45470
X4517 1 DigitalLDOLogic_VIA2 $T=14140 49780 0 0 $X=13670 $Y=49550
X4518 1 DigitalLDOLogic_VIA2 $T=14140 53860 0 0 $X=13670 $Y=53630
X4519 1 DigitalLDOLogic_VIA2 $T=14140 57940 0 0 $X=13670 $Y=57710
X4520 2 DigitalLDOLogic_VIA2 $T=17820 11700 0 0 $X=17350 $Y=11470
X4521 2 DigitalLDOLogic_VIA2 $T=17820 15780 0 0 $X=17350 $Y=15550
X4522 2 DigitalLDOLogic_VIA2 $T=17820 19860 0 0 $X=17350 $Y=19630
X4523 2 DigitalLDOLogic_VIA2 $T=17820 23940 0 0 $X=17350 $Y=23710
X4524 2 DigitalLDOLogic_VIA2 $T=17820 28020 0 0 $X=17350 $Y=27790
X4525 2 DigitalLDOLogic_VIA2 $T=17820 32100 0 0 $X=17350 $Y=31870
X4526 2 DigitalLDOLogic_VIA2 $T=17820 36180 0 0 $X=17350 $Y=35950
X4527 2 DigitalLDOLogic_VIA2 $T=17820 40260 0 0 $X=17350 $Y=40030
X4528 2 DigitalLDOLogic_VIA2 $T=17820 44340 0 0 $X=17350 $Y=44110
X4529 2 DigitalLDOLogic_VIA2 $T=17820 48420 0 0 $X=17350 $Y=48190
X4530 2 DigitalLDOLogic_VIA2 $T=17820 52500 0 0 $X=17350 $Y=52270
X4531 2 DigitalLDOLogic_VIA2 $T=17820 56580 0 0 $X=17350 $Y=56350
X4532 1 DigitalLDOLogic_VIA2 $T=19660 13060 0 0 $X=19190 $Y=12830
X4533 1 DigitalLDOLogic_VIA2 $T=19660 17140 0 0 $X=19190 $Y=16910
X4534 1 DigitalLDOLogic_VIA2 $T=19660 21220 0 0 $X=19190 $Y=20990
X4535 1 DigitalLDOLogic_VIA2 $T=19660 25300 0 0 $X=19190 $Y=25070
X4536 1 DigitalLDOLogic_VIA2 $T=19660 29380 0 0 $X=19190 $Y=29150
X4537 1 DigitalLDOLogic_VIA2 $T=19660 33460 0 0 $X=19190 $Y=33230
X4538 1 DigitalLDOLogic_VIA2 $T=19660 37540 0 0 $X=19190 $Y=37310
X4539 1 DigitalLDOLogic_VIA2 $T=19660 41620 0 0 $X=19190 $Y=41390
X4540 1 DigitalLDOLogic_VIA2 $T=19660 45700 0 0 $X=19190 $Y=45470
X4541 1 DigitalLDOLogic_VIA2 $T=19660 49780 0 0 $X=19190 $Y=49550
X4542 1 DigitalLDOLogic_VIA2 $T=19660 53860 0 0 $X=19190 $Y=53630
X4543 1 DigitalLDOLogic_VIA2 $T=19660 57940 0 0 $X=19190 $Y=57710
X4544 2 DigitalLDOLogic_VIA2 $T=23340 11700 0 0 $X=22870 $Y=11470
X4545 2 DigitalLDOLogic_VIA2 $T=23340 15780 0 0 $X=22870 $Y=15550
X4546 2 DigitalLDOLogic_VIA2 $T=23340 19860 0 0 $X=22870 $Y=19630
X4547 2 DigitalLDOLogic_VIA2 $T=23340 23940 0 0 $X=22870 $Y=23710
X4548 2 DigitalLDOLogic_VIA2 $T=23340 28020 0 0 $X=22870 $Y=27790
X4549 2 DigitalLDOLogic_VIA2 $T=23340 32100 0 0 $X=22870 $Y=31870
X4550 2 DigitalLDOLogic_VIA2 $T=23340 36180 0 0 $X=22870 $Y=35950
X4551 2 DigitalLDOLogic_VIA2 $T=23340 40260 0 0 $X=22870 $Y=40030
X4552 2 DigitalLDOLogic_VIA2 $T=23340 44340 0 0 $X=22870 $Y=44110
X4553 2 DigitalLDOLogic_VIA2 $T=23340 48420 0 0 $X=22870 $Y=48190
X4554 2 DigitalLDOLogic_VIA2 $T=23340 52500 0 0 $X=22870 $Y=52270
X4555 2 DigitalLDOLogic_VIA2 $T=23340 56580 0 0 $X=22870 $Y=56350
X4556 1 DigitalLDOLogic_VIA2 $T=25180 13060 0 0 $X=24710 $Y=12830
X4557 1 DigitalLDOLogic_VIA2 $T=25180 17140 0 0 $X=24710 $Y=16910
X4558 1 DigitalLDOLogic_VIA2 $T=25180 21220 0 0 $X=24710 $Y=20990
X4559 1 DigitalLDOLogic_VIA2 $T=25180 25300 0 0 $X=24710 $Y=25070
X4560 1 DigitalLDOLogic_VIA2 $T=25180 29380 0 0 $X=24710 $Y=29150
X4561 1 DigitalLDOLogic_VIA2 $T=25180 33460 0 0 $X=24710 $Y=33230
X4562 1 DigitalLDOLogic_VIA2 $T=25180 37540 0 0 $X=24710 $Y=37310
X4563 1 DigitalLDOLogic_VIA2 $T=25180 41620 0 0 $X=24710 $Y=41390
X4564 1 DigitalLDOLogic_VIA2 $T=25180 45700 0 0 $X=24710 $Y=45470
X4565 1 DigitalLDOLogic_VIA2 $T=25180 49780 0 0 $X=24710 $Y=49550
X4566 1 DigitalLDOLogic_VIA2 $T=25180 53860 0 0 $X=24710 $Y=53630
X4567 1 DigitalLDOLogic_VIA2 $T=25180 57940 0 0 $X=24710 $Y=57710
X4568 2 DigitalLDOLogic_VIA2 $T=28860 11700 0 0 $X=28390 $Y=11470
X4569 2 DigitalLDOLogic_VIA2 $T=28860 15780 0 0 $X=28390 $Y=15550
X4570 2 DigitalLDOLogic_VIA2 $T=28860 19860 0 0 $X=28390 $Y=19630
X4571 2 DigitalLDOLogic_VIA2 $T=28860 23940 0 0 $X=28390 $Y=23710
X4572 2 DigitalLDOLogic_VIA2 $T=28860 28020 0 0 $X=28390 $Y=27790
X4573 2 DigitalLDOLogic_VIA2 $T=28860 32100 0 0 $X=28390 $Y=31870
X4574 2 DigitalLDOLogic_VIA2 $T=28860 36180 0 0 $X=28390 $Y=35950
X4575 2 DigitalLDOLogic_VIA2 $T=28860 40260 0 0 $X=28390 $Y=40030
X4576 2 DigitalLDOLogic_VIA2 $T=28860 44340 0 0 $X=28390 $Y=44110
X4577 2 DigitalLDOLogic_VIA2 $T=28860 48420 0 0 $X=28390 $Y=48190
X4578 2 DigitalLDOLogic_VIA2 $T=28860 52500 0 0 $X=28390 $Y=52270
X4579 2 DigitalLDOLogic_VIA2 $T=28860 56580 0 0 $X=28390 $Y=56350
X4580 1 DigitalLDOLogic_VIA2 $T=30700 13060 0 0 $X=30230 $Y=12830
X4581 1 DigitalLDOLogic_VIA2 $T=30700 17140 0 0 $X=30230 $Y=16910
X4582 1 DigitalLDOLogic_VIA2 $T=30700 21220 0 0 $X=30230 $Y=20990
X4583 1 DigitalLDOLogic_VIA2 $T=30700 25300 0 0 $X=30230 $Y=25070
X4584 1 DigitalLDOLogic_VIA2 $T=30700 29380 0 0 $X=30230 $Y=29150
X4585 1 DigitalLDOLogic_VIA2 $T=30700 33460 0 0 $X=30230 $Y=33230
X4586 1 DigitalLDOLogic_VIA2 $T=30700 37540 0 0 $X=30230 $Y=37310
X4587 1 DigitalLDOLogic_VIA2 $T=30700 41620 0 0 $X=30230 $Y=41390
X4588 1 DigitalLDOLogic_VIA2 $T=30700 45700 0 0 $X=30230 $Y=45470
X4589 1 DigitalLDOLogic_VIA2 $T=30700 49780 0 0 $X=30230 $Y=49550
X4590 1 DigitalLDOLogic_VIA2 $T=30700 53860 0 0 $X=30230 $Y=53630
X4591 1 DigitalLDOLogic_VIA2 $T=30700 57940 0 0 $X=30230 $Y=57710
X4592 2 DigitalLDOLogic_VIA2 $T=34380 11700 0 0 $X=33910 $Y=11470
X4593 2 DigitalLDOLogic_VIA2 $T=34380 15780 0 0 $X=33910 $Y=15550
X4594 2 DigitalLDOLogic_VIA2 $T=34380 19860 0 0 $X=33910 $Y=19630
X4595 2 DigitalLDOLogic_VIA2 $T=34380 23940 0 0 $X=33910 $Y=23710
X4596 2 DigitalLDOLogic_VIA2 $T=34380 28020 0 0 $X=33910 $Y=27790
X4597 2 DigitalLDOLogic_VIA2 $T=34380 32100 0 0 $X=33910 $Y=31870
X4598 2 DigitalLDOLogic_VIA2 $T=34380 36180 0 0 $X=33910 $Y=35950
X4599 2 DigitalLDOLogic_VIA2 $T=34380 40260 0 0 $X=33910 $Y=40030
X4600 2 DigitalLDOLogic_VIA2 $T=34380 44340 0 0 $X=33910 $Y=44110
X4601 2 DigitalLDOLogic_VIA2 $T=34380 48420 0 0 $X=33910 $Y=48190
X4602 2 DigitalLDOLogic_VIA2 $T=34380 52500 0 0 $X=33910 $Y=52270
X4603 2 DigitalLDOLogic_VIA2 $T=34380 56580 0 0 $X=33910 $Y=56350
X4604 1 DigitalLDOLogic_VIA2 $T=36220 13060 0 0 $X=35750 $Y=12830
X4605 1 DigitalLDOLogic_VIA2 $T=36220 17140 0 0 $X=35750 $Y=16910
X4606 1 DigitalLDOLogic_VIA2 $T=36220 21220 0 0 $X=35750 $Y=20990
X4607 1 DigitalLDOLogic_VIA2 $T=36220 25300 0 0 $X=35750 $Y=25070
X4608 1 DigitalLDOLogic_VIA2 $T=36220 29380 0 0 $X=35750 $Y=29150
X4609 1 DigitalLDOLogic_VIA2 $T=36220 33460 0 0 $X=35750 $Y=33230
X4610 1 DigitalLDOLogic_VIA2 $T=36220 37540 0 0 $X=35750 $Y=37310
X4611 1 DigitalLDOLogic_VIA2 $T=36220 41620 0 0 $X=35750 $Y=41390
X4612 1 DigitalLDOLogic_VIA2 $T=36220 45700 0 0 $X=35750 $Y=45470
X4613 1 DigitalLDOLogic_VIA2 $T=36220 49780 0 0 $X=35750 $Y=49550
X4614 1 DigitalLDOLogic_VIA2 $T=36220 53860 0 0 $X=35750 $Y=53630
X4615 1 DigitalLDOLogic_VIA2 $T=36220 57940 0 0 $X=35750 $Y=57710
X4616 2 DigitalLDOLogic_VIA2 $T=39900 11700 0 0 $X=39430 $Y=11470
X4617 2 DigitalLDOLogic_VIA2 $T=39900 15780 0 0 $X=39430 $Y=15550
X4618 2 DigitalLDOLogic_VIA2 $T=39900 19860 0 0 $X=39430 $Y=19630
X4619 2 DigitalLDOLogic_VIA2 $T=39900 23940 0 0 $X=39430 $Y=23710
X4620 2 DigitalLDOLogic_VIA2 $T=39900 28020 0 0 $X=39430 $Y=27790
X4621 2 DigitalLDOLogic_VIA2 $T=39900 32100 0 0 $X=39430 $Y=31870
X4622 2 DigitalLDOLogic_VIA2 $T=39900 36180 0 0 $X=39430 $Y=35950
X4623 2 DigitalLDOLogic_VIA2 $T=39900 40260 0 0 $X=39430 $Y=40030
X4624 2 DigitalLDOLogic_VIA2 $T=39900 44340 0 0 $X=39430 $Y=44110
X4625 2 DigitalLDOLogic_VIA2 $T=39900 48420 0 0 $X=39430 $Y=48190
X4626 2 DigitalLDOLogic_VIA2 $T=39900 52500 0 0 $X=39430 $Y=52270
X4627 2 DigitalLDOLogic_VIA2 $T=39900 56580 0 0 $X=39430 $Y=56350
X4628 1 DigitalLDOLogic_VIA2 $T=41740 13060 0 0 $X=41270 $Y=12830
X4629 1 DigitalLDOLogic_VIA2 $T=41740 17140 0 0 $X=41270 $Y=16910
X4630 1 DigitalLDOLogic_VIA2 $T=41740 21220 0 0 $X=41270 $Y=20990
X4631 1 DigitalLDOLogic_VIA2 $T=41740 25300 0 0 $X=41270 $Y=25070
X4632 1 DigitalLDOLogic_VIA2 $T=41740 29380 0 0 $X=41270 $Y=29150
X4633 1 DigitalLDOLogic_VIA2 $T=41740 33460 0 0 $X=41270 $Y=33230
X4634 1 DigitalLDOLogic_VIA2 $T=41740 37540 0 0 $X=41270 $Y=37310
X4635 1 DigitalLDOLogic_VIA2 $T=41740 41620 0 0 $X=41270 $Y=41390
X4636 1 DigitalLDOLogic_VIA2 $T=41740 45700 0 0 $X=41270 $Y=45470
X4637 1 DigitalLDOLogic_VIA2 $T=41740 49780 0 0 $X=41270 $Y=49550
X4638 1 DigitalLDOLogic_VIA2 $T=41740 53860 0 0 $X=41270 $Y=53630
X4639 1 DigitalLDOLogic_VIA2 $T=41740 57940 0 0 $X=41270 $Y=57710
X4640 2 DigitalLDOLogic_VIA2 $T=45420 11700 0 0 $X=44950 $Y=11470
X4641 2 DigitalLDOLogic_VIA2 $T=45420 15780 0 0 $X=44950 $Y=15550
X4642 2 DigitalLDOLogic_VIA2 $T=45420 19860 0 0 $X=44950 $Y=19630
X4643 2 DigitalLDOLogic_VIA2 $T=45420 23940 0 0 $X=44950 $Y=23710
X4644 2 DigitalLDOLogic_VIA2 $T=45420 28020 0 0 $X=44950 $Y=27790
X4645 2 DigitalLDOLogic_VIA2 $T=45420 32100 0 0 $X=44950 $Y=31870
X4646 2 DigitalLDOLogic_VIA2 $T=45420 36180 0 0 $X=44950 $Y=35950
X4647 2 DigitalLDOLogic_VIA2 $T=45420 40260 0 0 $X=44950 $Y=40030
X4648 2 DigitalLDOLogic_VIA2 $T=45420 44340 0 0 $X=44950 $Y=44110
X4649 2 DigitalLDOLogic_VIA2 $T=45420 48420 0 0 $X=44950 $Y=48190
X4650 2 DigitalLDOLogic_VIA2 $T=45420 52500 0 0 $X=44950 $Y=52270
X4651 2 DigitalLDOLogic_VIA2 $T=45420 56580 0 0 $X=44950 $Y=56350
X4652 1 DigitalLDOLogic_VIA2 $T=47260 13060 0 0 $X=46790 $Y=12830
X4653 1 DigitalLDOLogic_VIA2 $T=47260 17140 0 0 $X=46790 $Y=16910
X4654 1 DigitalLDOLogic_VIA2 $T=47260 21220 0 0 $X=46790 $Y=20990
X4655 1 DigitalLDOLogic_VIA2 $T=47260 25300 0 0 $X=46790 $Y=25070
X4656 1 DigitalLDOLogic_VIA2 $T=47260 29380 0 0 $X=46790 $Y=29150
X4657 1 DigitalLDOLogic_VIA2 $T=47260 33460 0 0 $X=46790 $Y=33230
X4658 1 DigitalLDOLogic_VIA2 $T=47260 37540 0 0 $X=46790 $Y=37310
X4659 1 DigitalLDOLogic_VIA2 $T=47260 41620 0 0 $X=46790 $Y=41390
X4660 1 DigitalLDOLogic_VIA2 $T=47260 45700 0 0 $X=46790 $Y=45470
X4661 1 DigitalLDOLogic_VIA2 $T=47260 49780 0 0 $X=46790 $Y=49550
X4662 1 DigitalLDOLogic_VIA2 $T=47260 53860 0 0 $X=46790 $Y=53630
X4663 1 DigitalLDOLogic_VIA2 $T=47260 57940 0 0 $X=46790 $Y=57710
X4664 2 DigitalLDOLogic_VIA2 $T=50940 11700 0 0 $X=50470 $Y=11470
X4665 2 DigitalLDOLogic_VIA2 $T=50940 15780 0 0 $X=50470 $Y=15550
X4666 2 DigitalLDOLogic_VIA2 $T=50940 19860 0 0 $X=50470 $Y=19630
X4667 2 DigitalLDOLogic_VIA2 $T=50940 23940 0 0 $X=50470 $Y=23710
X4668 2 DigitalLDOLogic_VIA2 $T=50940 28020 0 0 $X=50470 $Y=27790
X4669 2 DigitalLDOLogic_VIA2 $T=50940 32100 0 0 $X=50470 $Y=31870
X4670 2 DigitalLDOLogic_VIA2 $T=50940 36180 0 0 $X=50470 $Y=35950
X4671 2 DigitalLDOLogic_VIA2 $T=50940 40260 0 0 $X=50470 $Y=40030
X4672 2 DigitalLDOLogic_VIA2 $T=50940 44340 0 0 $X=50470 $Y=44110
X4673 2 DigitalLDOLogic_VIA2 $T=50940 48420 0 0 $X=50470 $Y=48190
X4674 2 DigitalLDOLogic_VIA2 $T=50940 52500 0 0 $X=50470 $Y=52270
X4675 2 DigitalLDOLogic_VIA2 $T=50940 56580 0 0 $X=50470 $Y=56350
X4676 1 DigitalLDOLogic_VIA2 $T=52780 13060 0 0 $X=52310 $Y=12830
X4677 1 DigitalLDOLogic_VIA2 $T=52780 17140 0 0 $X=52310 $Y=16910
X4678 1 DigitalLDOLogic_VIA2 $T=52780 21220 0 0 $X=52310 $Y=20990
X4679 1 DigitalLDOLogic_VIA2 $T=52780 25300 0 0 $X=52310 $Y=25070
X4680 1 DigitalLDOLogic_VIA2 $T=52780 29380 0 0 $X=52310 $Y=29150
X4681 1 DigitalLDOLogic_VIA2 $T=52780 33460 0 0 $X=52310 $Y=33230
X4682 1 DigitalLDOLogic_VIA2 $T=52780 37540 0 0 $X=52310 $Y=37310
X4683 1 DigitalLDOLogic_VIA2 $T=52780 41620 0 0 $X=52310 $Y=41390
X4684 1 DigitalLDOLogic_VIA2 $T=52780 45700 0 0 $X=52310 $Y=45470
X4685 1 DigitalLDOLogic_VIA2 $T=52780 49780 0 0 $X=52310 $Y=49550
X4686 1 DigitalLDOLogic_VIA2 $T=52780 53860 0 0 $X=52310 $Y=53630
X4687 1 DigitalLDOLogic_VIA2 $T=52780 57940 0 0 $X=52310 $Y=57710
X4688 2 DigitalLDOLogic_VIA2 $T=56460 11700 0 0 $X=55990 $Y=11470
X4689 2 DigitalLDOLogic_VIA2 $T=56460 15780 0 0 $X=55990 $Y=15550
X4690 2 DigitalLDOLogic_VIA2 $T=56460 19860 0 0 $X=55990 $Y=19630
X4691 2 DigitalLDOLogic_VIA2 $T=56460 23940 0 0 $X=55990 $Y=23710
X4692 2 DigitalLDOLogic_VIA2 $T=56460 28020 0 0 $X=55990 $Y=27790
X4693 2 DigitalLDOLogic_VIA2 $T=56460 32100 0 0 $X=55990 $Y=31870
X4694 2 DigitalLDOLogic_VIA2 $T=56460 36180 0 0 $X=55990 $Y=35950
X4695 2 DigitalLDOLogic_VIA2 $T=56460 40260 0 0 $X=55990 $Y=40030
X4696 2 DigitalLDOLogic_VIA2 $T=56460 44340 0 0 $X=55990 $Y=44110
X4697 2 DigitalLDOLogic_VIA2 $T=56460 48420 0 0 $X=55990 $Y=48190
X4698 2 DigitalLDOLogic_VIA2 $T=56460 52500 0 0 $X=55990 $Y=52270
X4699 2 DigitalLDOLogic_VIA2 $T=56460 56580 0 0 $X=55990 $Y=56350
X4700 1 DigitalLDOLogic_VIA2 $T=58300 13060 0 0 $X=57830 $Y=12830
X4701 1 DigitalLDOLogic_VIA2 $T=58300 17140 0 0 $X=57830 $Y=16910
X4702 1 DigitalLDOLogic_VIA2 $T=58300 21220 0 0 $X=57830 $Y=20990
X4703 1 DigitalLDOLogic_VIA2 $T=58300 25300 0 0 $X=57830 $Y=25070
X4704 1 DigitalLDOLogic_VIA2 $T=58300 29380 0 0 $X=57830 $Y=29150
X4705 1 DigitalLDOLogic_VIA2 $T=58300 33460 0 0 $X=57830 $Y=33230
X4706 1 DigitalLDOLogic_VIA2 $T=58300 37540 0 0 $X=57830 $Y=37310
X4707 1 DigitalLDOLogic_VIA2 $T=58300 41620 0 0 $X=57830 $Y=41390
X4708 1 DigitalLDOLogic_VIA2 $T=58300 45700 0 0 $X=57830 $Y=45470
X4709 1 DigitalLDOLogic_VIA2 $T=58300 49780 0 0 $X=57830 $Y=49550
X4710 1 DigitalLDOLogic_VIA2 $T=58300 53860 0 0 $X=57830 $Y=53630
X4711 1 DigitalLDOLogic_VIA2 $T=58300 57940 0 0 $X=57830 $Y=57710
X4712 2 DigitalLDOLogic_VIA2 $T=61980 11700 0 0 $X=61510 $Y=11470
X4713 2 DigitalLDOLogic_VIA2 $T=61980 15780 0 0 $X=61510 $Y=15550
X4714 2 DigitalLDOLogic_VIA2 $T=61980 19860 0 0 $X=61510 $Y=19630
X4715 2 DigitalLDOLogic_VIA2 $T=61980 23940 0 0 $X=61510 $Y=23710
X4716 2 DigitalLDOLogic_VIA2 $T=61980 28020 0 0 $X=61510 $Y=27790
X4717 2 DigitalLDOLogic_VIA2 $T=61980 32100 0 0 $X=61510 $Y=31870
X4718 2 DigitalLDOLogic_VIA2 $T=61980 36180 0 0 $X=61510 $Y=35950
X4719 2 DigitalLDOLogic_VIA2 $T=61980 40260 0 0 $X=61510 $Y=40030
X4720 2 DigitalLDOLogic_VIA2 $T=61980 44340 0 0 $X=61510 $Y=44110
X4721 2 DigitalLDOLogic_VIA2 $T=61980 48420 0 0 $X=61510 $Y=48190
X4722 2 DigitalLDOLogic_VIA2 $T=61980 52500 0 0 $X=61510 $Y=52270
X4723 2 DigitalLDOLogic_VIA2 $T=61980 56580 0 0 $X=61510 $Y=56350
X4724 1 DigitalLDOLogic_VIA2 $T=63820 13060 0 0 $X=63350 $Y=12830
X4725 1 DigitalLDOLogic_VIA2 $T=63820 17140 0 0 $X=63350 $Y=16910
X4726 1 DigitalLDOLogic_VIA2 $T=63820 21220 0 0 $X=63350 $Y=20990
X4727 1 DigitalLDOLogic_VIA2 $T=63820 25300 0 0 $X=63350 $Y=25070
X4728 1 DigitalLDOLogic_VIA2 $T=63820 29380 0 0 $X=63350 $Y=29150
X4729 1 DigitalLDOLogic_VIA2 $T=63820 33460 0 0 $X=63350 $Y=33230
X4730 1 DigitalLDOLogic_VIA2 $T=63820 37540 0 0 $X=63350 $Y=37310
X4731 1 DigitalLDOLogic_VIA2 $T=63820 41620 0 0 $X=63350 $Y=41390
X4732 1 DigitalLDOLogic_VIA2 $T=63820 45700 0 0 $X=63350 $Y=45470
X4733 1 DigitalLDOLogic_VIA2 $T=63820 49780 0 0 $X=63350 $Y=49550
X4734 1 DigitalLDOLogic_VIA2 $T=63820 53860 0 0 $X=63350 $Y=53630
X4735 1 DigitalLDOLogic_VIA2 $T=63820 57940 0 0 $X=63350 $Y=57710
X4736 2 DigitalLDOLogic_VIA2 $T=67500 11700 0 0 $X=67030 $Y=11470
X4737 2 DigitalLDOLogic_VIA2 $T=67500 15780 0 0 $X=67030 $Y=15550
X4738 2 DigitalLDOLogic_VIA2 $T=67500 19860 0 0 $X=67030 $Y=19630
X4739 2 DigitalLDOLogic_VIA2 $T=67500 23940 0 0 $X=67030 $Y=23710
X4740 2 DigitalLDOLogic_VIA2 $T=67500 28020 0 0 $X=67030 $Y=27790
X4741 2 DigitalLDOLogic_VIA2 $T=67500 32100 0 0 $X=67030 $Y=31870
X4742 2 DigitalLDOLogic_VIA2 $T=67500 36180 0 0 $X=67030 $Y=35950
X4743 2 DigitalLDOLogic_VIA2 $T=67500 40260 0 0 $X=67030 $Y=40030
X4744 2 DigitalLDOLogic_VIA2 $T=67500 44340 0 0 $X=67030 $Y=44110
X4745 2 DigitalLDOLogic_VIA2 $T=67500 48420 0 0 $X=67030 $Y=48190
X4746 2 DigitalLDOLogic_VIA2 $T=67500 52500 0 0 $X=67030 $Y=52270
X4747 2 DigitalLDOLogic_VIA2 $T=67500 56580 0 0 $X=67030 $Y=56350
X4748 1 DigitalLDOLogic_VIA2 $T=69340 13060 0 0 $X=68870 $Y=12830
X4749 1 DigitalLDOLogic_VIA2 $T=69340 17140 0 0 $X=68870 $Y=16910
X4750 1 DigitalLDOLogic_VIA2 $T=69340 21220 0 0 $X=68870 $Y=20990
X4751 1 DigitalLDOLogic_VIA2 $T=69340 25300 0 0 $X=68870 $Y=25070
X4752 1 DigitalLDOLogic_VIA2 $T=69340 29380 0 0 $X=68870 $Y=29150
X4753 1 DigitalLDOLogic_VIA2 $T=69340 33460 0 0 $X=68870 $Y=33230
X4754 1 DigitalLDOLogic_VIA2 $T=69340 37540 0 0 $X=68870 $Y=37310
X4755 1 DigitalLDOLogic_VIA2 $T=69340 41620 0 0 $X=68870 $Y=41390
X4756 1 DigitalLDOLogic_VIA2 $T=69340 45700 0 0 $X=68870 $Y=45470
X4757 1 DigitalLDOLogic_VIA2 $T=69340 49780 0 0 $X=68870 $Y=49550
X4758 1 DigitalLDOLogic_VIA2 $T=69340 53860 0 0 $X=68870 $Y=53630
X4759 1 DigitalLDOLogic_VIA2 $T=69340 57940 0 0 $X=68870 $Y=57710
X4760 2 DigitalLDOLogic_VIA2 $T=73020 11700 0 0 $X=72550 $Y=11470
X4761 2 DigitalLDOLogic_VIA2 $T=73020 15780 0 0 $X=72550 $Y=15550
X4762 2 DigitalLDOLogic_VIA2 $T=73020 19860 0 0 $X=72550 $Y=19630
X4763 2 DigitalLDOLogic_VIA2 $T=73020 23940 0 0 $X=72550 $Y=23710
X4764 2 DigitalLDOLogic_VIA2 $T=73020 28020 0 0 $X=72550 $Y=27790
X4765 2 DigitalLDOLogic_VIA2 $T=73020 32100 0 0 $X=72550 $Y=31870
X4766 2 DigitalLDOLogic_VIA2 $T=73020 36180 0 0 $X=72550 $Y=35950
X4767 2 DigitalLDOLogic_VIA2 $T=73020 40260 0 0 $X=72550 $Y=40030
X4768 2 DigitalLDOLogic_VIA2 $T=73020 44340 0 0 $X=72550 $Y=44110
X4769 2 DigitalLDOLogic_VIA2 $T=73020 48420 0 0 $X=72550 $Y=48190
X4770 2 DigitalLDOLogic_VIA2 $T=73020 52500 0 0 $X=72550 $Y=52270
X4771 2 DigitalLDOLogic_VIA2 $T=73020 56580 0 0 $X=72550 $Y=56350
X4772 1 DigitalLDOLogic_VIA2 $T=74860 13060 0 0 $X=74390 $Y=12830
X4773 1 DigitalLDOLogic_VIA2 $T=74860 17140 0 0 $X=74390 $Y=16910
X4774 1 DigitalLDOLogic_VIA2 $T=74860 21220 0 0 $X=74390 $Y=20990
X4775 1 DigitalLDOLogic_VIA2 $T=74860 25300 0 0 $X=74390 $Y=25070
X4776 1 DigitalLDOLogic_VIA2 $T=74860 29380 0 0 $X=74390 $Y=29150
X4777 1 DigitalLDOLogic_VIA2 $T=74860 33460 0 0 $X=74390 $Y=33230
X4778 1 DigitalLDOLogic_VIA2 $T=74860 37540 0 0 $X=74390 $Y=37310
X4779 1 DigitalLDOLogic_VIA2 $T=74860 41620 0 0 $X=74390 $Y=41390
X4780 1 DigitalLDOLogic_VIA2 $T=74860 45700 0 0 $X=74390 $Y=45470
X4781 1 DigitalLDOLogic_VIA2 $T=74860 49780 0 0 $X=74390 $Y=49550
X4782 1 DigitalLDOLogic_VIA2 $T=74860 53860 0 0 $X=74390 $Y=53630
X4783 1 DigitalLDOLogic_VIA2 $T=74860 57940 0 0 $X=74390 $Y=57710
X4784 2 DigitalLDOLogic_VIA2 $T=78540 11700 0 0 $X=78070 $Y=11470
X4785 2 DigitalLDOLogic_VIA2 $T=78540 15780 0 0 $X=78070 $Y=15550
X4786 2 DigitalLDOLogic_VIA2 $T=78540 19860 0 0 $X=78070 $Y=19630
X4787 2 DigitalLDOLogic_VIA2 $T=78540 23940 0 0 $X=78070 $Y=23710
X4788 2 DigitalLDOLogic_VIA2 $T=78540 28020 0 0 $X=78070 $Y=27790
X4789 2 DigitalLDOLogic_VIA2 $T=78540 32100 0 0 $X=78070 $Y=31870
X4790 2 DigitalLDOLogic_VIA2 $T=78540 36180 0 0 $X=78070 $Y=35950
X4791 2 DigitalLDOLogic_VIA2 $T=78540 40260 0 0 $X=78070 $Y=40030
X4792 2 DigitalLDOLogic_VIA2 $T=78540 44340 0 0 $X=78070 $Y=44110
X4793 2 DigitalLDOLogic_VIA2 $T=78540 48420 0 0 $X=78070 $Y=48190
X4794 2 DigitalLDOLogic_VIA2 $T=78540 52500 0 0 $X=78070 $Y=52270
X4795 2 DigitalLDOLogic_VIA2 $T=78540 56580 0 0 $X=78070 $Y=56350
X4796 1 DigitalLDOLogic_VIA2 $T=80380 13060 0 0 $X=79910 $Y=12830
X4797 1 DigitalLDOLogic_VIA2 $T=80380 17140 0 0 $X=79910 $Y=16910
X4798 1 DigitalLDOLogic_VIA2 $T=80380 21220 0 0 $X=79910 $Y=20990
X4799 1 DigitalLDOLogic_VIA2 $T=80380 25300 0 0 $X=79910 $Y=25070
X4800 1 DigitalLDOLogic_VIA2 $T=80380 29380 0 0 $X=79910 $Y=29150
X4801 1 DigitalLDOLogic_VIA2 $T=80380 33460 0 0 $X=79910 $Y=33230
X4802 1 DigitalLDOLogic_VIA2 $T=80380 37540 0 0 $X=79910 $Y=37310
X4803 1 DigitalLDOLogic_VIA2 $T=80380 41620 0 0 $X=79910 $Y=41390
X4804 1 DigitalLDOLogic_VIA2 $T=80380 45700 0 0 $X=79910 $Y=45470
X4805 1 DigitalLDOLogic_VIA2 $T=80380 49780 0 0 $X=79910 $Y=49550
X4806 1 DigitalLDOLogic_VIA2 $T=80380 53860 0 0 $X=79910 $Y=53630
X4807 1 DigitalLDOLogic_VIA2 $T=80380 57940 0 0 $X=79910 $Y=57710
X4808 2 DigitalLDOLogic_VIA2 $T=84060 11700 0 0 $X=83590 $Y=11470
X4809 2 DigitalLDOLogic_VIA2 $T=84060 15780 0 0 $X=83590 $Y=15550
X4810 2 DigitalLDOLogic_VIA2 $T=84060 19860 0 0 $X=83590 $Y=19630
X4811 2 DigitalLDOLogic_VIA2 $T=84060 23940 0 0 $X=83590 $Y=23710
X4812 2 DigitalLDOLogic_VIA2 $T=84060 28020 0 0 $X=83590 $Y=27790
X4813 2 DigitalLDOLogic_VIA2 $T=84060 32100 0 0 $X=83590 $Y=31870
X4814 2 DigitalLDOLogic_VIA2 $T=84060 36180 0 0 $X=83590 $Y=35950
X4815 2 DigitalLDOLogic_VIA2 $T=84060 40260 0 0 $X=83590 $Y=40030
X4816 2 DigitalLDOLogic_VIA2 $T=84060 44340 0 0 $X=83590 $Y=44110
X4817 2 DigitalLDOLogic_VIA2 $T=84060 48420 0 0 $X=83590 $Y=48190
X4818 2 DigitalLDOLogic_VIA2 $T=84060 52500 0 0 $X=83590 $Y=52270
X4819 2 DigitalLDOLogic_VIA2 $T=84060 56580 0 0 $X=83590 $Y=56350
X4820 1 DigitalLDOLogic_VIA2 $T=85900 13060 0 0 $X=85430 $Y=12830
X4821 1 DigitalLDOLogic_VIA2 $T=85900 17140 0 0 $X=85430 $Y=16910
X4822 1 DigitalLDOLogic_VIA2 $T=85900 21220 0 0 $X=85430 $Y=20990
X4823 1 DigitalLDOLogic_VIA2 $T=85900 25300 0 0 $X=85430 $Y=25070
X4824 1 DigitalLDOLogic_VIA2 $T=85900 29380 0 0 $X=85430 $Y=29150
X4825 1 DigitalLDOLogic_VIA2 $T=85900 33460 0 0 $X=85430 $Y=33230
X4826 1 DigitalLDOLogic_VIA2 $T=85900 37540 0 0 $X=85430 $Y=37310
X4827 1 DigitalLDOLogic_VIA2 $T=85900 41620 0 0 $X=85430 $Y=41390
X4828 1 DigitalLDOLogic_VIA2 $T=85900 45700 0 0 $X=85430 $Y=45470
X4829 1 DigitalLDOLogic_VIA2 $T=85900 49780 0 0 $X=85430 $Y=49550
X4830 1 DigitalLDOLogic_VIA2 $T=85900 53860 0 0 $X=85430 $Y=53630
X4831 1 DigitalLDOLogic_VIA2 $T=85900 57940 0 0 $X=85430 $Y=57710
X4832 2 DigitalLDOLogic_VIA2 $T=89580 11700 0 0 $X=89110 $Y=11470
X4833 2 DigitalLDOLogic_VIA2 $T=89580 15780 0 0 $X=89110 $Y=15550
X4834 2 DigitalLDOLogic_VIA2 $T=89580 19860 0 0 $X=89110 $Y=19630
X4835 2 DigitalLDOLogic_VIA2 $T=89580 23940 0 0 $X=89110 $Y=23710
X4836 2 DigitalLDOLogic_VIA2 $T=89580 28020 0 0 $X=89110 $Y=27790
X4837 2 DigitalLDOLogic_VIA2 $T=89580 32100 0 0 $X=89110 $Y=31870
X4838 2 DigitalLDOLogic_VIA2 $T=89580 36180 0 0 $X=89110 $Y=35950
X4839 2 DigitalLDOLogic_VIA2 $T=89580 40260 0 0 $X=89110 $Y=40030
X4840 2 DigitalLDOLogic_VIA2 $T=89580 44340 0 0 $X=89110 $Y=44110
X4841 2 DigitalLDOLogic_VIA2 $T=89580 48420 0 0 $X=89110 $Y=48190
X4842 2 DigitalLDOLogic_VIA2 $T=89580 52500 0 0 $X=89110 $Y=52270
X4843 2 DigitalLDOLogic_VIA2 $T=89580 56580 0 0 $X=89110 $Y=56350
X4844 1 DigitalLDOLogic_VIA2 $T=91420 13060 0 0 $X=90950 $Y=12830
X4845 1 DigitalLDOLogic_VIA2 $T=91420 17140 0 0 $X=90950 $Y=16910
X4846 1 DigitalLDOLogic_VIA2 $T=91420 21220 0 0 $X=90950 $Y=20990
X4847 1 DigitalLDOLogic_VIA2 $T=91420 25300 0 0 $X=90950 $Y=25070
X4848 1 DigitalLDOLogic_VIA2 $T=91420 29380 0 0 $X=90950 $Y=29150
X4849 1 DigitalLDOLogic_VIA2 $T=91420 33460 0 0 $X=90950 $Y=33230
X4850 1 DigitalLDOLogic_VIA2 $T=91420 37540 0 0 $X=90950 $Y=37310
X4851 1 DigitalLDOLogic_VIA2 $T=91420 41620 0 0 $X=90950 $Y=41390
X4852 1 DigitalLDOLogic_VIA2 $T=91420 45700 0 0 $X=90950 $Y=45470
X4853 1 DigitalLDOLogic_VIA2 $T=91420 49780 0 0 $X=90950 $Y=49550
X4854 1 DigitalLDOLogic_VIA2 $T=91420 53860 0 0 $X=90950 $Y=53630
X4855 1 DigitalLDOLogic_VIA2 $T=91420 57940 0 0 $X=90950 $Y=57710
X4856 2 DigitalLDOLogic_VIA2 $T=95100 11700 0 0 $X=94630 $Y=11470
X4857 2 DigitalLDOLogic_VIA2 $T=95100 15780 0 0 $X=94630 $Y=15550
X4858 2 DigitalLDOLogic_VIA2 $T=95100 19860 0 0 $X=94630 $Y=19630
X4859 2 DigitalLDOLogic_VIA2 $T=95100 23940 0 0 $X=94630 $Y=23710
X4860 2 DigitalLDOLogic_VIA2 $T=95100 28020 0 0 $X=94630 $Y=27790
X4861 2 DigitalLDOLogic_VIA2 $T=95100 32100 0 0 $X=94630 $Y=31870
X4862 2 DigitalLDOLogic_VIA2 $T=95100 36180 0 0 $X=94630 $Y=35950
X4863 2 DigitalLDOLogic_VIA2 $T=95100 40260 0 0 $X=94630 $Y=40030
X4864 2 DigitalLDOLogic_VIA2 $T=95100 44340 0 0 $X=94630 $Y=44110
X4865 2 DigitalLDOLogic_VIA2 $T=95100 48420 0 0 $X=94630 $Y=48190
X4866 2 DigitalLDOLogic_VIA2 $T=95100 52500 0 0 $X=94630 $Y=52270
X4867 2 DigitalLDOLogic_VIA2 $T=95100 56580 0 0 $X=94630 $Y=56350
X4868 1 DigitalLDOLogic_VIA2 $T=96940 13060 0 0 $X=96470 $Y=12830
X4869 1 DigitalLDOLogic_VIA2 $T=96940 17140 0 0 $X=96470 $Y=16910
X4870 1 DigitalLDOLogic_VIA2 $T=96940 21220 0 0 $X=96470 $Y=20990
X4871 1 DigitalLDOLogic_VIA2 $T=96940 25300 0 0 $X=96470 $Y=25070
X4872 1 DigitalLDOLogic_VIA2 $T=96940 29380 0 0 $X=96470 $Y=29150
X4873 1 DigitalLDOLogic_VIA2 $T=96940 33460 0 0 $X=96470 $Y=33230
X4874 1 DigitalLDOLogic_VIA2 $T=96940 37540 0 0 $X=96470 $Y=37310
X4875 1 DigitalLDOLogic_VIA2 $T=96940 41620 0 0 $X=96470 $Y=41390
X4876 1 DigitalLDOLogic_VIA2 $T=96940 45700 0 0 $X=96470 $Y=45470
X4877 1 DigitalLDOLogic_VIA2 $T=96940 49780 0 0 $X=96470 $Y=49550
X4878 1 DigitalLDOLogic_VIA2 $T=96940 53860 0 0 $X=96470 $Y=53630
X4879 1 DigitalLDOLogic_VIA2 $T=96940 57940 0 0 $X=96470 $Y=57710
X4880 2 DigitalLDOLogic_VIA2 $T=100620 11700 0 0 $X=100150 $Y=11470
X4881 2 DigitalLDOLogic_VIA2 $T=100620 15780 0 0 $X=100150 $Y=15550
X4882 2 DigitalLDOLogic_VIA2 $T=100620 19860 0 0 $X=100150 $Y=19630
X4883 2 DigitalLDOLogic_VIA2 $T=100620 23940 0 0 $X=100150 $Y=23710
X4884 2 DigitalLDOLogic_VIA2 $T=100620 28020 0 0 $X=100150 $Y=27790
X4885 2 DigitalLDOLogic_VIA2 $T=100620 32100 0 0 $X=100150 $Y=31870
X4886 2 DigitalLDOLogic_VIA2 $T=100620 36180 0 0 $X=100150 $Y=35950
X4887 2 DigitalLDOLogic_VIA2 $T=100620 40260 0 0 $X=100150 $Y=40030
X4888 2 DigitalLDOLogic_VIA2 $T=100620 44340 0 0 $X=100150 $Y=44110
X4889 2 DigitalLDOLogic_VIA2 $T=100620 48420 0 0 $X=100150 $Y=48190
X4890 2 DigitalLDOLogic_VIA2 $T=100620 52500 0 0 $X=100150 $Y=52270
X4891 2 DigitalLDOLogic_VIA2 $T=100620 56580 0 0 $X=100150 $Y=56350
X4892 1 DigitalLDOLogic_VIA2 $T=102460 13060 0 0 $X=101990 $Y=12830
X4893 1 DigitalLDOLogic_VIA2 $T=102460 17140 0 0 $X=101990 $Y=16910
X4894 1 DigitalLDOLogic_VIA2 $T=102460 21220 0 0 $X=101990 $Y=20990
X4895 1 DigitalLDOLogic_VIA2 $T=102460 25300 0 0 $X=101990 $Y=25070
X4896 1 DigitalLDOLogic_VIA2 $T=102460 29380 0 0 $X=101990 $Y=29150
X4897 1 DigitalLDOLogic_VIA2 $T=102460 33460 0 0 $X=101990 $Y=33230
X4898 1 DigitalLDOLogic_VIA2 $T=102460 37540 0 0 $X=101990 $Y=37310
X4899 1 DigitalLDOLogic_VIA2 $T=102460 41620 0 0 $X=101990 $Y=41390
X4900 1 DigitalLDOLogic_VIA2 $T=102460 45700 0 0 $X=101990 $Y=45470
X4901 1 DigitalLDOLogic_VIA2 $T=102460 49780 0 0 $X=101990 $Y=49550
X4902 1 DigitalLDOLogic_VIA2 $T=102460 53860 0 0 $X=101990 $Y=53630
X4903 1 DigitalLDOLogic_VIA2 $T=102460 57940 0 0 $X=101990 $Y=57710
X4904 2 DigitalLDOLogic_VIA2 $T=106140 11700 0 0 $X=105670 $Y=11470
X4905 2 DigitalLDOLogic_VIA2 $T=106140 15780 0 0 $X=105670 $Y=15550
X4906 2 DigitalLDOLogic_VIA2 $T=106140 19860 0 0 $X=105670 $Y=19630
X4907 2 DigitalLDOLogic_VIA2 $T=106140 23940 0 0 $X=105670 $Y=23710
X4908 2 DigitalLDOLogic_VIA2 $T=106140 28020 0 0 $X=105670 $Y=27790
X4909 2 DigitalLDOLogic_VIA2 $T=106140 32100 0 0 $X=105670 $Y=31870
X4910 2 DigitalLDOLogic_VIA2 $T=106140 36180 0 0 $X=105670 $Y=35950
X4911 2 DigitalLDOLogic_VIA2 $T=106140 40260 0 0 $X=105670 $Y=40030
X4912 2 DigitalLDOLogic_VIA2 $T=106140 44340 0 0 $X=105670 $Y=44110
X4913 2 DigitalLDOLogic_VIA2 $T=106140 48420 0 0 $X=105670 $Y=48190
X4914 2 DigitalLDOLogic_VIA2 $T=106140 52500 0 0 $X=105670 $Y=52270
X4915 2 DigitalLDOLogic_VIA2 $T=106140 56580 0 0 $X=105670 $Y=56350
X4916 1 DigitalLDOLogic_VIA2 $T=107980 13060 0 0 $X=107510 $Y=12830
X4917 1 DigitalLDOLogic_VIA2 $T=107980 17140 0 0 $X=107510 $Y=16910
X4918 1 DigitalLDOLogic_VIA2 $T=107980 21220 0 0 $X=107510 $Y=20990
X4919 1 DigitalLDOLogic_VIA2 $T=107980 25300 0 0 $X=107510 $Y=25070
X4920 1 DigitalLDOLogic_VIA2 $T=107980 29380 0 0 $X=107510 $Y=29150
X4921 1 DigitalLDOLogic_VIA2 $T=107980 33460 0 0 $X=107510 $Y=33230
X4922 1 DigitalLDOLogic_VIA2 $T=107980 37540 0 0 $X=107510 $Y=37310
X4923 1 DigitalLDOLogic_VIA2 $T=107980 41620 0 0 $X=107510 $Y=41390
X4924 1 DigitalLDOLogic_VIA2 $T=107980 45700 0 0 $X=107510 $Y=45470
X4925 1 DigitalLDOLogic_VIA2 $T=107980 49780 0 0 $X=107510 $Y=49550
X4926 1 DigitalLDOLogic_VIA2 $T=107980 53860 0 0 $X=107510 $Y=53630
X4927 1 DigitalLDOLogic_VIA2 $T=107980 57940 0 0 $X=107510 $Y=57710
X4928 2 DigitalLDOLogic_VIA2 $T=111660 11700 0 0 $X=111190 $Y=11470
X4929 2 DigitalLDOLogic_VIA2 $T=111660 15780 0 0 $X=111190 $Y=15550
X4930 2 DigitalLDOLogic_VIA2 $T=111660 19860 0 0 $X=111190 $Y=19630
X4931 2 DigitalLDOLogic_VIA2 $T=111660 23940 0 0 $X=111190 $Y=23710
X4932 2 DigitalLDOLogic_VIA2 $T=111660 28020 0 0 $X=111190 $Y=27790
X4933 2 DigitalLDOLogic_VIA2 $T=111660 32100 0 0 $X=111190 $Y=31870
X4934 2 DigitalLDOLogic_VIA2 $T=111660 36180 0 0 $X=111190 $Y=35950
X4935 2 DigitalLDOLogic_VIA2 $T=111660 40260 0 0 $X=111190 $Y=40030
X4936 2 DigitalLDOLogic_VIA2 $T=111660 44340 0 0 $X=111190 $Y=44110
X4937 2 DigitalLDOLogic_VIA2 $T=111660 48420 0 0 $X=111190 $Y=48190
X4938 2 DigitalLDOLogic_VIA2 $T=111660 52500 0 0 $X=111190 $Y=52270
X4939 2 DigitalLDOLogic_VIA2 $T=111660 56580 0 0 $X=111190 $Y=56350
X4940 1 DigitalLDOLogic_VIA2 $T=113500 13060 0 0 $X=113030 $Y=12830
X4941 1 DigitalLDOLogic_VIA2 $T=113500 17140 0 0 $X=113030 $Y=16910
X4942 1 DigitalLDOLogic_VIA2 $T=113500 21220 0 0 $X=113030 $Y=20990
X4943 1 DigitalLDOLogic_VIA2 $T=113500 25300 0 0 $X=113030 $Y=25070
X4944 1 DigitalLDOLogic_VIA2 $T=113500 29380 0 0 $X=113030 $Y=29150
X4945 1 DigitalLDOLogic_VIA2 $T=113500 33460 0 0 $X=113030 $Y=33230
X4946 1 DigitalLDOLogic_VIA2 $T=113500 37540 0 0 $X=113030 $Y=37310
X4947 1 DigitalLDOLogic_VIA2 $T=113500 41620 0 0 $X=113030 $Y=41390
X4948 1 DigitalLDOLogic_VIA2 $T=113500 45700 0 0 $X=113030 $Y=45470
X4949 1 DigitalLDOLogic_VIA2 $T=113500 49780 0 0 $X=113030 $Y=49550
X4950 1 DigitalLDOLogic_VIA2 $T=113500 53860 0 0 $X=113030 $Y=53630
X4951 1 DigitalLDOLogic_VIA2 $T=113500 57940 0 0 $X=113030 $Y=57710
X4952 2 DigitalLDOLogic_VIA2 $T=117180 11700 0 0 $X=116710 $Y=11470
X4953 2 DigitalLDOLogic_VIA2 $T=117180 15780 0 0 $X=116710 $Y=15550
X4954 2 DigitalLDOLogic_VIA2 $T=117180 19860 0 0 $X=116710 $Y=19630
X4955 2 DigitalLDOLogic_VIA2 $T=117180 23940 0 0 $X=116710 $Y=23710
X4956 2 DigitalLDOLogic_VIA2 $T=117180 28020 0 0 $X=116710 $Y=27790
X4957 2 DigitalLDOLogic_VIA2 $T=117180 32100 0 0 $X=116710 $Y=31870
X4958 2 DigitalLDOLogic_VIA2 $T=117180 36180 0 0 $X=116710 $Y=35950
X4959 2 DigitalLDOLogic_VIA2 $T=117180 40260 0 0 $X=116710 $Y=40030
X4960 2 DigitalLDOLogic_VIA2 $T=117180 44340 0 0 $X=116710 $Y=44110
X4961 2 DigitalLDOLogic_VIA2 $T=117180 48420 0 0 $X=116710 $Y=48190
X4962 2 DigitalLDOLogic_VIA2 $T=117180 52500 0 0 $X=116710 $Y=52270
X4963 2 DigitalLDOLogic_VIA2 $T=117180 56580 0 0 $X=116710 $Y=56350
X4964 1 DigitalLDOLogic_VIA2 $T=119020 13060 0 0 $X=118550 $Y=12830
X4965 1 DigitalLDOLogic_VIA2 $T=119020 17140 0 0 $X=118550 $Y=16910
X4966 1 DigitalLDOLogic_VIA2 $T=119020 21220 0 0 $X=118550 $Y=20990
X4967 1 DigitalLDOLogic_VIA2 $T=119020 25300 0 0 $X=118550 $Y=25070
X4968 1 DigitalLDOLogic_VIA2 $T=119020 29380 0 0 $X=118550 $Y=29150
X4969 1 DigitalLDOLogic_VIA2 $T=119020 33460 0 0 $X=118550 $Y=33230
X4970 1 DigitalLDOLogic_VIA2 $T=119020 37540 0 0 $X=118550 $Y=37310
X4971 1 DigitalLDOLogic_VIA2 $T=119020 41620 0 0 $X=118550 $Y=41390
X4972 1 DigitalLDOLogic_VIA2 $T=119020 45700 0 0 $X=118550 $Y=45470
X4973 1 DigitalLDOLogic_VIA2 $T=119020 49780 0 0 $X=118550 $Y=49550
X4974 1 DigitalLDOLogic_VIA2 $T=119020 53860 0 0 $X=118550 $Y=53630
X4975 1 DigitalLDOLogic_VIA2 $T=119020 57940 0 0 $X=118550 $Y=57710
X4976 2 DigitalLDOLogic_VIA2 $T=122700 11700 0 0 $X=122230 $Y=11470
X4977 2 DigitalLDOLogic_VIA2 $T=122700 15780 0 0 $X=122230 $Y=15550
X4978 2 DigitalLDOLogic_VIA2 $T=122700 19860 0 0 $X=122230 $Y=19630
X4979 2 DigitalLDOLogic_VIA2 $T=122700 23940 0 0 $X=122230 $Y=23710
X4980 2 DigitalLDOLogic_VIA2 $T=122700 28020 0 0 $X=122230 $Y=27790
X4981 2 DigitalLDOLogic_VIA2 $T=122700 32100 0 0 $X=122230 $Y=31870
X4982 2 DigitalLDOLogic_VIA2 $T=122700 36180 0 0 $X=122230 $Y=35950
X4983 2 DigitalLDOLogic_VIA2 $T=122700 40260 0 0 $X=122230 $Y=40030
X4984 2 DigitalLDOLogic_VIA2 $T=122700 44340 0 0 $X=122230 $Y=44110
X4985 2 DigitalLDOLogic_VIA2 $T=122700 48420 0 0 $X=122230 $Y=48190
X4986 2 DigitalLDOLogic_VIA2 $T=122700 52500 0 0 $X=122230 $Y=52270
X4987 2 DigitalLDOLogic_VIA2 $T=122700 56580 0 0 $X=122230 $Y=56350
X4988 1 DigitalLDOLogic_VIA2 $T=124540 13060 0 0 $X=124070 $Y=12830
X4989 1 DigitalLDOLogic_VIA2 $T=124540 17140 0 0 $X=124070 $Y=16910
X4990 1 DigitalLDOLogic_VIA2 $T=124540 21220 0 0 $X=124070 $Y=20990
X4991 1 DigitalLDOLogic_VIA2 $T=124540 25300 0 0 $X=124070 $Y=25070
X4992 1 DigitalLDOLogic_VIA2 $T=124540 29380 0 0 $X=124070 $Y=29150
X4993 1 DigitalLDOLogic_VIA2 $T=124540 33460 0 0 $X=124070 $Y=33230
X4994 1 DigitalLDOLogic_VIA2 $T=124540 37540 0 0 $X=124070 $Y=37310
X4995 1 DigitalLDOLogic_VIA2 $T=124540 41620 0 0 $X=124070 $Y=41390
X4996 1 DigitalLDOLogic_VIA2 $T=124540 45700 0 0 $X=124070 $Y=45470
X4997 1 DigitalLDOLogic_VIA2 $T=124540 49780 0 0 $X=124070 $Y=49550
X4998 1 DigitalLDOLogic_VIA2 $T=124540 53860 0 0 $X=124070 $Y=53630
X4999 1 DigitalLDOLogic_VIA2 $T=124540 57940 0 0 $X=124070 $Y=57710
X5000 2 DigitalLDOLogic_VIA2 $T=128220 11700 0 0 $X=127750 $Y=11470
X5001 2 DigitalLDOLogic_VIA2 $T=128220 15780 0 0 $X=127750 $Y=15550
X5002 2 DigitalLDOLogic_VIA2 $T=128220 19860 0 0 $X=127750 $Y=19630
X5003 2 DigitalLDOLogic_VIA2 $T=128220 23940 0 0 $X=127750 $Y=23710
X5004 2 DigitalLDOLogic_VIA2 $T=128220 28020 0 0 $X=127750 $Y=27790
X5005 2 DigitalLDOLogic_VIA2 $T=128220 32100 0 0 $X=127750 $Y=31870
X5006 2 DigitalLDOLogic_VIA2 $T=128220 36180 0 0 $X=127750 $Y=35950
X5007 2 DigitalLDOLogic_VIA2 $T=128220 40260 0 0 $X=127750 $Y=40030
X5008 2 DigitalLDOLogic_VIA2 $T=128220 44340 0 0 $X=127750 $Y=44110
X5009 2 DigitalLDOLogic_VIA2 $T=128220 48420 0 0 $X=127750 $Y=48190
X5010 2 DigitalLDOLogic_VIA2 $T=128220 52500 0 0 $X=127750 $Y=52270
X5011 2 DigitalLDOLogic_VIA2 $T=128220 56580 0 0 $X=127750 $Y=56350
X5012 1 DigitalLDOLogic_VIA2 $T=130060 13060 0 0 $X=129590 $Y=12830
X5013 1 DigitalLDOLogic_VIA2 $T=130060 17140 0 0 $X=129590 $Y=16910
X5014 1 DigitalLDOLogic_VIA2 $T=130060 21220 0 0 $X=129590 $Y=20990
X5015 1 DigitalLDOLogic_VIA2 $T=130060 25300 0 0 $X=129590 $Y=25070
X5016 1 DigitalLDOLogic_VIA2 $T=130060 29380 0 0 $X=129590 $Y=29150
X5017 1 DigitalLDOLogic_VIA2 $T=130060 33460 0 0 $X=129590 $Y=33230
X5018 1 DigitalLDOLogic_VIA2 $T=130060 37540 0 0 $X=129590 $Y=37310
X5019 1 DigitalLDOLogic_VIA2 $T=130060 41620 0 0 $X=129590 $Y=41390
X5020 1 DigitalLDOLogic_VIA2 $T=130060 45700 0 0 $X=129590 $Y=45470
X5021 1 DigitalLDOLogic_VIA2 $T=130060 49780 0 0 $X=129590 $Y=49550
X5022 1 DigitalLDOLogic_VIA2 $T=130060 53860 0 0 $X=129590 $Y=53630
X5023 1 DigitalLDOLogic_VIA2 $T=130060 57940 0 0 $X=129590 $Y=57710
X5024 2 DigitalLDOLogic_VIA2 $T=133740 11700 0 0 $X=133270 $Y=11470
X5025 2 DigitalLDOLogic_VIA2 $T=133740 15780 0 0 $X=133270 $Y=15550
X5026 2 DigitalLDOLogic_VIA2 $T=133740 19860 0 0 $X=133270 $Y=19630
X5027 2 DigitalLDOLogic_VIA2 $T=133740 23940 0 0 $X=133270 $Y=23710
X5028 2 DigitalLDOLogic_VIA2 $T=133740 28020 0 0 $X=133270 $Y=27790
X5029 2 DigitalLDOLogic_VIA2 $T=133740 32100 0 0 $X=133270 $Y=31870
X5030 2 DigitalLDOLogic_VIA2 $T=133740 36180 0 0 $X=133270 $Y=35950
X5031 2 DigitalLDOLogic_VIA2 $T=133740 40260 0 0 $X=133270 $Y=40030
X5032 2 DigitalLDOLogic_VIA2 $T=133740 44340 0 0 $X=133270 $Y=44110
X5033 2 DigitalLDOLogic_VIA2 $T=133740 48420 0 0 $X=133270 $Y=48190
X5034 2 DigitalLDOLogic_VIA2 $T=133740 52500 0 0 $X=133270 $Y=52270
X5035 2 DigitalLDOLogic_VIA2 $T=133740 56580 0 0 $X=133270 $Y=56350
X5036 1 DigitalLDOLogic_VIA2 $T=135580 13060 0 0 $X=135110 $Y=12830
X5037 1 DigitalLDOLogic_VIA2 $T=135580 17140 0 0 $X=135110 $Y=16910
X5038 1 DigitalLDOLogic_VIA2 $T=135580 21220 0 0 $X=135110 $Y=20990
X5039 1 DigitalLDOLogic_VIA2 $T=135580 25300 0 0 $X=135110 $Y=25070
X5040 1 DigitalLDOLogic_VIA2 $T=135580 29380 0 0 $X=135110 $Y=29150
X5041 1 DigitalLDOLogic_VIA2 $T=135580 33460 0 0 $X=135110 $Y=33230
X5042 1 DigitalLDOLogic_VIA2 $T=135580 37540 0 0 $X=135110 $Y=37310
X5043 1 DigitalLDOLogic_VIA2 $T=135580 41620 0 0 $X=135110 $Y=41390
X5044 1 DigitalLDOLogic_VIA2 $T=135580 45700 0 0 $X=135110 $Y=45470
X5045 1 DigitalLDOLogic_VIA2 $T=135580 49780 0 0 $X=135110 $Y=49550
X5046 1 DigitalLDOLogic_VIA2 $T=135580 53860 0 0 $X=135110 $Y=53630
X5047 1 DigitalLDOLogic_VIA2 $T=135580 57940 0 0 $X=135110 $Y=57710
X5048 2 DigitalLDOLogic_VIA2 $T=139260 11700 0 0 $X=138790 $Y=11470
X5049 2 DigitalLDOLogic_VIA2 $T=139260 15780 0 0 $X=138790 $Y=15550
X5050 2 DigitalLDOLogic_VIA2 $T=139260 19860 0 0 $X=138790 $Y=19630
X5051 2 DigitalLDOLogic_VIA2 $T=139260 23940 0 0 $X=138790 $Y=23710
X5052 2 DigitalLDOLogic_VIA2 $T=139260 28020 0 0 $X=138790 $Y=27790
X5053 2 DigitalLDOLogic_VIA2 $T=139260 32100 0 0 $X=138790 $Y=31870
X5054 2 DigitalLDOLogic_VIA2 $T=139260 36180 0 0 $X=138790 $Y=35950
X5055 2 DigitalLDOLogic_VIA2 $T=139260 40260 0 0 $X=138790 $Y=40030
X5056 2 DigitalLDOLogic_VIA2 $T=139260 44340 0 0 $X=138790 $Y=44110
X5057 2 DigitalLDOLogic_VIA2 $T=139260 48420 0 0 $X=138790 $Y=48190
X5058 2 DigitalLDOLogic_VIA2 $T=139260 52500 0 0 $X=138790 $Y=52270
X5059 2 DigitalLDOLogic_VIA2 $T=139260 56580 0 0 $X=138790 $Y=56350
X5060 1 DigitalLDOLogic_VIA2 $T=141100 13060 0 0 $X=140630 $Y=12830
X5061 1 DigitalLDOLogic_VIA2 $T=141100 17140 0 0 $X=140630 $Y=16910
X5062 1 DigitalLDOLogic_VIA2 $T=141100 21220 0 0 $X=140630 $Y=20990
X5063 1 DigitalLDOLogic_VIA2 $T=141100 25300 0 0 $X=140630 $Y=25070
X5064 1 DigitalLDOLogic_VIA2 $T=141100 29380 0 0 $X=140630 $Y=29150
X5065 1 DigitalLDOLogic_VIA2 $T=141100 33460 0 0 $X=140630 $Y=33230
X5066 1 DigitalLDOLogic_VIA2 $T=141100 37540 0 0 $X=140630 $Y=37310
X5067 1 DigitalLDOLogic_VIA2 $T=141100 41620 0 0 $X=140630 $Y=41390
X5068 1 DigitalLDOLogic_VIA2 $T=141100 45700 0 0 $X=140630 $Y=45470
X5069 1 DigitalLDOLogic_VIA2 $T=141100 49780 0 0 $X=140630 $Y=49550
X5070 1 DigitalLDOLogic_VIA2 $T=141100 53860 0 0 $X=140630 $Y=53630
X5071 1 DigitalLDOLogic_VIA2 $T=141100 57940 0 0 $X=140630 $Y=57710
X5072 2 DigitalLDOLogic_VIA2 $T=144780 11700 0 0 $X=144310 $Y=11470
X5073 2 DigitalLDOLogic_VIA2 $T=144780 15780 0 0 $X=144310 $Y=15550
X5074 2 DigitalLDOLogic_VIA2 $T=144780 19860 0 0 $X=144310 $Y=19630
X5075 2 DigitalLDOLogic_VIA2 $T=144780 23940 0 0 $X=144310 $Y=23710
X5076 2 DigitalLDOLogic_VIA2 $T=144780 28020 0 0 $X=144310 $Y=27790
X5077 2 DigitalLDOLogic_VIA2 $T=144780 32100 0 0 $X=144310 $Y=31870
X5078 2 DigitalLDOLogic_VIA2 $T=144780 36180 0 0 $X=144310 $Y=35950
X5079 2 DigitalLDOLogic_VIA2 $T=144780 40260 0 0 $X=144310 $Y=40030
X5080 2 DigitalLDOLogic_VIA2 $T=144780 44340 0 0 $X=144310 $Y=44110
X5081 2 DigitalLDOLogic_VIA2 $T=144780 48420 0 0 $X=144310 $Y=48190
X5082 2 DigitalLDOLogic_VIA2 $T=144780 52500 0 0 $X=144310 $Y=52270
X5083 2 DigitalLDOLogic_VIA2 $T=144780 56580 0 0 $X=144310 $Y=56350
X5084 1 DigitalLDOLogic_VIA2 $T=146620 13060 0 0 $X=146150 $Y=12830
X5085 1 DigitalLDOLogic_VIA2 $T=146620 17140 0 0 $X=146150 $Y=16910
X5086 1 DigitalLDOLogic_VIA2 $T=146620 21220 0 0 $X=146150 $Y=20990
X5087 1 DigitalLDOLogic_VIA2 $T=146620 25300 0 0 $X=146150 $Y=25070
X5088 1 DigitalLDOLogic_VIA2 $T=146620 29380 0 0 $X=146150 $Y=29150
X5089 1 DigitalLDOLogic_VIA2 $T=146620 33460 0 0 $X=146150 $Y=33230
X5090 1 DigitalLDOLogic_VIA2 $T=146620 37540 0 0 $X=146150 $Y=37310
X5091 1 DigitalLDOLogic_VIA2 $T=146620 41620 0 0 $X=146150 $Y=41390
X5092 1 DigitalLDOLogic_VIA2 $T=146620 45700 0 0 $X=146150 $Y=45470
X5093 1 DigitalLDOLogic_VIA2 $T=146620 49780 0 0 $X=146150 $Y=49550
X5094 1 DigitalLDOLogic_VIA2 $T=146620 53860 0 0 $X=146150 $Y=53630
X5095 1 DigitalLDOLogic_VIA2 $T=146620 57940 0 0 $X=146150 $Y=57710
X5096 2 DigitalLDOLogic_VIA2 $T=150300 11700 0 0 $X=149830 $Y=11470
X5097 2 DigitalLDOLogic_VIA2 $T=150300 15780 0 0 $X=149830 $Y=15550
X5098 2 DigitalLDOLogic_VIA2 $T=150300 19860 0 0 $X=149830 $Y=19630
X5099 2 DigitalLDOLogic_VIA2 $T=150300 23940 0 0 $X=149830 $Y=23710
X5100 2 DigitalLDOLogic_VIA2 $T=150300 28020 0 0 $X=149830 $Y=27790
X5101 2 DigitalLDOLogic_VIA2 $T=150300 32100 0 0 $X=149830 $Y=31870
X5102 2 DigitalLDOLogic_VIA2 $T=150300 36180 0 0 $X=149830 $Y=35950
X5103 2 DigitalLDOLogic_VIA2 $T=150300 40260 0 0 $X=149830 $Y=40030
X5104 2 DigitalLDOLogic_VIA2 $T=150300 44340 0 0 $X=149830 $Y=44110
X5105 2 DigitalLDOLogic_VIA2 $T=150300 48420 0 0 $X=149830 $Y=48190
X5106 2 DigitalLDOLogic_VIA2 $T=150300 52500 0 0 $X=149830 $Y=52270
X5107 2 DigitalLDOLogic_VIA2 $T=150300 56580 0 0 $X=149830 $Y=56350
X5108 1 DigitalLDOLogic_VIA2 $T=152140 13060 0 0 $X=151670 $Y=12830
X5109 1 DigitalLDOLogic_VIA2 $T=152140 17140 0 0 $X=151670 $Y=16910
X5110 1 DigitalLDOLogic_VIA2 $T=152140 21220 0 0 $X=151670 $Y=20990
X5111 1 DigitalLDOLogic_VIA2 $T=152140 25300 0 0 $X=151670 $Y=25070
X5112 1 DigitalLDOLogic_VIA2 $T=152140 29380 0 0 $X=151670 $Y=29150
X5113 1 DigitalLDOLogic_VIA2 $T=152140 33460 0 0 $X=151670 $Y=33230
X5114 1 DigitalLDOLogic_VIA2 $T=152140 37540 0 0 $X=151670 $Y=37310
X5115 1 DigitalLDOLogic_VIA2 $T=152140 41620 0 0 $X=151670 $Y=41390
X5116 1 DigitalLDOLogic_VIA2 $T=152140 45700 0 0 $X=151670 $Y=45470
X5117 1 DigitalLDOLogic_VIA2 $T=152140 49780 0 0 $X=151670 $Y=49550
X5118 1 DigitalLDOLogic_VIA2 $T=152140 53860 0 0 $X=151670 $Y=53630
X5119 1 DigitalLDOLogic_VIA2 $T=152140 57940 0 0 $X=151670 $Y=57710
X5120 2 DigitalLDOLogic_VIA2 $T=155820 11700 0 0 $X=155350 $Y=11470
X5121 2 DigitalLDOLogic_VIA2 $T=155820 15780 0 0 $X=155350 $Y=15550
X5122 2 DigitalLDOLogic_VIA2 $T=155820 19860 0 0 $X=155350 $Y=19630
X5123 2 DigitalLDOLogic_VIA2 $T=155820 23940 0 0 $X=155350 $Y=23710
X5124 2 DigitalLDOLogic_VIA2 $T=155820 28020 0 0 $X=155350 $Y=27790
X5125 2 DigitalLDOLogic_VIA2 $T=155820 32100 0 0 $X=155350 $Y=31870
X5126 2 DigitalLDOLogic_VIA2 $T=155820 36180 0 0 $X=155350 $Y=35950
X5127 2 DigitalLDOLogic_VIA2 $T=155820 40260 0 0 $X=155350 $Y=40030
X5128 2 DigitalLDOLogic_VIA2 $T=155820 44340 0 0 $X=155350 $Y=44110
X5129 2 DigitalLDOLogic_VIA2 $T=155820 48420 0 0 $X=155350 $Y=48190
X5130 2 DigitalLDOLogic_VIA2 $T=155820 52500 0 0 $X=155350 $Y=52270
X5131 2 DigitalLDOLogic_VIA2 $T=155820 56580 0 0 $X=155350 $Y=56350
X5132 1 DigitalLDOLogic_VIA2 $T=157660 13060 0 0 $X=157190 $Y=12830
X5133 1 DigitalLDOLogic_VIA2 $T=157660 17140 0 0 $X=157190 $Y=16910
X5134 1 DigitalLDOLogic_VIA2 $T=157660 21220 0 0 $X=157190 $Y=20990
X5135 1 DigitalLDOLogic_VIA2 $T=157660 25300 0 0 $X=157190 $Y=25070
X5136 1 DigitalLDOLogic_VIA2 $T=157660 29380 0 0 $X=157190 $Y=29150
X5137 1 DigitalLDOLogic_VIA2 $T=157660 33460 0 0 $X=157190 $Y=33230
X5138 1 DigitalLDOLogic_VIA2 $T=157660 37540 0 0 $X=157190 $Y=37310
X5139 1 DigitalLDOLogic_VIA2 $T=157660 41620 0 0 $X=157190 $Y=41390
X5140 1 DigitalLDOLogic_VIA2 $T=157660 45700 0 0 $X=157190 $Y=45470
X5141 1 DigitalLDOLogic_VIA2 $T=157660 49780 0 0 $X=157190 $Y=49550
X5142 1 DigitalLDOLogic_VIA2 $T=157660 53860 0 0 $X=157190 $Y=53630
X5143 1 DigitalLDOLogic_VIA2 $T=157660 57940 0 0 $X=157190 $Y=57710
X5144 2 DigitalLDOLogic_VIA2 $T=161340 11700 0 0 $X=160870 $Y=11470
X5145 2 DigitalLDOLogic_VIA2 $T=161340 15780 0 0 $X=160870 $Y=15550
X5146 2 DigitalLDOLogic_VIA2 $T=161340 19860 0 0 $X=160870 $Y=19630
X5147 2 DigitalLDOLogic_VIA2 $T=161340 23940 0 0 $X=160870 $Y=23710
X5148 2 DigitalLDOLogic_VIA2 $T=161340 28020 0 0 $X=160870 $Y=27790
X5149 2 DigitalLDOLogic_VIA2 $T=161340 32100 0 0 $X=160870 $Y=31870
X5150 2 DigitalLDOLogic_VIA2 $T=161340 36180 0 0 $X=160870 $Y=35950
X5151 2 DigitalLDOLogic_VIA2 $T=161340 40260 0 0 $X=160870 $Y=40030
X5152 2 DigitalLDOLogic_VIA2 $T=161340 44340 0 0 $X=160870 $Y=44110
X5153 2 DigitalLDOLogic_VIA2 $T=161340 48420 0 0 $X=160870 $Y=48190
X5154 2 DigitalLDOLogic_VIA2 $T=161340 52500 0 0 $X=160870 $Y=52270
X5155 2 DigitalLDOLogic_VIA2 $T=161340 56580 0 0 $X=160870 $Y=56350
X5156 1 DigitalLDOLogic_VIA2 $T=163180 13060 0 0 $X=162710 $Y=12830
X5157 1 DigitalLDOLogic_VIA2 $T=163180 17140 0 0 $X=162710 $Y=16910
X5158 1 DigitalLDOLogic_VIA2 $T=163180 21220 0 0 $X=162710 $Y=20990
X5159 1 DigitalLDOLogic_VIA2 $T=163180 25300 0 0 $X=162710 $Y=25070
X5160 1 DigitalLDOLogic_VIA2 $T=163180 29380 0 0 $X=162710 $Y=29150
X5161 1 DigitalLDOLogic_VIA2 $T=163180 33460 0 0 $X=162710 $Y=33230
X5162 1 DigitalLDOLogic_VIA2 $T=163180 37540 0 0 $X=162710 $Y=37310
X5163 1 DigitalLDOLogic_VIA2 $T=163180 41620 0 0 $X=162710 $Y=41390
X5164 1 DigitalLDOLogic_VIA2 $T=163180 45700 0 0 $X=162710 $Y=45470
X5165 1 DigitalLDOLogic_VIA2 $T=163180 49780 0 0 $X=162710 $Y=49550
X5166 1 DigitalLDOLogic_VIA2 $T=163180 53860 0 0 $X=162710 $Y=53630
X5167 1 DigitalLDOLogic_VIA2 $T=163180 57940 0 0 $X=162710 $Y=57710
X5168 2 DigitalLDOLogic_VIA2 $T=166860 11700 0 0 $X=166390 $Y=11470
X5169 2 DigitalLDOLogic_VIA2 $T=166860 15780 0 0 $X=166390 $Y=15550
X5170 2 DigitalLDOLogic_VIA2 $T=166860 19860 0 0 $X=166390 $Y=19630
X5171 2 DigitalLDOLogic_VIA2 $T=166860 23940 0 0 $X=166390 $Y=23710
X5172 2 DigitalLDOLogic_VIA2 $T=166860 28020 0 0 $X=166390 $Y=27790
X5173 2 DigitalLDOLogic_VIA2 $T=166860 32100 0 0 $X=166390 $Y=31870
X5174 2 DigitalLDOLogic_VIA2 $T=166860 36180 0 0 $X=166390 $Y=35950
X5175 2 DigitalLDOLogic_VIA2 $T=166860 40260 0 0 $X=166390 $Y=40030
X5176 2 DigitalLDOLogic_VIA2 $T=166860 44340 0 0 $X=166390 $Y=44110
X5177 2 DigitalLDOLogic_VIA2 $T=166860 48420 0 0 $X=166390 $Y=48190
X5178 2 DigitalLDOLogic_VIA2 $T=166860 52500 0 0 $X=166390 $Y=52270
X5179 2 DigitalLDOLogic_VIA2 $T=166860 56580 0 0 $X=166390 $Y=56350
X5180 1 DigitalLDOLogic_VIA2 $T=168700 13060 0 0 $X=168230 $Y=12830
X5181 1 DigitalLDOLogic_VIA2 $T=168700 17140 0 0 $X=168230 $Y=16910
X5182 1 DigitalLDOLogic_VIA2 $T=168700 21220 0 0 $X=168230 $Y=20990
X5183 1 DigitalLDOLogic_VIA2 $T=168700 25300 0 0 $X=168230 $Y=25070
X5184 1 DigitalLDOLogic_VIA2 $T=168700 29380 0 0 $X=168230 $Y=29150
X5185 1 DigitalLDOLogic_VIA2 $T=168700 33460 0 0 $X=168230 $Y=33230
X5186 1 DigitalLDOLogic_VIA2 $T=168700 37540 0 0 $X=168230 $Y=37310
X5187 1 DigitalLDOLogic_VIA2 $T=168700 41620 0 0 $X=168230 $Y=41390
X5188 1 DigitalLDOLogic_VIA2 $T=168700 45700 0 0 $X=168230 $Y=45470
X5189 1 DigitalLDOLogic_VIA2 $T=168700 49780 0 0 $X=168230 $Y=49550
X5190 1 DigitalLDOLogic_VIA2 $T=168700 53860 0 0 $X=168230 $Y=53630
X5191 1 DigitalLDOLogic_VIA2 $T=168700 57940 0 0 $X=168230 $Y=57710
X5192 2 DigitalLDOLogic_VIA2 $T=172380 11700 0 0 $X=171910 $Y=11470
X5193 2 DigitalLDOLogic_VIA2 $T=172380 15780 0 0 $X=171910 $Y=15550
X5194 2 DigitalLDOLogic_VIA2 $T=172380 19860 0 0 $X=171910 $Y=19630
X5195 2 DigitalLDOLogic_VIA2 $T=172380 23940 0 0 $X=171910 $Y=23710
X5196 2 DigitalLDOLogic_VIA2 $T=172380 28020 0 0 $X=171910 $Y=27790
X5197 2 DigitalLDOLogic_VIA2 $T=172380 32100 0 0 $X=171910 $Y=31870
X5198 2 DigitalLDOLogic_VIA2 $T=172380 36180 0 0 $X=171910 $Y=35950
X5199 2 DigitalLDOLogic_VIA2 $T=172380 40260 0 0 $X=171910 $Y=40030
X5200 2 DigitalLDOLogic_VIA2 $T=172380 44340 0 0 $X=171910 $Y=44110
X5201 2 DigitalLDOLogic_VIA2 $T=172380 48420 0 0 $X=171910 $Y=48190
X5202 2 DigitalLDOLogic_VIA2 $T=172380 52500 0 0 $X=171910 $Y=52270
X5203 2 DigitalLDOLogic_VIA2 $T=172380 56580 0 0 $X=171910 $Y=56350
X5204 1 DigitalLDOLogic_VIA2 $T=174220 13060 0 0 $X=173750 $Y=12830
X5205 1 DigitalLDOLogic_VIA2 $T=174220 17140 0 0 $X=173750 $Y=16910
X5206 1 DigitalLDOLogic_VIA2 $T=174220 21220 0 0 $X=173750 $Y=20990
X5207 1 DigitalLDOLogic_VIA2 $T=174220 25300 0 0 $X=173750 $Y=25070
X5208 1 DigitalLDOLogic_VIA2 $T=174220 29380 0 0 $X=173750 $Y=29150
X5209 1 DigitalLDOLogic_VIA2 $T=174220 33460 0 0 $X=173750 $Y=33230
X5210 1 DigitalLDOLogic_VIA2 $T=174220 37540 0 0 $X=173750 $Y=37310
X5211 1 DigitalLDOLogic_VIA2 $T=174220 41620 0 0 $X=173750 $Y=41390
X5212 1 DigitalLDOLogic_VIA2 $T=174220 45700 0 0 $X=173750 $Y=45470
X5213 1 DigitalLDOLogic_VIA2 $T=174220 49780 0 0 $X=173750 $Y=49550
X5214 1 DigitalLDOLogic_VIA2 $T=174220 53860 0 0 $X=173750 $Y=53630
X5215 1 DigitalLDOLogic_VIA2 $T=174220 57940 0 0 $X=173750 $Y=57710
X5216 2 DigitalLDOLogic_VIA2 $T=177900 11700 0 0 $X=177430 $Y=11470
X5217 2 DigitalLDOLogic_VIA2 $T=177900 15780 0 0 $X=177430 $Y=15550
X5218 2 DigitalLDOLogic_VIA2 $T=177900 19860 0 0 $X=177430 $Y=19630
X5219 2 DigitalLDOLogic_VIA2 $T=177900 23940 0 0 $X=177430 $Y=23710
X5220 2 DigitalLDOLogic_VIA2 $T=177900 28020 0 0 $X=177430 $Y=27790
X5221 2 DigitalLDOLogic_VIA2 $T=177900 32100 0 0 $X=177430 $Y=31870
X5222 2 DigitalLDOLogic_VIA2 $T=177900 36180 0 0 $X=177430 $Y=35950
X5223 2 DigitalLDOLogic_VIA2 $T=177900 40260 0 0 $X=177430 $Y=40030
X5224 2 DigitalLDOLogic_VIA2 $T=177900 44340 0 0 $X=177430 $Y=44110
X5225 2 DigitalLDOLogic_VIA2 $T=177900 48420 0 0 $X=177430 $Y=48190
X5226 2 DigitalLDOLogic_VIA2 $T=177900 52500 0 0 $X=177430 $Y=52270
X5227 2 DigitalLDOLogic_VIA2 $T=177900 56580 0 0 $X=177430 $Y=56350
X5228 1 DigitalLDOLogic_VIA2 $T=179740 13060 0 0 $X=179270 $Y=12830
X5229 1 DigitalLDOLogic_VIA2 $T=179740 17140 0 0 $X=179270 $Y=16910
X5230 1 DigitalLDOLogic_VIA2 $T=179740 21220 0 0 $X=179270 $Y=20990
X5231 1 DigitalLDOLogic_VIA2 $T=179740 25300 0 0 $X=179270 $Y=25070
X5232 1 DigitalLDOLogic_VIA2 $T=179740 29380 0 0 $X=179270 $Y=29150
X5233 1 DigitalLDOLogic_VIA2 $T=179740 33460 0 0 $X=179270 $Y=33230
X5234 1 DigitalLDOLogic_VIA2 $T=179740 37540 0 0 $X=179270 $Y=37310
X5235 1 DigitalLDOLogic_VIA2 $T=179740 41620 0 0 $X=179270 $Y=41390
X5236 1 DigitalLDOLogic_VIA2 $T=179740 45700 0 0 $X=179270 $Y=45470
X5237 1 DigitalLDOLogic_VIA2 $T=179740 49780 0 0 $X=179270 $Y=49550
X5238 1 DigitalLDOLogic_VIA2 $T=179740 53860 0 0 $X=179270 $Y=53630
X5239 1 DigitalLDOLogic_VIA2 $T=179740 57940 0 0 $X=179270 $Y=57710
X5240 2 DigitalLDOLogic_VIA2 $T=183420 11700 0 0 $X=182950 $Y=11470
X5241 2 DigitalLDOLogic_VIA2 $T=183420 15780 0 0 $X=182950 $Y=15550
X5242 2 DigitalLDOLogic_VIA2 $T=183420 19860 0 0 $X=182950 $Y=19630
X5243 2 DigitalLDOLogic_VIA2 $T=183420 23940 0 0 $X=182950 $Y=23710
X5244 2 DigitalLDOLogic_VIA2 $T=183420 28020 0 0 $X=182950 $Y=27790
X5245 2 DigitalLDOLogic_VIA2 $T=183420 32100 0 0 $X=182950 $Y=31870
X5246 2 DigitalLDOLogic_VIA2 $T=183420 36180 0 0 $X=182950 $Y=35950
X5247 2 DigitalLDOLogic_VIA2 $T=183420 40260 0 0 $X=182950 $Y=40030
X5248 2 DigitalLDOLogic_VIA2 $T=183420 44340 0 0 $X=182950 $Y=44110
X5249 2 DigitalLDOLogic_VIA2 $T=183420 48420 0 0 $X=182950 $Y=48190
X5250 2 DigitalLDOLogic_VIA2 $T=183420 52500 0 0 $X=182950 $Y=52270
X5251 2 DigitalLDOLogic_VIA2 $T=183420 56580 0 0 $X=182950 $Y=56350
X5252 1 DigitalLDOLogic_VIA2 $T=185260 13060 0 0 $X=184790 $Y=12830
X5253 1 DigitalLDOLogic_VIA2 $T=185260 17140 0 0 $X=184790 $Y=16910
X5254 1 DigitalLDOLogic_VIA2 $T=185260 21220 0 0 $X=184790 $Y=20990
X5255 1 DigitalLDOLogic_VIA2 $T=185260 25300 0 0 $X=184790 $Y=25070
X5256 1 DigitalLDOLogic_VIA2 $T=185260 29380 0 0 $X=184790 $Y=29150
X5257 1 DigitalLDOLogic_VIA2 $T=185260 33460 0 0 $X=184790 $Y=33230
X5258 1 DigitalLDOLogic_VIA2 $T=185260 37540 0 0 $X=184790 $Y=37310
X5259 1 DigitalLDOLogic_VIA2 $T=185260 41620 0 0 $X=184790 $Y=41390
X5260 1 DigitalLDOLogic_VIA2 $T=185260 45700 0 0 $X=184790 $Y=45470
X5261 1 DigitalLDOLogic_VIA2 $T=185260 49780 0 0 $X=184790 $Y=49550
X5262 1 DigitalLDOLogic_VIA2 $T=185260 53860 0 0 $X=184790 $Y=53630
X5263 1 DigitalLDOLogic_VIA2 $T=185260 57940 0 0 $X=184790 $Y=57710
X5264 2 DigitalLDOLogic_VIA2 $T=188940 11700 0 0 $X=188470 $Y=11470
X5265 2 DigitalLDOLogic_VIA2 $T=188940 15780 0 0 $X=188470 $Y=15550
X5266 2 DigitalLDOLogic_VIA2 $T=188940 19860 0 0 $X=188470 $Y=19630
X5267 2 DigitalLDOLogic_VIA2 $T=188940 23940 0 0 $X=188470 $Y=23710
X5268 2 DigitalLDOLogic_VIA2 $T=188940 28020 0 0 $X=188470 $Y=27790
X5269 2 DigitalLDOLogic_VIA2 $T=188940 32100 0 0 $X=188470 $Y=31870
X5270 2 DigitalLDOLogic_VIA2 $T=188940 36180 0 0 $X=188470 $Y=35950
X5271 2 DigitalLDOLogic_VIA2 $T=188940 40260 0 0 $X=188470 $Y=40030
X5272 2 DigitalLDOLogic_VIA2 $T=188940 44340 0 0 $X=188470 $Y=44110
X5273 2 DigitalLDOLogic_VIA2 $T=188940 48420 0 0 $X=188470 $Y=48190
X5274 2 DigitalLDOLogic_VIA2 $T=188940 52500 0 0 $X=188470 $Y=52270
X5275 2 DigitalLDOLogic_VIA2 $T=188940 56580 0 0 $X=188470 $Y=56350
X5276 2 DigitalLDOLogic_VIA3 $T=12300 18500 0 0 $X=11590 $Y=17500
X5277 2 DigitalLDOLogic_VIA3 $T=12300 38900 0 0 $X=11590 $Y=37900
X5278 2 DigitalLDOLogic_VIA3 $T=17820 18500 0 0 $X=17110 $Y=17500
X5279 2 DigitalLDOLogic_VIA3 $T=17820 38900 0 0 $X=17110 $Y=37900
X5280 2 DigitalLDOLogic_VIA3 $T=23340 18500 0 0 $X=22630 $Y=17500
X5281 2 DigitalLDOLogic_VIA3 $T=23340 38900 0 0 $X=22630 $Y=37900
X5282 2 DigitalLDOLogic_VIA3 $T=28860 18500 0 0 $X=28150 $Y=17500
X5283 2 DigitalLDOLogic_VIA3 $T=28860 38900 0 0 $X=28150 $Y=37900
X5284 2 DigitalLDOLogic_VIA3 $T=34380 18500 0 0 $X=33670 $Y=17500
X5285 2 DigitalLDOLogic_VIA3 $T=34380 38900 0 0 $X=33670 $Y=37900
X5286 2 DigitalLDOLogic_VIA3 $T=39900 18500 0 0 $X=39190 $Y=17500
X5287 2 DigitalLDOLogic_VIA3 $T=39900 38900 0 0 $X=39190 $Y=37900
X5288 2 DigitalLDOLogic_VIA3 $T=45420 18500 0 0 $X=44710 $Y=17500
X5289 2 DigitalLDOLogic_VIA3 $T=45420 38900 0 0 $X=44710 $Y=37900
X5290 2 DigitalLDOLogic_VIA3 $T=50940 18500 0 0 $X=50230 $Y=17500
X5291 2 DigitalLDOLogic_VIA3 $T=50940 38900 0 0 $X=50230 $Y=37900
X5292 2 DigitalLDOLogic_VIA3 $T=56460 18500 0 0 $X=55750 $Y=17500
X5293 2 DigitalLDOLogic_VIA3 $T=56460 38900 0 0 $X=55750 $Y=37900
X5294 2 DigitalLDOLogic_VIA3 $T=61980 18500 0 0 $X=61270 $Y=17500
X5295 2 DigitalLDOLogic_VIA3 $T=61980 38900 0 0 $X=61270 $Y=37900
X5296 2 DigitalLDOLogic_VIA3 $T=67500 18500 0 0 $X=66790 $Y=17500
X5297 2 DigitalLDOLogic_VIA3 $T=67500 38900 0 0 $X=66790 $Y=37900
X5298 2 DigitalLDOLogic_VIA3 $T=73020 18500 0 0 $X=72310 $Y=17500
X5299 2 DigitalLDOLogic_VIA3 $T=73020 38900 0 0 $X=72310 $Y=37900
X5300 2 DigitalLDOLogic_VIA3 $T=78540 18500 0 0 $X=77830 $Y=17500
X5301 2 DigitalLDOLogic_VIA3 $T=78540 38900 0 0 $X=77830 $Y=37900
X5302 2 DigitalLDOLogic_VIA3 $T=84060 18500 0 0 $X=83350 $Y=17500
X5303 2 DigitalLDOLogic_VIA3 $T=84060 38900 0 0 $X=83350 $Y=37900
X5304 2 DigitalLDOLogic_VIA3 $T=89580 18500 0 0 $X=88870 $Y=17500
X5305 2 DigitalLDOLogic_VIA3 $T=89580 38900 0 0 $X=88870 $Y=37900
X5306 2 DigitalLDOLogic_VIA3 $T=95100 18500 0 0 $X=94390 $Y=17500
X5307 2 DigitalLDOLogic_VIA3 $T=95100 38900 0 0 $X=94390 $Y=37900
X5308 2 DigitalLDOLogic_VIA3 $T=100620 18500 0 0 $X=99910 $Y=17500
X5309 2 DigitalLDOLogic_VIA3 $T=100620 38900 0 0 $X=99910 $Y=37900
X5310 2 DigitalLDOLogic_VIA3 $T=106140 18500 0 0 $X=105430 $Y=17500
X5311 2 DigitalLDOLogic_VIA3 $T=106140 38900 0 0 $X=105430 $Y=37900
X5312 2 DigitalLDOLogic_VIA3 $T=111660 18500 0 0 $X=110950 $Y=17500
X5313 2 DigitalLDOLogic_VIA3 $T=111660 38900 0 0 $X=110950 $Y=37900
X5314 2 DigitalLDOLogic_VIA3 $T=117180 18500 0 0 $X=116470 $Y=17500
X5315 2 DigitalLDOLogic_VIA3 $T=117180 38900 0 0 $X=116470 $Y=37900
X5316 2 DigitalLDOLogic_VIA3 $T=122700 18500 0 0 $X=121990 $Y=17500
X5317 2 DigitalLDOLogic_VIA3 $T=122700 38900 0 0 $X=121990 $Y=37900
X5318 2 DigitalLDOLogic_VIA3 $T=128220 18500 0 0 $X=127510 $Y=17500
X5319 2 DigitalLDOLogic_VIA3 $T=128220 38900 0 0 $X=127510 $Y=37900
X5320 2 DigitalLDOLogic_VIA3 $T=133740 18500 0 0 $X=133030 $Y=17500
X5321 2 DigitalLDOLogic_VIA3 $T=133740 38900 0 0 $X=133030 $Y=37900
X5322 2 DigitalLDOLogic_VIA3 $T=139260 18500 0 0 $X=138550 $Y=17500
X5323 2 DigitalLDOLogic_VIA3 $T=139260 38900 0 0 $X=138550 $Y=37900
X5324 2 DigitalLDOLogic_VIA3 $T=144780 18500 0 0 $X=144070 $Y=17500
X5325 2 DigitalLDOLogic_VIA3 $T=144780 38900 0 0 $X=144070 $Y=37900
X5326 2 DigitalLDOLogic_VIA3 $T=150300 18500 0 0 $X=149590 $Y=17500
X5327 2 DigitalLDOLogic_VIA3 $T=150300 38900 0 0 $X=149590 $Y=37900
X5328 2 DigitalLDOLogic_VIA3 $T=155820 18500 0 0 $X=155110 $Y=17500
X5329 2 DigitalLDOLogic_VIA3 $T=155820 38900 0 0 $X=155110 $Y=37900
X5330 2 DigitalLDOLogic_VIA3 $T=161340 18500 0 0 $X=160630 $Y=17500
X5331 2 DigitalLDOLogic_VIA3 $T=161340 38900 0 0 $X=160630 $Y=37900
X5332 2 DigitalLDOLogic_VIA3 $T=166860 18500 0 0 $X=166150 $Y=17500
X5333 2 DigitalLDOLogic_VIA3 $T=166860 38900 0 0 $X=166150 $Y=37900
X5334 2 DigitalLDOLogic_VIA3 $T=172380 18500 0 0 $X=171670 $Y=17500
X5335 2 DigitalLDOLogic_VIA3 $T=172380 38900 0 0 $X=171670 $Y=37900
X5336 2 DigitalLDOLogic_VIA3 $T=177900 18500 0 0 $X=177190 $Y=17500
X5337 2 DigitalLDOLogic_VIA3 $T=177900 38900 0 0 $X=177190 $Y=37900
X5338 2 DigitalLDOLogic_VIA3 $T=183420 18500 0 0 $X=182710 $Y=17500
X5339 2 DigitalLDOLogic_VIA3 $T=183420 38900 0 0 $X=182710 $Y=37900
X5340 2 DigitalLDOLogic_VIA3 $T=188940 18500 0 0 $X=188230 $Y=17500
X5341 2 DigitalLDOLogic_VIA3 $T=188940 38900 0 0 $X=188230 $Y=37900
X5342 1 DigitalLDOLogic_VIA4 $T=12070 10110 0 0 $X=11820 $Y=9980
X5343 1 DigitalLDOLogic_VIA4 $T=14830 10110 0 0 $X=14580 $Y=9980
X5344 1 DigitalLDOLogic_VIA4 $T=17590 10110 0 0 $X=17340 $Y=9980
X5345 1 DigitalLDOLogic_VIA4 $T=20350 10110 0 0 $X=20100 $Y=9980
X5346 1 DigitalLDOLogic_VIA4 $T=23110 10110 0 0 $X=22860 $Y=9980
X5347 1 DigitalLDOLogic_VIA4 $T=25870 10110 0 0 $X=25620 $Y=9980
X5348 1 DigitalLDOLogic_VIA4 $T=28630 10110 0 0 $X=28380 $Y=9980
X5349 1 DigitalLDOLogic_VIA4 $T=31390 10110 0 0 $X=31140 $Y=9980
X5350 1 DigitalLDOLogic_VIA4 $T=34150 10110 0 0 $X=33900 $Y=9980
X5351 1 DigitalLDOLogic_VIA4 $T=36910 10110 0 0 $X=36660 $Y=9980
X5352 1 DigitalLDOLogic_VIA4 $T=39670 10110 0 0 $X=39420 $Y=9980
X5353 1 DigitalLDOLogic_VIA4 $T=42430 10110 0 0 $X=42180 $Y=9980
X5354 1 DigitalLDOLogic_VIA4 $T=45190 10110 0 0 $X=44940 $Y=9980
X5355 1 DigitalLDOLogic_VIA4 $T=47950 10110 0 0 $X=47700 $Y=9980
X5356 1 DigitalLDOLogic_VIA4 $T=50710 10110 0 0 $X=50460 $Y=9980
X5357 1 DigitalLDOLogic_VIA4 $T=53470 10110 0 0 $X=53220 $Y=9980
X5358 1 DigitalLDOLogic_VIA4 $T=56230 10110 0 0 $X=55980 $Y=9980
X5359 1 DigitalLDOLogic_VIA4 $T=58990 10110 0 0 $X=58740 $Y=9980
X5360 1 DigitalLDOLogic_VIA4 $T=61750 10110 0 0 $X=61500 $Y=9980
X5361 1 DigitalLDOLogic_VIA4 $T=64510 10110 0 0 $X=64260 $Y=9980
X5362 1 DigitalLDOLogic_VIA4 $T=67270 10110 0 0 $X=67020 $Y=9980
X5363 1 DigitalLDOLogic_VIA4 $T=70030 10110 0 0 $X=69780 $Y=9980
X5364 1 DigitalLDOLogic_VIA4 $T=72790 10110 0 0 $X=72540 $Y=9980
X5365 1 DigitalLDOLogic_VIA4 $T=75550 10110 0 0 $X=75300 $Y=9980
X5366 1 DigitalLDOLogic_VIA4 $T=78310 10110 0 0 $X=78060 $Y=9980
X5367 1 DigitalLDOLogic_VIA4 $T=81070 10110 0 0 $X=80820 $Y=9980
X5368 1 DigitalLDOLogic_VIA4 $T=83830 10110 0 0 $X=83580 $Y=9980
X5369 1 DigitalLDOLogic_VIA4 $T=86590 10110 0 0 $X=86340 $Y=9980
X5370 1 DigitalLDOLogic_VIA4 $T=89350 10110 0 0 $X=89100 $Y=9980
X5371 1 DigitalLDOLogic_VIA4 $T=92110 10110 0 0 $X=91860 $Y=9980
X5372 1 DigitalLDOLogic_VIA4 $T=94870 10110 0 0 $X=94620 $Y=9980
X5373 1 DigitalLDOLogic_VIA4 $T=97630 10110 0 0 $X=97380 $Y=9980
X5374 1 DigitalLDOLogic_VIA4 $T=100390 10110 0 0 $X=100140 $Y=9980
X5375 1 DigitalLDOLogic_VIA4 $T=103150 10110 0 0 $X=102900 $Y=9980
X5376 1 DigitalLDOLogic_VIA4 $T=105910 10110 0 0 $X=105660 $Y=9980
X5377 1 DigitalLDOLogic_VIA4 $T=108670 10110 0 0 $X=108420 $Y=9980
X5378 1 DigitalLDOLogic_VIA4 $T=111430 10110 0 0 $X=111180 $Y=9980
X5379 1 DigitalLDOLogic_VIA4 $T=114190 10110 0 0 $X=113940 $Y=9980
X5380 1 DigitalLDOLogic_VIA4 $T=116950 10110 0 0 $X=116700 $Y=9980
X5381 1 DigitalLDOLogic_VIA4 $T=119710 10110 0 0 $X=119460 $Y=9980
X5382 1 DigitalLDOLogic_VIA4 $T=122470 10110 0 0 $X=122220 $Y=9980
X5383 1 DigitalLDOLogic_VIA4 $T=125230 10110 0 0 $X=124980 $Y=9980
X5384 1 DigitalLDOLogic_VIA4 $T=127990 10110 0 0 $X=127740 $Y=9980
X5385 1 DigitalLDOLogic_VIA4 $T=130750 10110 0 0 $X=130500 $Y=9980
X5386 1 DigitalLDOLogic_VIA4 $T=133510 10110 0 0 $X=133260 $Y=9980
X5387 1 DigitalLDOLogic_VIA4 $T=136270 10110 0 0 $X=136020 $Y=9980
X5388 1 DigitalLDOLogic_VIA4 $T=139030 10110 0 0 $X=138780 $Y=9980
X5389 1 DigitalLDOLogic_VIA4 $T=141790 10110 0 0 $X=141540 $Y=9980
X5390 1 DigitalLDOLogic_VIA4 $T=144550 10110 0 0 $X=144300 $Y=9980
X5391 1 DigitalLDOLogic_VIA4 $T=147310 10110 0 0 $X=147060 $Y=9980
X5392 1 DigitalLDOLogic_VIA4 $T=150070 10110 0 0 $X=149820 $Y=9980
X5393 1 DigitalLDOLogic_VIA4 $T=152830 10110 0 0 $X=152580 $Y=9980
X5394 1 DigitalLDOLogic_VIA4 $T=155590 10110 0 0 $X=155340 $Y=9980
X5395 1 DigitalLDOLogic_VIA4 $T=158350 10110 0 0 $X=158100 $Y=9980
X5396 1 DigitalLDOLogic_VIA4 $T=161110 10110 0 0 $X=160860 $Y=9980
X5397 1 DigitalLDOLogic_VIA4 $T=163870 10110 0 0 $X=163620 $Y=9980
X5398 1 DigitalLDOLogic_VIA4 $T=166630 10110 0 0 $X=166380 $Y=9980
X5399 1 DigitalLDOLogic_VIA4 $T=169390 10110 0 0 $X=169140 $Y=9980
X5400 1 DigitalLDOLogic_VIA4 $T=172150 10110 0 0 $X=171900 $Y=9980
X5401 1 DigitalLDOLogic_VIA4 $T=174910 10110 0 0 $X=174660 $Y=9980
X5402 1 DigitalLDOLogic_VIA4 $T=177670 10110 0 0 $X=177420 $Y=9980
X5403 1 DigitalLDOLogic_VIA4 $T=180430 10110 0 0 $X=180180 $Y=9980
X5404 1 DigitalLDOLogic_VIA4 $T=183190 10110 0 0 $X=182940 $Y=9980
X5405 1 DigitalLDOLogic_VIA4 $T=185950 10110 0 0 $X=185700 $Y=9980
X5406 1 DigitalLDOLogic_VIA4 $T=188710 10110 0 0 $X=188460 $Y=9980
X5407 1 2 MASCO__Y3 $T=13430 24300 0 0 $X=13430 $Y=24300
X5408 1 2 MASCO__Y3 $T=13430 44700 0 0 $X=13430 $Y=44700
X5409 1 2 MASCO__Y3 $T=57590 24300 0 0 $X=57590 $Y=24300
X5410 1 2 MASCO__Y3 $T=57590 44700 0 0 $X=57590 $Y=44700
X5411 1 2 MASCO__Y3 $T=101750 24300 0 0 $X=101750 $Y=24300
X5412 1 2 MASCO__Y3 $T=101750 44700 0 0 $X=101750 $Y=44700
X5413 1 2 MASCO__Y3 $T=145910 24300 0 0 $X=145910 $Y=24300
X5414 1 2 MASCO__Y3 $T=145910 44700 0 0 $X=145910 $Y=44700
X5415 1 2 MASCO__B94 $T=29130 26080 0 0 $X=29130 $Y=26080
X5416 1 2 MASCO__B94 $T=29130 31520 0 0 $X=29130 $Y=31520
X5417 1 2 MASCO__B94 $T=29130 36960 0 0 $X=29130 $Y=36960
X5418 1 2 MASCO__B94 $T=29130 42400 0 0 $X=29130 $Y=42400
X5419 1 2 MASCO__B94 $T=29130 47840 0 0 $X=29130 $Y=47840
X5420 1 2 MASCO__B94 $T=29130 53280 0 0 $X=29130 $Y=53280
X5421 1 2 MASCO__B94 $T=58570 31520 0 0 $X=58570 $Y=31520
X5422 1 2 MASCO__B94 $T=58570 36960 0 0 $X=58570 $Y=36960
X5423 1 2 MASCO__B94 $T=58570 42400 0 0 $X=58570 $Y=42400
X5424 1 2 MASCO__B94 $T=58570 47840 0 0 $X=58570 $Y=47840
X5425 1 2 MASCO__B94 $T=58570 53280 0 0 $X=58570 $Y=53280
X5426 1 2 MASCO__B94 $T=88010 31520 0 0 $X=88010 $Y=31520
X5427 1 2 MASCO__B94 $T=88010 36960 0 0 $X=88010 $Y=36960
X5428 1 2 MASCO__B94 $T=88010 42400 0 0 $X=88010 $Y=42400
X5429 1 2 MASCO__B94 $T=88010 47840 0 0 $X=88010 $Y=47840
X5430 1 2 MASCO__B94 $T=88010 53280 0 0 $X=88010 $Y=53280
X5431 1 2 MASCO__B94 $T=102730 20640 0 0 $X=102730 $Y=20640
X5432 1 2 MASCO__B94 $T=146890 26080 0 0 $X=146890 $Y=26080
X5433 1 2 MASCO__B94 $T=176330 9760 0 0 $X=176330 $Y=9760
X5434 1 2 MASCO__B94 $T=176330 26080 0 0 $X=176330 $Y=26080
X5435 1 2 MASCO__B97 $T=25910 26080 0 0 $X=25910 $Y=26080
X5436 1 2 MASCO__B97 $T=25910 31520 0 0 $X=25910 $Y=31520
X5437 1 2 MASCO__B97 $T=25910 36960 0 0 $X=25910 $Y=36960
X5438 1 2 MASCO__B97 $T=25910 42400 0 0 $X=25910 $Y=42400
X5439 1 2 MASCO__B97 $T=25910 47840 0 0 $X=25910 $Y=47840
X5440 1 2 MASCO__B97 $T=25910 53280 0 0 $X=25910 $Y=53280
X5441 1 2 MASCO__B97 $T=84790 31520 0 0 $X=84790 $Y=31520
X5442 1 2 MASCO__B97 $T=84790 36960 0 0 $X=84790 $Y=36960
X5443 1 2 MASCO__B97 $T=84790 42400 0 0 $X=84790 $Y=42400
X5444 1 2 MASCO__B97 $T=84790 47840 0 0 $X=84790 $Y=47840
X5445 1 2 MASCO__B97 $T=84790 53280 0 0 $X=84790 $Y=53280
X5446 1 2 MASCO__B97 $T=114230 26080 0 0 $X=114230 $Y=26080
X5447 1 2 MASCO__B97 $T=114230 31520 0 0 $X=114230 $Y=31520
X5448 1 2 MASCO__B97 $T=114230 36960 0 0 $X=114230 $Y=36960
X5449 1 2 MASCO__B97 $T=114230 42400 0 0 $X=114230 $Y=42400
X5450 1 2 MASCO__B97 $T=114230 47840 0 0 $X=114230 $Y=47840
X5451 1 2 MASCO__B97 $T=114230 53280 0 0 $X=114230 $Y=53280
X5452 1 2 MASCO__B97 $T=173110 26080 0 0 $X=173110 $Y=26080
X5453 1 2 MASCO__B101 $T=13030 9760 0 0 $X=13030 $Y=9760
X5454 1 2 MASCO__B101 $T=13030 15200 0 0 $X=13030 $Y=15200
X5455 1 2 MASCO__B101 $T=13030 20640 0 0 $X=13030 $Y=20640
X5456 1 2 MASCO__B101 $T=13030 26080 0 0 $X=13030 $Y=26080
X5457 1 2 MASCO__B101 $T=13030 31520 0 0 $X=13030 $Y=31520
X5458 1 2 MASCO__B101 $T=13030 36960 0 0 $X=13030 $Y=36960
X5459 1 2 MASCO__B101 $T=13030 42400 0 0 $X=13030 $Y=42400
X5460 1 2 MASCO__B101 $T=13030 47840 0 0 $X=13030 $Y=47840
X5461 1 2 MASCO__B101 $T=13030 53280 0 0 $X=13030 $Y=53280
X5462 1 2 MASCO__B101 $T=42470 9760 0 0 $X=42470 $Y=9760
X5463 1 2 MASCO__B101 $T=42470 26080 0 0 $X=42470 $Y=26080
X5464 1 2 MASCO__B101 $T=42470 31520 0 0 $X=42470 $Y=31520
X5465 1 2 MASCO__B101 $T=42470 36960 0 0 $X=42470 $Y=36960
X5466 1 2 MASCO__B101 $T=42470 42400 0 0 $X=42470 $Y=42400
X5467 1 2 MASCO__B101 $T=42470 47840 0 0 $X=42470 $Y=47840
X5468 1 2 MASCO__B101 $T=42470 53280 0 0 $X=42470 $Y=53280
X5469 1 2 MASCO__B101 $T=71910 31520 0 0 $X=71910 $Y=31520
X5470 1 2 MASCO__B101 $T=71910 36960 0 0 $X=71910 $Y=36960
X5471 1 2 MASCO__B101 $T=71910 42400 0 0 $X=71910 $Y=42400
X5472 1 2 MASCO__B101 $T=71910 47840 0 0 $X=71910 $Y=47840
X5473 1 2 MASCO__B101 $T=71910 53280 0 0 $X=71910 $Y=53280
X5474 1 2 MASCO__B101 $T=101350 31520 0 0 $X=101350 $Y=31520
X5475 1 2 MASCO__B101 $T=101350 36960 0 0 $X=101350 $Y=36960
X5476 1 2 MASCO__B101 $T=101350 42400 0 0 $X=101350 $Y=42400
X5477 1 2 MASCO__B101 $T=101350 47840 0 0 $X=101350 $Y=47840
X5478 1 2 MASCO__B101 $T=101350 53280 0 0 $X=101350 $Y=53280
X5479 1 2 MASCO__B101 $T=130790 15200 0 0 $X=130790 $Y=15200
X5480 1 2 MASCO__B101 $T=160230 26080 0 0 $X=160230 $Y=26080
.ends DigitalLDOLogic

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_736670542250                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_736670542250 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_736670542250

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_736670542251                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_736670542251 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_736670542251

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_730310354533                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_730310354533 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=0
.ends nfet_01v8_CDNS_730310354533

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_730310354534                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_730310354534 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=1.6e-06 $X=0 $Y=0 $dt=1
.ends pfet_01v8_CDNS_730310354534

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nwellTap_CDNS_730310354531                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nwellTap_CDNS_730310354531 1
** N=1 EP=1 FDC=0
.ends nwellTap_CDNS_730310354531

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: subTap_CDNS_730310354532                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt subTap_CDNS_730310354532 1
** N=1 EP=1 FDC=0
.ends subTap_CDNS_730310354532

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inverter                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inverter 1 2 3 4
** N=4 EP=4 FDC=2
X0 3 L1M1_C_CDNS_736670542250 $T=2665 780 0 0 $X=2550 $Y=615
X1 2 L1M1_C_CDNS_736670542250 $T=2665 6690 0 0 $X=2550 $Y=6525
X2 4 L1M1_C_CDNS_736670542250 $T=3095 2830 0 0 $X=2980 $Y=2665
X3 2 M1M2_C_CDNS_736670542251 $T=-710 7295 0 0 $X=-840 $Y=6975
X4 3 M1M2_C_CDNS_736670542251 $T=5890 105 0 0 $X=5760 $Y=-215
X5 3 4 1 nfet_01v8_CDNS_730310354533 $T=2805 1285 0 0 $X=2540 $Y=1135
X6 2 4 1 pfet_01v8_CDNS_730310354534 $T=2805 4555 0 0 $X=2360 $Y=4375
X7 2 nwellTap_CDNS_730310354531 $T=2920 7265 0 0 $X=2475 $Y=6880
X8 3 subTap_CDNS_730310354532 $T=2735 130 0 0 $X=2440 $Y=-75
.ends inverter

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: polyConn_CDNS_729836244780                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt polyConn_CDNS_729836244780 1
** N=1 EP=1 FDC=0
.ends polyConn_CDNS_729836244780

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_729836244780                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_729836244780 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_729836244780

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_729836244781                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_729836244781 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_729836244781

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nwellTap_CDNS_729836244781                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nwellTap_CDNS_729836244781 1
** N=1 EP=1 FDC=0
.ends nwellTap_CDNS_729836244781

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nwellTap_CDNS_729836244782                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nwellTap_CDNS_729836244782 1
** N=1 EP=1 FDC=0
.ends nwellTap_CDNS_729836244782

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_729836244783                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_729836244783 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.5e-07 W=1.2e-06 $X=0 $Y=0 $dt=1
.ends pfet_01v8_CDNS_729836244783

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pass_transistors                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pass_transistors 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35
** N=35 EP=35 FDC=32
X0 1 polyConn_CDNS_729836244780 $T=2745 10060 0 0 $X=2610 $Y=9895
X1 2 polyConn_CDNS_729836244780 $T=3180 -2295 0 0 $X=3045 $Y=-2460
X2 3 polyConn_CDNS_729836244780 $T=3800 10050 0 0 $X=3665 $Y=9885
X3 4 polyConn_CDNS_729836244780 $T=4240 -2275 0 0 $X=4105 $Y=-2440
X4 5 polyConn_CDNS_729836244780 $T=4860 10060 0 0 $X=4725 $Y=9895
X5 6 polyConn_CDNS_729836244780 $T=5305 -2265 0 0 $X=5170 $Y=-2430
X6 7 polyConn_CDNS_729836244780 $T=5930 10065 0 0 $X=5795 $Y=9900
X7 8 polyConn_CDNS_729836244780 $T=6355 -2270 0 0 $X=6220 $Y=-2435
X8 9 polyConn_CDNS_729836244780 $T=6985 10070 0 0 $X=6850 $Y=9905
X9 10 polyConn_CDNS_729836244780 $T=7415 -2275 0 0 $X=7280 $Y=-2440
X10 11 polyConn_CDNS_729836244780 $T=8045 10070 0 0 $X=7910 $Y=9905
X11 12 polyConn_CDNS_729836244780 $T=8480 -2275 0 0 $X=8345 $Y=-2440
X12 13 polyConn_CDNS_729836244780 $T=9100 10070 0 0 $X=8965 $Y=9905
X13 14 polyConn_CDNS_729836244780 $T=9540 -2285 0 0 $X=9405 $Y=-2450
X14 15 polyConn_CDNS_729836244780 $T=10950 10065 0 0 $X=10815 $Y=9900
X15 16 polyConn_CDNS_729836244780 $T=11155 -2285 0 0 $X=11020 $Y=-2450
X16 17 polyConn_CDNS_729836244780 $T=12010 10075 0 0 $X=11875 $Y=9910
X17 18 polyConn_CDNS_729836244780 $T=12210 -2270 0 0 $X=12075 $Y=-2435
X18 19 polyConn_CDNS_729836244780 $T=13070 10075 0 0 $X=12935 $Y=9910
X19 20 polyConn_CDNS_729836244780 $T=13265 -2265 0 0 $X=13130 $Y=-2430
X20 21 polyConn_CDNS_729836244780 $T=14125 10090 0 0 $X=13990 $Y=9925
X21 22 polyConn_CDNS_729836244780 $T=14320 -2265 0 0 $X=14185 $Y=-2430
X22 23 polyConn_CDNS_729836244780 $T=15175 10080 0 0 $X=15040 $Y=9915
X23 24 polyConn_CDNS_729836244780 $T=15380 -2275 0 0 $X=15245 $Y=-2440
X24 25 polyConn_CDNS_729836244780 $T=16230 10080 0 0 $X=16095 $Y=9915
X25 26 polyConn_CDNS_729836244780 $T=16445 -2270 0 0 $X=16310 $Y=-2435
X26 27 polyConn_CDNS_729836244780 $T=18100 10090 0 0 $X=17965 $Y=9925
X27 28 polyConn_CDNS_729836244780 $T=18115 -2295 0 0 $X=17980 $Y=-2460
X28 29 polyConn_CDNS_729836244780 $T=19155 10080 0 0 $X=19020 $Y=9915
X29 30 polyConn_CDNS_729836244780 $T=19175 -2285 0 0 $X=19040 $Y=-2450
X30 31 polyConn_CDNS_729836244780 $T=20220 10080 0 0 $X=20085 $Y=9915
X31 32 polyConn_CDNS_729836244780 $T=20235 -2290 0 0 $X=20100 $Y=-2455
X32 33 M1M2_C_CDNS_729836244780 $T=485 12610 0 0 $X=355 $Y=12290
X33 33 M1M2_C_CDNS_729836244780 $T=490 285 0 0 $X=360 $Y=-35
X34 34 M1M2_C_CDNS_729836244780 $T=22800 13950 0 0 $X=22670 $Y=13630
X35 34 M1M2_C_CDNS_729836244780 $T=22865 1745 0 0 $X=22735 $Y=1425
X36 33 L1M1_C_CDNS_729836244781 $T=2480 12060 0 0 $X=2365 $Y=11895
X37 33 L1M1_C_CDNS_729836244781 $T=2915 -255 0 0 $X=2800 $Y=-420
X38 34 L1M1_C_CDNS_729836244781 $T=3010 13260 0 0 $X=2895 $Y=13095
X39 34 L1M1_C_CDNS_729836244781 $T=3445 1045 0 0 $X=3330 $Y=880
X40 33 L1M1_C_CDNS_729836244781 $T=3540 12065 0 0 $X=3425 $Y=11900
X41 3 L1M1_C_CDNS_729836244781 $T=3800 9600 0 0 $X=3685 $Y=9435
X42 33 L1M1_C_CDNS_729836244781 $T=3975 -255 0 0 $X=3860 $Y=-420
X43 34 L1M1_C_CDNS_729836244781 $T=4070 13275 0 0 $X=3955 $Y=13110
X44 4 L1M1_C_CDNS_729836244781 $T=4240 -2730 0 0 $X=4125 $Y=-2895
X45 34 L1M1_C_CDNS_729836244781 $T=4505 1055 0 0 $X=4390 $Y=890
X46 33 L1M1_C_CDNS_729836244781 $T=4600 12065 0 0 $X=4485 $Y=11900
X47 5 L1M1_C_CDNS_729836244781 $T=4860 9140 0 0 $X=4745 $Y=8975
X48 33 L1M1_C_CDNS_729836244781 $T=5035 -255 0 0 $X=4920 $Y=-420
X49 34 L1M1_C_CDNS_729836244781 $T=5130 13260 0 0 $X=5015 $Y=13095
X50 6 L1M1_C_CDNS_729836244781 $T=5305 -3175 0 0 $X=5190 $Y=-3340
X51 34 L1M1_C_CDNS_729836244781 $T=5565 1050 0 0 $X=5450 $Y=885
X52 33 L1M1_C_CDNS_729836244781 $T=5660 12080 0 0 $X=5545 $Y=11915
X53 7 L1M1_C_CDNS_729836244781 $T=5930 8685 0 0 $X=5815 $Y=8520
X54 33 L1M1_C_CDNS_729836244781 $T=6090 -255 0 0 $X=5975 $Y=-420
X55 34 L1M1_C_CDNS_729836244781 $T=6190 13265 0 0 $X=6075 $Y=13100
X56 8 L1M1_C_CDNS_729836244781 $T=6355 -3660 0 0 $X=6240 $Y=-3825
X57 34 L1M1_C_CDNS_729836244781 $T=6620 1050 0 0 $X=6505 $Y=885
X58 33 L1M1_C_CDNS_729836244781 $T=6720 12080 0 0 $X=6605 $Y=11915
X59 9 L1M1_C_CDNS_729836244781 $T=6985 8235 0 0 $X=6870 $Y=8070
X60 33 L1M1_C_CDNS_729836244781 $T=7150 -255 0 0 $X=7035 $Y=-420
X61 34 L1M1_C_CDNS_729836244781 $T=7250 13265 0 0 $X=7135 $Y=13100
X62 10 L1M1_C_CDNS_729836244781 $T=7415 -4105 0 0 $X=7300 $Y=-4270
X63 34 L1M1_C_CDNS_729836244781 $T=7680 1050 0 0 $X=7565 $Y=885
X64 33 L1M1_C_CDNS_729836244781 $T=7775 12085 0 0 $X=7660 $Y=11920
X65 11 L1M1_C_CDNS_729836244781 $T=8045 7760 0 0 $X=7930 $Y=7595
X66 33 L1M1_C_CDNS_729836244781 $T=8210 -255 0 0 $X=8095 $Y=-420
X67 34 L1M1_C_CDNS_729836244781 $T=8305 13265 0 0 $X=8190 $Y=13100
X68 12 L1M1_C_CDNS_729836244781 $T=8480 -4575 0 0 $X=8365 $Y=-4740
X69 34 L1M1_C_CDNS_729836244781 $T=8740 1050 0 0 $X=8625 $Y=885
X70 33 L1M1_C_CDNS_729836244781 $T=8830 12085 0 0 $X=8715 $Y=11920
X71 13 L1M1_C_CDNS_729836244781 $T=9100 7300 0 0 $X=8985 $Y=7135
X72 33 L1M1_C_CDNS_729836244781 $T=9270 -250 0 0 $X=9155 $Y=-415
X73 34 L1M1_C_CDNS_729836244781 $T=9360 13265 0 0 $X=9245 $Y=13100
X74 14 L1M1_C_CDNS_729836244781 $T=9540 -5050 0 0 $X=9425 $Y=-5215
X75 34 L1M1_C_CDNS_729836244781 $T=9800 1050 0 0 $X=9685 $Y=885
X76 33 L1M1_C_CDNS_729836244781 $T=10685 12075 0 0 $X=10570 $Y=11910
X77 33 L1M1_C_CDNS_729836244781 $T=10885 -255 0 0 $X=10770 $Y=-420
X78 15 L1M1_C_CDNS_729836244781 $T=10950 6805 0 0 $X=10835 $Y=6640
X79 16 L1M1_C_CDNS_729836244781 $T=11155 -5545 0 0 $X=11040 $Y=-5710
X80 34 L1M1_C_CDNS_729836244781 $T=11215 13255 0 0 $X=11100 $Y=13090
X81 34 L1M1_C_CDNS_729836244781 $T=11415 1050 0 0 $X=11300 $Y=885
X82 33 L1M1_C_CDNS_729836244781 $T=11745 12075 0 0 $X=11630 $Y=11910
X83 33 L1M1_C_CDNS_729836244781 $T=11940 -255 0 0 $X=11825 $Y=-420
X84 17 L1M1_C_CDNS_729836244781 $T=12010 6285 0 0 $X=11895 $Y=6120
X85 18 L1M1_C_CDNS_729836244781 $T=12210 -6055 0 0 $X=12095 $Y=-6220
X86 34 L1M1_C_CDNS_729836244781 $T=12275 13265 0 0 $X=12160 $Y=13100
X87 34 L1M1_C_CDNS_729836244781 $T=12470 1050 0 0 $X=12355 $Y=885
X88 33 L1M1_C_CDNS_729836244781 $T=12800 12075 0 0 $X=12685 $Y=11910
X89 33 L1M1_C_CDNS_729836244781 $T=12995 -255 0 0 $X=12880 $Y=-420
X90 19 L1M1_C_CDNS_729836244781 $T=13070 5735 0 0 $X=12955 $Y=5570
X91 20 L1M1_C_CDNS_729836244781 $T=13265 -6605 0 0 $X=13150 $Y=-6770
X92 34 L1M1_C_CDNS_729836244781 $T=13330 13265 0 0 $X=13215 $Y=13100
X93 34 L1M1_C_CDNS_729836244781 $T=13525 1050 0 0 $X=13410 $Y=885
X94 33 L1M1_C_CDNS_729836244781 $T=13855 12075 0 0 $X=13740 $Y=11910
X95 33 L1M1_C_CDNS_729836244781 $T=14055 -255 0 0 $X=13940 $Y=-420
X96 21 L1M1_C_CDNS_729836244781 $T=14125 5295 0 0 $X=14010 $Y=5130
X97 22 L1M1_C_CDNS_729836244781 $T=14320 -7055 0 0 $X=14205 $Y=-7220
X98 34 L1M1_C_CDNS_729836244781 $T=14385 13265 0 0 $X=14270 $Y=13100
X99 34 L1M1_C_CDNS_729836244781 $T=14585 1050 0 0 $X=14470 $Y=885
X100 33 L1M1_C_CDNS_729836244781 $T=14905 12065 0 0 $X=14790 $Y=11900
X101 33 L1M1_C_CDNS_729836244781 $T=15115 -260 0 0 $X=15000 $Y=-425
X102 23 L1M1_C_CDNS_729836244781 $T=15175 4755 0 0 $X=15060 $Y=4590
X103 24 L1M1_C_CDNS_729836244781 $T=15380 -7595 0 0 $X=15265 $Y=-7760
X104 34 L1M1_C_CDNS_729836244781 $T=15435 13260 0 0 $X=15320 $Y=13095
X105 34 L1M1_C_CDNS_729836244781 $T=15645 1045 0 0 $X=15530 $Y=880
X106 33 L1M1_C_CDNS_729836244781 $T=15965 12075 0 0 $X=15850 $Y=11910
X107 33 L1M1_C_CDNS_729836244781 $T=16175 -260 0 0 $X=16060 $Y=-425
X108 25 L1M1_C_CDNS_729836244781 $T=16230 4185 0 0 $X=16115 $Y=4020
X109 26 L1M1_C_CDNS_729836244781 $T=16445 -8160 0 0 $X=16330 $Y=-8325
X110 34 L1M1_C_CDNS_729836244781 $T=16495 13260 0 0 $X=16380 $Y=13095
X111 34 L1M1_C_CDNS_729836244781 $T=16705 1045 0 0 $X=16590 $Y=880
X112 33 L1M1_C_CDNS_729836244781 $T=17830 12075 0 0 $X=17715 $Y=11910
X113 33 L1M1_C_CDNS_729836244781 $T=17850 -260 0 0 $X=17735 $Y=-425
X114 27 L1M1_C_CDNS_729836244781 $T=18100 3650 0 0 $X=17985 $Y=3485
X115 28 L1M1_C_CDNS_729836244781 $T=18115 -8740 0 0 $X=18000 $Y=-8905
X116 34 L1M1_C_CDNS_729836244781 $T=18360 13255 0 0 $X=18245 $Y=13090
X117 34 L1M1_C_CDNS_729836244781 $T=18380 1020 0 0 $X=18265 $Y=855
X118 33 L1M1_C_CDNS_729836244781 $T=18890 12095 0 0 $X=18775 $Y=11930
X119 33 L1M1_C_CDNS_729836244781 $T=18910 -260 0 0 $X=18795 $Y=-425
X120 29 L1M1_C_CDNS_729836244781 $T=19155 3160 0 0 $X=19040 $Y=2995
X121 30 L1M1_C_CDNS_729836244781 $T=19175 -9235 0 0 $X=19060 $Y=-9400
X122 34 L1M1_C_CDNS_729836244781 $T=19420 13260 0 0 $X=19305 $Y=13095
X123 34 L1M1_C_CDNS_729836244781 $T=19440 1020 0 0 $X=19325 $Y=855
X124 33 L1M1_C_CDNS_729836244781 $T=19950 12080 0 0 $X=19835 $Y=11915
X125 33 L1M1_C_CDNS_729836244781 $T=19965 -260 0 0 $X=19850 $Y=-425
X126 31 L1M1_C_CDNS_729836244781 $T=20220 2685 0 0 $X=20105 $Y=2520
X127 32 L1M1_C_CDNS_729836244781 $T=20235 -9705 0 0 $X=20120 $Y=-9870
X128 34 L1M1_C_CDNS_729836244781 $T=20480 13240 0 0 $X=20365 $Y=13075
X129 34 L1M1_C_CDNS_729836244781 $T=20495 1020 0 0 $X=20380 $Y=855
X130 33 nwellTap_CDNS_729836244781 $T=1780 12560 0 0 $X=1335 $Y=12175
X131 33 nwellTap_CDNS_729836244781 $T=2175 195 0 0 $X=1730 $Y=-190
X132 33 nwellTap_CDNS_729836244781 $T=21155 12545 0 0 $X=20710 $Y=12160
X133 33 nwellTap_CDNS_729836244781 $T=21200 -5 0 0 $X=20755 $Y=-390
X134 33 nwellTap_CDNS_729836244782 $T=10020 11065 0 0 $X=9755 $Y=10500
X135 33 nwellTap_CDNS_729836244782 $T=10390 -1250 0 0 $X=10125 $Y=-1815
X136 33 nwellTap_CDNS_729836244782 $T=17170 11125 0 0 $X=16905 $Y=10560
X137 33 nwellTap_CDNS_729836244782 $T=17300 -1255 0 0 $X=17035 $Y=-1820
X138 33 34 1 pfet_01v8_CDNS_729836244783 $T=2620 10485 0 0 $X=2175 $Y=10305
X139 33 34 2 pfet_01v8_CDNS_729836244783 $T=3055 -1865 0 0 $X=2610 $Y=-2045
X140 33 34 3 pfet_01v8_CDNS_729836244783 $T=3680 10485 0 0 $X=3235 $Y=10305
X141 33 34 4 pfet_01v8_CDNS_729836244783 $T=4115 -1865 0 0 $X=3670 $Y=-2045
X142 33 34 5 pfet_01v8_CDNS_729836244783 $T=4740 10485 0 0 $X=4295 $Y=10305
X143 33 34 6 pfet_01v8_CDNS_729836244783 $T=5175 -1865 0 0 $X=4730 $Y=-2045
X144 33 34 7 pfet_01v8_CDNS_729836244783 $T=5800 10485 0 0 $X=5355 $Y=10305
X145 33 34 8 pfet_01v8_CDNS_729836244783 $T=6230 -1865 0 0 $X=5785 $Y=-2045
X146 33 34 9 pfet_01v8_CDNS_729836244783 $T=6860 10485 0 0 $X=6415 $Y=10305
X147 33 34 10 pfet_01v8_CDNS_729836244783 $T=7290 -1865 0 0 $X=6845 $Y=-2045
X148 33 34 11 pfet_01v8_CDNS_729836244783 $T=7915 10485 0 0 $X=7470 $Y=10305
X149 33 34 12 pfet_01v8_CDNS_729836244783 $T=8350 -1865 0 0 $X=7905 $Y=-2045
X150 33 34 13 pfet_01v8_CDNS_729836244783 $T=8970 10485 0 0 $X=8525 $Y=10305
X151 33 34 14 pfet_01v8_CDNS_729836244783 $T=9410 -1865 0 0 $X=8965 $Y=-2045
X152 33 34 15 pfet_01v8_CDNS_729836244783 $T=10825 10485 0 0 $X=10380 $Y=10305
X153 33 34 16 pfet_01v8_CDNS_729836244783 $T=11025 -1865 0 0 $X=10580 $Y=-2045
X154 33 34 17 pfet_01v8_CDNS_729836244783 $T=11885 10485 0 0 $X=11440 $Y=10305
X155 33 34 18 pfet_01v8_CDNS_729836244783 $T=12080 -1865 0 0 $X=11635 $Y=-2045
X156 33 34 19 pfet_01v8_CDNS_729836244783 $T=12940 10485 0 0 $X=12495 $Y=10305
X157 33 34 20 pfet_01v8_CDNS_729836244783 $T=13135 -1865 0 0 $X=12690 $Y=-2045
X158 33 34 21 pfet_01v8_CDNS_729836244783 $T=13995 10485 0 0 $X=13550 $Y=10305
X159 33 34 22 pfet_01v8_CDNS_729836244783 $T=14195 -1865 0 0 $X=13750 $Y=-2045
X160 33 34 23 pfet_01v8_CDNS_729836244783 $T=15045 10480 0 0 $X=14600 $Y=10300
X161 33 34 24 pfet_01v8_CDNS_729836244783 $T=15255 -1870 0 0 $X=14810 $Y=-2050
X162 33 34 25 pfet_01v8_CDNS_729836244783 $T=16105 10480 0 0 $X=15660 $Y=10300
X163 33 34 26 pfet_01v8_CDNS_729836244783 $T=16315 -1870 0 0 $X=15870 $Y=-2050
X164 33 34 27 pfet_01v8_CDNS_729836244783 $T=17970 10480 0 0 $X=17525 $Y=10300
X165 33 34 28 pfet_01v8_CDNS_729836244783 $T=17990 -1870 0 0 $X=17545 $Y=-2050
X166 33 34 29 pfet_01v8_CDNS_729836244783 $T=19030 10480 0 0 $X=18585 $Y=10300
X167 33 34 30 pfet_01v8_CDNS_729836244783 $T=19050 -1870 0 0 $X=18605 $Y=-2050
X168 33 34 31 pfet_01v8_CDNS_729836244783 $T=20090 10480 0 0 $X=19645 $Y=10300
X169 33 34 32 pfet_01v8_CDNS_729836244783 $T=20105 -1870 0 0 $X=19660 $Y=-2050
.ends pass_transistors

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_736669032860                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_736669032860 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_736669032860

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_736669032861                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_736669032861 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_736669032861

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_730309971733                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_730309971733 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=1
.ends pfet_01v8_CDNS_730309971733

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_730309971734                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_730309971734 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=0
.ends nfet_01v8_CDNS_730309971734

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_730309971735                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_730309971735 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=1.6e-06 $X=0 $Y=0 $dt=1
.ends pfet_01v8_CDNS_730309971735

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: polyConn_CDNS_730309971730                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt polyConn_CDNS_730309971730 1
** N=1 EP=1 FDC=0
.ends polyConn_CDNS_730309971730

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nwellTap_CDNS_730309971731                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nwellTap_CDNS_730309971731 1
** N=1 EP=1 FDC=0
.ends nwellTap_CDNS_730309971731

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: subTap_CDNS_730309971732                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt subTap_CDNS_730309971732 1
** N=1 EP=1 FDC=0
.ends subTap_CDNS_730309971732

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rs_latch_new                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rs_latch_new 1 2 3 4 5 6
** N=8 EP=6 FDC=8
X0 6 L1M1_C_CDNS_736669032860 $T=1035 -1950 0 0 $X=920 $Y=-2115
X1 5 L1M1_C_CDNS_736669032860 $T=1035 3960 0 0 $X=920 $Y=3795
X2 7 L1M1_C_CDNS_736669032860 $T=1465 100 0 0 $X=1350 $Y=-65
X3 6 L1M1_C_CDNS_736669032860 $T=3435 -2000 0 0 $X=3320 $Y=-2165
X4 5 L1M1_C_CDNS_736669032860 $T=3435 4050 0 0 $X=3320 $Y=3885
X5 3 L1M1_C_CDNS_736669032860 $T=3865 2045 0 0 $X=3750 $Y=1880
X6 6 L1M1_C_CDNS_736669032860 $T=6430 -2010 0 0 $X=6315 $Y=-2175
X7 5 L1M1_C_CDNS_736669032860 $T=6430 4075 0 0 $X=6315 $Y=3910
X8 2 L1M1_C_CDNS_736669032860 $T=6860 1595 0 0 $X=6745 $Y=1430
X9 6 L1M1_C_CDNS_736669032860 $T=8840 -1950 0 0 $X=8725 $Y=-2115
X10 5 L1M1_C_CDNS_736669032860 $T=8840 3960 0 0 $X=8725 $Y=3795
X11 8 L1M1_C_CDNS_736669032860 $T=9270 105 0 0 $X=9155 $Y=-60
X12 5 M1M2_C_CDNS_736669032861 $T=-1945 4595 0 0 $X=-2075 $Y=4275
X13 6 M1M2_C_CDNS_736669032861 $T=13505 -2615 0 0 $X=13375 $Y=-2935
X14 5 3 2 pfet_01v8_CDNS_730309971733 $T=3575 2425 0 0 $X=3130 $Y=2245
X15 5 2 3 pfet_01v8_CDNS_730309971733 $T=6570 2425 0 0 $X=6125 $Y=2245
X16 6 7 1 nfet_01v8_CDNS_730309971734 $T=1175 -1445 0 0 $X=910 $Y=-1595
X17 6 3 7 nfet_01v8_CDNS_730309971734 $T=3575 -1455 0 0 $X=3310 $Y=-1605
X18 6 2 8 nfet_01v8_CDNS_730309971734 $T=6570 -1455 0 0 $X=6305 $Y=-1605
X19 6 8 4 nfet_01v8_CDNS_730309971734 $T=8980 -1445 0 0 $X=8715 $Y=-1595
X20 5 7 1 pfet_01v8_CDNS_730309971735 $T=1175 1825 0 0 $X=730 $Y=1645
X21 5 8 4 pfet_01v8_CDNS_730309971735 $T=8980 1825 0 0 $X=8535 $Y=1645
X22 1 polyConn_CDNS_730309971730 $T=640 830 0 0 $X=505 $Y=665
X23 7 polyConn_CDNS_730309971730 $T=3230 100 0 0 $X=3095 $Y=-65
X24 2 polyConn_CDNS_730309971730 $T=4295 1595 0 0 $X=4160 $Y=1430
X25 3 polyConn_CDNS_730309971730 $T=6190 2045 0 0 $X=6055 $Y=1880
X26 8 polyConn_CDNS_730309971730 $T=7500 105 0 0 $X=7365 $Y=-60
X27 4 polyConn_CDNS_730309971730 $T=10025 980 0 0 $X=9890 $Y=815
X28 5 nwellTap_CDNS_730309971731 $T=2460 2925 0 0 $X=2195 $Y=2360
X29 5 nwellTap_CDNS_730309971731 $T=7840 2925 0 0 $X=7575 $Y=2360
X30 6 subTap_CDNS_730309971732 $T=2480 -955 0 0 $X=2365 $Y=-1340
X31 6 subTap_CDNS_730309971732 $T=7880 -970 0 0 $X=7765 $Y=-1355
.ends rs_latch_new

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ptap_tile                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ptap_tile 1
** N=1 EP=1 FDC=0
.ends ptap_tile

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ntap_tile                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ntap_tile 1
** N=1 EP=1 FDC=0
.ends ntap_tile

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=6.5e-06 $X=570 $Y=0 $dt=0
M1 1 3 2 4 nfet_01v8 L=1.5e-07 W=6.5e-06 $X=1000 $Y=0 $dt=0
.ends two_finger_mos_tile

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile_1                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile_1 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1e-06 $X=570 $Y=0 $dt=0
M1 1 3 2 4 nfet_01v8 L=1.5e-07 W=1e-06 $X=1000 $Y=0 $dt=0
.ends two_finger_mos_tile_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile_2                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile_2 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1.1e-05 $X=570 $Y=0 $dt=0
M1 1 3 2 4 nfet_01v8 L=1.5e-07 W=1.1e-05 $X=1000 $Y=0 $dt=0
.ends two_finger_mos_tile_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile_3                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile_3 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 pfet_01v8 L=1.5e-07 W=1e-06 $X=570 $Y=0 $dt=1
M1 1 3 2 4 pfet_01v8 L=1.5e-07 W=1e-06 $X=1000 $Y=0 $dt=1
.ends two_finger_mos_tile_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile_4                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile_4 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 pfet_01v8 L=1.5e-07 W=4.2e-07 $X=570 $Y=0 $dt=1
M1 1 3 2 4 pfet_01v8 L=1.5e-07 W=4.2e-07 $X=1000 $Y=0 $dt=1
.ends two_finger_mos_tile_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: strong_arm_half                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt strong_arm_half 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 FDC=36
X0 3 ptap_tile $T=0 -35640 0 0 $X=-205 $Y=-35790
X1 4 ntap_tile $T=0 0 0 0 $X=-430 $Y=-540
X2 3 3 3 3 two_finger_mos_tile $T=-430 -32940 0 0 $X=-215 $Y=-34175
X3 3 6 5 3 two_finger_mos_tile $T=1290 -32940 0 0 $X=1505 $Y=-34175
X4 3 6 5 3 two_finger_mos_tile $T=3010 -32940 0 0 $X=3225 $Y=-34175
X5 3 3 3 3 two_finger_mos_tile_1 $T=-430 -24300 0 0 $X=-215 $Y=-25535
X6 6 7 8 3 two_finger_mos_tile_1 $T=1290 -24300 0 0 $X=1505 $Y=-25535
X7 6 9 10 3 two_finger_mos_tile_1 $T=3010 -24300 0 0 $X=3225 $Y=-25535
X8 3 3 3 3 two_finger_mos_tile_2 $T=-430 -21060 0 0 $X=-215 $Y=-22295
X9 7 1 2 3 two_finger_mos_tile_2 $T=1290 -21060 0 0 $X=1505 $Y=-22295
X10 9 2 1 3 two_finger_mos_tile_2 $T=3010 -21060 0 0 $X=3225 $Y=-22295
X11 4 4 4 4 two_finger_mos_tile_3 $T=-430 -7560 0 0 $X=-430 $Y=-9180
X12 4 1 2 4 two_finger_mos_tile_3 $T=1290 -7560 0 0 $X=1290 $Y=-9180
X13 4 2 1 4 two_finger_mos_tile_3 $T=3010 -7560 0 0 $X=3010 $Y=-9180
X14 4 4 4 4 two_finger_mos_tile_4 $T=-430 -4320 0 0 $X=-430 $Y=-5940
X15 4 4 4 4 two_finger_mos_tile_4 $T=-430 -1620 0 0 $X=-430 $Y=-3240
X16 4 7 5 4 two_finger_mos_tile_4 $T=1290 -4320 0 0 $X=1290 $Y=-5940
X17 4 1 5 4 two_finger_mos_tile_4 $T=1290 -1620 0 0 $X=1290 $Y=-3240
X18 4 9 5 4 two_finger_mos_tile_4 $T=3010 -4320 0 0 $X=3010 $Y=-5940
X19 4 2 5 4 two_finger_mos_tile_4 $T=3010 -1620 0 0 $X=3010 $Y=-3240
.ends strong_arm_half

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: strong_arm                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt strong_arm 1 2 3 4 5 6 7
** N=11 EP=7 FDC=72
X0 6 4 1 2 7 8 9 3 10 5 strong_arm_half $T=0 0 0 0 $X=-430 $Y=-35790
X1 6 4 1 2 7 8 9 3 11 5 strong_arm_half $T=9460 0 1 180 $X=4730 $Y=-35790
.ends strong_arm

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__mux2_1                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__mux2_1 1 2 3 4 5 6 7 8
** N=18 EP=8 FDC=12
M0 3 9 1 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=395 $Y=235 $dt=0
M1 13 4 3 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=940 $Y=235 $dt=0
M2 9 5 13 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1420 $Y=235 $dt=0
M3 14 6 9 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=2045 $Y=235 $dt=0
M4 3 10 14 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=2525 $Y=235 $dt=0
M5 10 4 3 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=3365 $Y=235 $dt=0
M6 2 9 1 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=395 $Y=1485 $dt=2
M7 11 4 2 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=940 $Y=1870 $dt=2
M8 9 6 11 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=1455 $Y=1870 $dt=2
M9 12 5 9 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=2525 $Y=1870 $dt=2
M10 2 10 12 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=2885 $Y=1870 $dt=2
M11 10 4 2 8 pfet_01v8_hvt L=1.5e-07 W=4.2e-07 $X=3365 $Y=1870 $dt=2
.ends sky130_fd_sc_hd__mux2_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__mux2_2                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__mux2_2 1 2 3 4 5 6 7 8
** N=18 EP=8 FDC=14
M0 1 9 3 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=395 $Y=235 $dt=0
M1 3 9 1 7 nfet_01v8 L=1.5e-07 W=6.5e-07 $X=815 $Y=235 $dt=0
M2 13 10 3 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1290 $Y=235 $dt=0
M3 9 4 13 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=1765 $Y=235 $dt=0
M4 14 5 9 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=2740 $Y=235 $dt=0
M5 3 6 14 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=3165 $Y=235 $dt=0
M6 10 6 3 7 nfet_01v8 L=1.5e-07 W=4.2e-07 $X=3585 $Y=235 $dt=0
M7 1 9 2 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=395 $Y=1485 $dt=2
M8 2 9 1 8 pfet_01v8_hvt L=1.5e-07 W=1e-06 $X=815 $Y=1485 $dt=2
M9 11 10 2 8 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=1380 $Y=1845 $dt=2
M10 9 5 11 8 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=2245 $Y=1845 $dt=2
M11 12 4 9 8 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=2805 $Y=1845 $dt=2
M12 2 6 12 8 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=3165 $Y=1845 $dt=2
M13 10 6 2 8 pfet_01v8_hvt L=1.5e-07 W=6.4e-07 $X=3585 $Y=1845 $dt=2
.ends sky130_fd_sc_hd__mux2_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__tap_1                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__tap_1 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__tap_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__tapvpwrvgnd_1                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 1 2
** N=2 EP=2 FDC=0
.ends sky130_fd_sc_hd__tapvpwrvgnd_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_6                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_6 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=1.97e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=1.97e-06 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_3                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_3 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=5.9e-07 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=5.9e-07 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_12                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_12 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=4.73e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=4.73e-06 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_4                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_4 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=1.05e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=1.05e-06 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__decap_8                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__decap_8 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 1 2 3 nfet_01v8 L=2.89e-06 W=5.5e-07 $X=395 $Y=235 $dt=0
M1 1 2 1 4 pfet_01v8_hvt L=2.89e-06 W=8.7e-07 $X=395 $Y=1615 $dt=2
.ends sky130_fd_sc_hd__decap_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__fill_2                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__fill_2 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__fill_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: sky130_fd_sc_hd__fill_1                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt sky130_fd_sc_hd__fill_1 1 2 3 4
** N=4 EP=4 FDC=0
.ends sky130_fd_sc_hd__fill_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2M3_PR                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2M3_PR 1
** N=1 EP=1 FDC=0
.ends M2M3_PR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_PR                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_PR 1
** N=1 EP=1 FDC=0
.ends M1M2_PR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_PR                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_PR 1
** N=1 EP=1 FDC=0
.ends L1M1_PR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3M4_PR                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3M4_PR 1
** N=1 EP=1 FDC=0
.ends M3M4_PR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA0                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA0 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA1                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA1 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA2                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA2 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA3                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA3 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA4                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA4 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA5                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA5 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA7                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA7 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA8                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA8 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA9                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA9 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA10                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA10 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA11                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA11 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA12                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA12 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA13                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA13 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA15                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA15 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA16                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA16 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top_VIA18                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top_VIA18 1
** N=1 EP=1 FDC=0
.ends digital_ldo_top_VIA18

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y1 1
** N=1 EP=1 FDC=0
X0 1 digital_ldo_top_VIA12 $T=710 1000 0 0 $X=0 $Y=0
X1 1 digital_ldo_top_VIA12 $T=6230 1000 0 0 $X=5520 $Y=0
X2 1 digital_ldo_top_VIA12 $T=11750 1000 0 0 $X=11040 $Y=0
X3 1 digital_ldo_top_VIA12 $T=17270 1000 0 0 $X=16560 $Y=0
X4 1 digital_ldo_top_VIA12 $T=22790 1000 0 0 $X=22080 $Y=0
X5 1 digital_ldo_top_VIA12 $T=28310 1000 0 0 $X=27600 $Y=0
X6 1 digital_ldo_top_VIA12 $T=33830 1000 0 0 $X=33120 $Y=0
.ends MASCO__Y1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y2 1
** N=1 EP=1 FDC=0
X0 1 digital_ldo_top_VIA12 $T=710 1000 0 0 $X=0 $Y=0
X1 1 digital_ldo_top_VIA12 $T=6230 1000 0 0 $X=5520 $Y=0
X2 1 digital_ldo_top_VIA12 $T=11750 1000 0 0 $X=11040 $Y=0
X3 1 digital_ldo_top_VIA12 $T=17270 1000 0 0 $X=16560 $Y=0
X4 1 digital_ldo_top_VIA12 $T=22790 1000 0 0 $X=22080 $Y=0
X5 1 digital_ldo_top_VIA12 $T=28310 1000 0 0 $X=27600 $Y=0
X6 1 digital_ldo_top_VIA12 $T=33830 1000 0 0 $X=33120 $Y=0
X7 1 digital_ldo_top_VIA12 $T=39350 1000 0 0 $X=38640 $Y=0
X8 1 digital_ldo_top_VIA12 $T=44870 1000 0 0 $X=44160 $Y=0
X9 1 digital_ldo_top_VIA12 $T=50390 1000 0 0 $X=49680 $Y=0
X10 1 digital_ldo_top_VIA12 $T=55910 1000 0 0 $X=55200 $Y=0
X11 1 digital_ldo_top_VIA12 $T=61430 1000 0 0 $X=60720 $Y=0
.ends MASCO__Y2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B31                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B31 1 2
** N=2 EP=2 FDC=4
X0 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=1570 2960 1 0 $X=1380 $Y=0
X1 1 2 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=1570 2960 0 0 $X=1380 $Y=2720
X2 1 2 2 1 sky130_fd_sc_hd__decap_3 $T=190 2960 1 0 $X=0 $Y=0
X3 1 2 2 1 sky130_fd_sc_hd__decap_3 $T=190 2960 0 0 $X=0 $Y=2720
.ends MASCO__B31

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B32                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B32 1 2
** N=2 EP=2 FDC=8
X0 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 2960 1 0 $X=0 $Y=0
X1 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 2960 0 0 $X=0 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_8 $T=5710 2960 1 0 $X=5520 $Y=0
X3 2 1 1 2 sky130_fd_sc_hd__decap_8 $T=5710 2960 0 0 $X=5520 $Y=2720
.ends MASCO__B32

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B33                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B33 1 2
** N=2 EP=2 FDC=4
X0 2 1 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=190 240 0 0 $X=0 $Y=0
X1 2 1 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=190 5680 1 0 $X=0 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=650 240 0 0 $X=460 $Y=0
X3 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=650 5680 1 0 $X=460 $Y=2720
.ends MASCO__B33

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B35                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B35 1 2
** N=2 EP=2 FDC=8
X0 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 2960 1 0 $X=0 $Y=0
X1 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 2960 0 0 $X=0 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=5710 2960 1 0 $X=5520 $Y=0
X3 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=5710 2960 0 0 $X=5520 $Y=2720
.ends MASCO__B35

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B37                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B37 1 2
** N=2 EP=2 FDC=4
X0 2 1 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=190 2960 1 0 $X=0 $Y=0
X1 2 1 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=190 2960 0 0 $X=0 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=650 2960 1 0 $X=460 $Y=0
X3 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=650 2960 0 0 $X=460 $Y=2720
.ends MASCO__B37

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B39                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B39 1 2
** N=2 EP=2 FDC=4
X0 2 1 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=1570 240 0 0 $X=1380 $Y=0
X1 2 1 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=1570 5680 1 0 $X=1380 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=190 240 0 0 $X=0 $Y=0
X3 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=190 5680 1 0 $X=0 $Y=2720
.ends MASCO__B39

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B40                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B40 1 2
** N=2 EP=2 FDC=8
X0 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 240 0 0 $X=0 $Y=0
X1 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 5680 1 0 $X=0 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=5710 240 0 0 $X=5520 $Y=0
X3 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=5710 5680 1 0 $X=5520 $Y=2720
.ends MASCO__B40

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B63                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B63 1 2
** N=2 EP=2 FDC=32
X0 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=13070 240 0 0 $X=12880 $Y=0
X1 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=13070 5680 1 0 $X=12880 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=13070 5680 0 0 $X=12880 $Y=5440
X3 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=13070 11120 1 0 $X=12880 $Y=8160
X4 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 240 0 0 $X=0 $Y=0
X5 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 5680 1 0 $X=0 $Y=2720
X6 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 5680 0 0 $X=0 $Y=5440
X7 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 11120 1 0 $X=0 $Y=8160
X8 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=5710 240 0 0 $X=5520 $Y=0
X9 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=5710 5680 1 0 $X=5520 $Y=2720
X10 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=5710 5680 0 0 $X=5520 $Y=5440
X11 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=5710 11120 1 0 $X=5520 $Y=8160
X12 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=11230 240 0 0 $X=11040 $Y=0
X13 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=11230 5680 1 0 $X=11040 $Y=2720
X14 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=11230 5680 0 0 $X=11040 $Y=5440
X15 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=11230 11120 1 0 $X=11040 $Y=8160
.ends MASCO__B63

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B64                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B64 1 2
** N=2 EP=2 FDC=24
X0 1 2 MASCO__B35 $T=5980 0 0 0 $X=5980 $Y=0
X1 1 2 MASCO__B35 $T=5980 5440 0 0 $X=5980 $Y=5440
X2 1 2 MASCO__B37 $T=0 0 0 0 $X=0 $Y=0
X3 1 2 MASCO__B37 $T=0 5440 0 0 $X=0 $Y=5440
.ends MASCO__B64

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B65                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B65 1 2
** N=2 EP=2 FDC=24
X0 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=2030 2960 1 0 $X=1840 $Y=0
X1 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=2030 2960 0 0 $X=1840 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=2030 8400 1 0 $X=1840 $Y=5440
X3 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=2030 8400 0 0 $X=1840 $Y=8160
X4 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=7550 2960 1 0 $X=7360 $Y=0
X5 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=7550 2960 0 0 $X=7360 $Y=2720
X6 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=7550 8400 1 0 $X=7360 $Y=5440
X7 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=7550 8400 0 0 $X=7360 $Y=8160
X8 2 1 MASCO__B31 $T=0 0 0 0 $X=0 $Y=0
X9 2 1 MASCO__B31 $T=0 5440 0 0 $X=0 $Y=5440
.ends MASCO__B65

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B66                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B66 1 2
** N=2 EP=2 FDC=32
X0 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=13070 2960 1 0 $X=12880 $Y=0
X1 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=13070 2960 0 0 $X=12880 $Y=2720
X2 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=13070 8400 1 0 $X=12880 $Y=5440
X3 2 1 1 2 sky130_fd_sc_hd__decap_3 $T=13070 8400 0 0 $X=12880 $Y=8160
X4 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 2960 1 0 $X=0 $Y=0
X5 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 2960 0 0 $X=0 $Y=2720
X6 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 8400 1 0 $X=0 $Y=5440
X7 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=190 8400 0 0 $X=0 $Y=8160
X8 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=5710 2960 1 0 $X=5520 $Y=0
X9 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=5710 2960 0 0 $X=5520 $Y=2720
X10 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=5710 8400 1 0 $X=5520 $Y=5440
X11 2 1 1 2 sky130_fd_sc_hd__decap_12 $T=5710 8400 0 0 $X=5520 $Y=8160
X12 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=11230 2960 1 0 $X=11040 $Y=0
X13 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=11230 2960 0 0 $X=11040 $Y=2720
X14 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=11230 8400 1 0 $X=11040 $Y=5440
X15 2 1 1 2 sky130_fd_sc_hd__decap_4 $T=11230 8400 0 0 $X=11040 $Y=8160
.ends MASCO__B66

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B67                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B67 1 2
** N=2 EP=2 FDC=24
X0 2 1 MASCO__B31 $T=7360 0 0 0 $X=7360 $Y=0
X1 2 1 MASCO__B31 $T=7360 5440 0 0 $X=7360 $Y=5440
X2 1 2 MASCO__B35 $T=0 0 0 0 $X=0 $Y=0
X3 1 2 MASCO__B35 $T=0 5440 0 0 $X=0 $Y=5440
.ends MASCO__B67

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: digital_ldo_top                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt digital_ldo_top 130 143 144 131 132 145 2 3 133 146
+ 134 147 122 148 135 149 136 123 45 124
+ 150 137 125 138 151 8 139 152 126 153
+ 140 10 127 154 141 128 129 155 142
** N=332 EP=39 FDC=9490
X0 1 2 3 3 2 sky130_fd_sc_hd__diode_2 $T=352240 12720 0 0 $X=352050 $Y=12480
X1 2 4 3 5 3 2 sky130_fd_sc_hd__clkbuf_1 $T=53700 50800 0 0 $X=53510 $Y=50560
X2 2 6 3 7 3 2 sky130_fd_sc_hd__clkbuf_1 $T=55080 23600 0 0 $X=54890 $Y=23360
X3 2 7 3 5 3 2 sky130_fd_sc_hd__clkbuf_1 $T=95560 23600 0 0 $X=95370 $Y=23360
X4 2 5 3 8 3 2 sky130_fd_sc_hd__clkbuf_1 $T=98320 23600 0 0 $X=98130 $Y=23360
X5 2 9 3 7 3 2 sky130_fd_sc_hd__clkbuf_1 $T=100160 23600 0 0 $X=99970 $Y=23360
X6 2 10 3 11 3 12 2 sky130_fd_sc_hd__buf_8 $T=36220 12720 1 0 $X=36030 $Y=9760
X7 2 3 13 14 15 16 17 18 19 20
+ 21 22 23 9 24 25 26 27 28 29
+ 30 31 32 33 34 35 36 1 37 38
+ 39 40 41 42 43 44 45 46 47 48
+ 49 50 51 52 53 54 55 56 57 58
+ 59 60 61 62 63 64 65 66 67 68
+ 69 70 71 72 73 74 75 76 77 78
+ 79 80 81 82 83 DigitalLDOLogic $T=105000 25000 0 0 $X=105000 $Y=25000
X8 6 2 3 84 inverter $T=20915 20215 0 0 $X=20000 $Y=20000
X9 85 2 3 37 inverter $T=80915 20215 0 0 $X=80000 $Y=20000
X10 86 2 3 87 inverter $T=80915 30215 0 0 $X=80000 $Y=30000
X11 88 89 90 91 92 93 94 95 96 97
+ 98 99 100 101 102 103 104 105 106 107
+ 108 109 110 111 112 113 114 115 116 117
+ 118 119 2 11 3 pass_transistors $T=324695 29870 0 0 $X=325000 $Y=20000
X12 120 86 85 121 2 3 rs_latch_new $T=62095 22970 0 0 $X=60000 $Y=20000
X13 3 2 122 120 11 121 4 strong_arm $T=40430 55790 0 0 $X=40000 $Y=20000
X14 94 2 3 123 124 21 3 2 sky130_fd_sc_hd__mux2_1 $T=145240 12720 0 180 $X=140910 $Y=9760
X15 97 2 3 123 125 24 3 2 sky130_fd_sc_hd__mux2_1 $T=170540 18160 0 180 $X=166210 $Y=15200
X16 96 2 3 123 126 23 3 2 sky130_fd_sc_hd__mux2_1 $T=175140 12720 1 180 $X=170810 $Y=12480
X17 98 2 3 123 127 25 3 2 sky130_fd_sc_hd__mux2_1 $T=176060 12720 0 180 $X=171730 $Y=9760
X18 100 2 3 123 128 28 3 2 sky130_fd_sc_hd__mux2_1 $T=178360 18160 1 0 $X=178170 $Y=15200
X19 99 2 3 123 129 26 3 2 sky130_fd_sc_hd__mux2_1 $T=186640 18160 0 180 $X=182310 $Y=15200
X20 102 2 3 123 130 29 3 2 sky130_fd_sc_hd__mux2_1 $T=203660 12720 1 180 $X=199330 $Y=12480
X21 101 2 3 123 131 30 3 2 sky130_fd_sc_hd__mux2_1 $T=201820 12720 1 0 $X=201630 $Y=9760
X22 104 2 3 123 132 31 3 2 sky130_fd_sc_hd__mux2_1 $T=201820 18160 1 0 $X=201630 $Y=15200
X23 106 2 3 123 133 33 3 2 sky130_fd_sc_hd__mux2_1 $T=211020 12720 1 180 $X=206690 $Y=12480
X24 108 2 3 123 134 35 3 2 sky130_fd_sc_hd__mux2_1 $T=216540 18160 1 0 $X=216350 $Y=15200
X25 110 2 3 123 135 36 3 2 sky130_fd_sc_hd__mux2_1 $T=234020 12720 0 180 $X=229690 $Y=9760
X26 103 2 3 123 136 32 3 2 sky130_fd_sc_hd__mux2_1 $T=230340 18160 1 0 $X=230150 $Y=15200
X27 112 2 3 123 137 38 3 2 sky130_fd_sc_hd__mux2_1 $T=248280 12720 1 180 $X=243950 $Y=12480
X28 105 2 3 123 138 34 3 2 sky130_fd_sc_hd__mux2_1 $T=263000 12720 0 180 $X=258670 $Y=9760
X29 114 2 3 123 139 40 3 2 sky130_fd_sc_hd__mux2_1 $T=263000 12720 1 180 $X=258670 $Y=12480
X30 116 2 3 123 140 42 3 2 sky130_fd_sc_hd__mux2_1 $T=284160 12720 1 180 $X=279830 $Y=12480
X31 117 2 3 123 141 47 3 2 sky130_fd_sc_hd__mux2_1 $T=290140 18160 1 0 $X=289950 $Y=15200
X32 107 2 3 123 142 1 3 2 sky130_fd_sc_hd__mux2_1 $T=307160 12720 0 180 $X=302830 $Y=9760
X33 118 2 3 123 143 43 3 2 sky130_fd_sc_hd__mux2_1 $T=307160 18160 0 180 $X=302830 $Y=15200
X34 109 2 3 123 144 39 3 2 sky130_fd_sc_hd__mux2_1 $T=318200 18160 0 180 $X=313870 $Y=15200
X35 111 2 3 123 145 41 3 2 sky130_fd_sc_hd__mux2_1 $T=334760 12720 0 180 $X=330430 $Y=9760
X36 115 2 3 123 146 46 3 2 sky130_fd_sc_hd__mux2_1 $T=341660 12720 1 0 $X=341470 $Y=9760
X37 113 2 3 123 147 44 3 2 sky130_fd_sc_hd__mux2_1 $T=345800 12720 1 0 $X=345610 $Y=9760
X38 119 2 3 14 148 123 3 2 sky130_fd_sc_hd__mux2_2 $T=95100 18160 0 180 $X=90770 $Y=15200
X39 91 2 3 16 149 123 3 2 sky130_fd_sc_hd__mux2_2 $T=117640 12720 1 180 $X=113310 $Y=12480
X40 89 2 3 13 150 123 3 2 sky130_fd_sc_hd__mux2_2 $T=117640 18160 0 180 $X=113310 $Y=15200
X41 93 2 3 18 151 123 3 2 sky130_fd_sc_hd__mux2_2 $T=122240 18160 0 180 $X=117910 $Y=15200
X42 88 2 3 15 152 123 3 2 sky130_fd_sc_hd__mux2_2 $T=124080 18160 1 0 $X=123890 $Y=15200
X43 90 2 3 17 153 123 3 2 sky130_fd_sc_hd__mux2_2 $T=128220 18160 1 0 $X=128030 $Y=15200
X44 92 2 3 19 154 123 3 2 sky130_fd_sc_hd__mux2_2 $T=141100 12720 1 180 $X=136770 $Y=12480
X45 95 2 3 22 155 123 3 2 sky130_fd_sc_hd__mux2_2 $T=155820 18160 0 180 $X=151490 $Y=15200
X46 156 157 2 3 sky130_fd_sc_hd__tap_1 $T=10000 12720 1 0 $X=9810 $Y=9760
X47 158 159 2 3 sky130_fd_sc_hd__tap_1 $T=10000 12720 0 0 $X=9810 $Y=12480
X48 160 161 2 3 sky130_fd_sc_hd__tap_1 $T=10000 18160 1 0 $X=9810 $Y=15200
X49 162 163 2 3 sky130_fd_sc_hd__tap_1 $T=10000 18160 0 0 $X=9810 $Y=17920
X50 164 165 2 3 sky130_fd_sc_hd__tap_1 $T=10000 23600 1 0 $X=9810 $Y=20640
X51 166 167 2 3 sky130_fd_sc_hd__tap_1 $T=10000 23600 0 0 $X=9810 $Y=23360
X52 168 169 2 3 sky130_fd_sc_hd__tap_1 $T=10000 29040 1 0 $X=9810 $Y=26080
X53 170 171 2 3 sky130_fd_sc_hd__tap_1 $T=10000 29040 0 0 $X=9810 $Y=28800
X54 172 173 2 3 sky130_fd_sc_hd__tap_1 $T=10000 34480 1 0 $X=9810 $Y=31520
X55 174 175 2 3 sky130_fd_sc_hd__tap_1 $T=10000 34480 0 0 $X=9810 $Y=34240
X56 176 177 2 3 sky130_fd_sc_hd__tap_1 $T=10000 39920 1 0 $X=9810 $Y=36960
X57 178 179 2 3 sky130_fd_sc_hd__tap_1 $T=10000 39920 0 0 $X=9810 $Y=39680
X58 180 181 2 3 sky130_fd_sc_hd__tap_1 $T=10000 45360 1 0 $X=9810 $Y=42400
X59 182 183 2 3 sky130_fd_sc_hd__tap_1 $T=10000 45360 0 0 $X=9810 $Y=45120
X60 184 185 2 3 sky130_fd_sc_hd__tap_1 $T=10000 50800 1 0 $X=9810 $Y=47840
X61 186 187 2 3 sky130_fd_sc_hd__tap_1 $T=10000 50800 0 0 $X=9810 $Y=50560
X62 188 189 2 3 sky130_fd_sc_hd__tap_1 $T=10000 56240 1 0 $X=9810 $Y=53280
X63 190 191 2 3 sky130_fd_sc_hd__tap_1 $T=10000 56240 0 0 $X=9810 $Y=56000
X64 192 193 2 3 sky130_fd_sc_hd__tap_1 $T=10000 61680 1 0 $X=9810 $Y=58720
X65 194 195 2 3 sky130_fd_sc_hd__tap_1 $T=10000 61680 0 0 $X=9810 $Y=61440
X66 196 197 2 3 sky130_fd_sc_hd__tap_1 $T=10000 67120 1 0 $X=9810 $Y=64160
X67 198 199 2 3 sky130_fd_sc_hd__tap_1 $T=10000 67120 0 0 $X=9810 $Y=66880
X68 200 201 2 3 sky130_fd_sc_hd__tap_1 $T=10000 72560 1 0 $X=9810 $Y=69600
X69 202 203 2 3 sky130_fd_sc_hd__tap_1 $T=10000 72560 0 0 $X=9810 $Y=72320
X70 204 205 2 3 sky130_fd_sc_hd__tap_1 $T=10000 78000 1 0 $X=9810 $Y=75040
X71 206 207 2 3 sky130_fd_sc_hd__tap_1 $T=10000 78000 0 0 $X=9810 $Y=77760
X72 208 209 2 3 sky130_fd_sc_hd__tap_1 $T=10000 83440 1 0 $X=9810 $Y=80480
X73 210 211 2 3 sky130_fd_sc_hd__tap_1 $T=10000 83440 0 0 $X=9810 $Y=83200
X74 212 213 2 3 sky130_fd_sc_hd__tap_1 $T=10000 88880 1 0 $X=9810 $Y=85920
X75 214 215 2 3 sky130_fd_sc_hd__tap_1 $T=10000 88880 0 0 $X=9810 $Y=88640
X76 216 217 2 3 sky130_fd_sc_hd__tap_1 $T=10000 94320 1 0 $X=9810 $Y=91360
X77 218 219 2 3 sky130_fd_sc_hd__tap_1 $T=10000 94320 0 0 $X=9810 $Y=94080
X78 220 221 2 3 sky130_fd_sc_hd__tap_1 $T=10000 99760 1 0 $X=9810 $Y=96800
X79 222 223 2 3 sky130_fd_sc_hd__tap_1 $T=10000 99760 0 0 $X=9810 $Y=99520
X80 224 225 2 3 sky130_fd_sc_hd__tap_1 $T=10000 105200 1 0 $X=9810 $Y=102240
X81 226 227 2 3 sky130_fd_sc_hd__tap_1 $T=10000 105200 0 0 $X=9810 $Y=104960
X82 228 229 2 3 sky130_fd_sc_hd__tap_1 $T=10000 110640 1 0 $X=9810 $Y=107680
X83 230 231 2 3 sky130_fd_sc_hd__tap_1 $T=10000 110640 0 0 $X=9810 $Y=110400
X84 232 233 2 3 sky130_fd_sc_hd__tap_1 $T=10000 116080 1 0 $X=9810 $Y=113120
X85 234 235 2 3 sky130_fd_sc_hd__tap_1 $T=10000 116080 0 0 $X=9810 $Y=115840
X86 236 237 2 3 sky130_fd_sc_hd__tap_1 $T=10000 121520 1 0 $X=9810 $Y=118560
X87 238 239 2 3 sky130_fd_sc_hd__tap_1 $T=10000 121520 0 0 $X=9810 $Y=121280
X88 240 241 2 3 sky130_fd_sc_hd__tap_1 $T=10000 126960 1 0 $X=9810 $Y=124000
X89 242 243 2 3 sky130_fd_sc_hd__tap_1 $T=10000 126960 0 0 $X=9810 $Y=126720
X90 244 245 2 3 sky130_fd_sc_hd__tap_1 $T=379840 12720 0 180 $X=379190 $Y=9760
X91 246 247 2 3 sky130_fd_sc_hd__tap_1 $T=379840 12720 1 180 $X=379190 $Y=12480
X92 248 249 2 3 sky130_fd_sc_hd__tap_1 $T=379840 18160 0 180 $X=379190 $Y=15200
X93 250 251 2 3 sky130_fd_sc_hd__tap_1 $T=379840 18160 1 180 $X=379190 $Y=17920
X94 252 253 2 3 sky130_fd_sc_hd__tap_1 $T=379840 23600 0 180 $X=379190 $Y=20640
X95 254 255 2 3 sky130_fd_sc_hd__tap_1 $T=379840 23600 1 180 $X=379190 $Y=23360
X96 256 257 2 3 sky130_fd_sc_hd__tap_1 $T=379840 29040 0 180 $X=379190 $Y=26080
X97 258 259 2 3 sky130_fd_sc_hd__tap_1 $T=379840 29040 1 180 $X=379190 $Y=28800
X98 260 261 2 3 sky130_fd_sc_hd__tap_1 $T=379840 34480 0 180 $X=379190 $Y=31520
X99 262 263 2 3 sky130_fd_sc_hd__tap_1 $T=379840 34480 1 180 $X=379190 $Y=34240
X100 264 265 2 3 sky130_fd_sc_hd__tap_1 $T=379840 39920 0 180 $X=379190 $Y=36960
X101 266 267 2 3 sky130_fd_sc_hd__tap_1 $T=379840 39920 1 180 $X=379190 $Y=39680
X102 268 269 2 3 sky130_fd_sc_hd__tap_1 $T=379840 45360 0 180 $X=379190 $Y=42400
X103 270 271 2 3 sky130_fd_sc_hd__tap_1 $T=379840 45360 1 180 $X=379190 $Y=45120
X104 272 273 2 3 sky130_fd_sc_hd__tap_1 $T=379840 50800 0 180 $X=379190 $Y=47840
X105 274 275 2 3 sky130_fd_sc_hd__tap_1 $T=379840 50800 1 180 $X=379190 $Y=50560
X106 276 277 2 3 sky130_fd_sc_hd__tap_1 $T=379840 56240 0 180 $X=379190 $Y=53280
X107 278 279 2 3 sky130_fd_sc_hd__tap_1 $T=379840 56240 1 180 $X=379190 $Y=56000
X108 280 281 2 3 sky130_fd_sc_hd__tap_1 $T=379840 61680 0 180 $X=379190 $Y=58720
X109 282 283 2 3 sky130_fd_sc_hd__tap_1 $T=379840 61680 1 180 $X=379190 $Y=61440
X110 284 285 2 3 sky130_fd_sc_hd__tap_1 $T=379840 67120 0 180 $X=379190 $Y=64160
X111 286 287 2 3 sky130_fd_sc_hd__tap_1 $T=379840 67120 1 180 $X=379190 $Y=66880
X112 288 289 2 3 sky130_fd_sc_hd__tap_1 $T=379840 72560 0 180 $X=379190 $Y=69600
X113 290 291 2 3 sky130_fd_sc_hd__tap_1 $T=379840 72560 1 180 $X=379190 $Y=72320
X114 292 293 2 3 sky130_fd_sc_hd__tap_1 $T=379840 78000 0 180 $X=379190 $Y=75040
X115 294 295 2 3 sky130_fd_sc_hd__tap_1 $T=379840 78000 1 180 $X=379190 $Y=77760
X116 296 297 2 3 sky130_fd_sc_hd__tap_1 $T=379840 83440 0 180 $X=379190 $Y=80480
X117 298 299 2 3 sky130_fd_sc_hd__tap_1 $T=379840 83440 1 180 $X=379190 $Y=83200
X118 300 301 2 3 sky130_fd_sc_hd__tap_1 $T=379840 88880 0 180 $X=379190 $Y=85920
X119 302 303 2 3 sky130_fd_sc_hd__tap_1 $T=379840 88880 1 180 $X=379190 $Y=88640
X120 304 305 2 3 sky130_fd_sc_hd__tap_1 $T=379840 94320 0 180 $X=379190 $Y=91360
X121 306 307 2 3 sky130_fd_sc_hd__tap_1 $T=379840 94320 1 180 $X=379190 $Y=94080
X122 308 309 2 3 sky130_fd_sc_hd__tap_1 $T=379840 99760 0 180 $X=379190 $Y=96800
X123 310 311 2 3 sky130_fd_sc_hd__tap_1 $T=379840 99760 1 180 $X=379190 $Y=99520
X124 312 313 2 3 sky130_fd_sc_hd__tap_1 $T=379840 105200 0 180 $X=379190 $Y=102240
X125 314 315 2 3 sky130_fd_sc_hd__tap_1 $T=379840 105200 1 180 $X=379190 $Y=104960
X126 316 317 2 3 sky130_fd_sc_hd__tap_1 $T=379840 110640 0 180 $X=379190 $Y=107680
X127 318 319 2 3 sky130_fd_sc_hd__tap_1 $T=379840 110640 1 180 $X=379190 $Y=110400
X128 320 321 2 3 sky130_fd_sc_hd__tap_1 $T=379840 116080 0 180 $X=379190 $Y=113120
X129 322 323 2 3 sky130_fd_sc_hd__tap_1 $T=379840 116080 1 180 $X=379190 $Y=115840
X130 324 325 2 3 sky130_fd_sc_hd__tap_1 $T=379840 121520 0 180 $X=379190 $Y=118560
X131 326 327 2 3 sky130_fd_sc_hd__tap_1 $T=379840 121520 1 180 $X=379190 $Y=121280
X132 328 329 2 3 sky130_fd_sc_hd__tap_1 $T=379840 126960 0 180 $X=379190 $Y=124000
X133 330 331 2 3 sky130_fd_sc_hd__tap_1 $T=379840 126960 1 180 $X=379190 $Y=126720
X134 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=29320 12720 1 0 $X=29130 $Y=9760
X135 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=29320 126960 0 0 $X=29130 $Y=126720
X136 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=30700 12720 0 0 $X=30510 $Y=12480
X137 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=30700 18160 1 0 $X=30510 $Y=15200
X138 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=30700 18160 0 0 $X=30510 $Y=17920
X139 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=30700 23600 1 0 $X=30510 $Y=20640
X140 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=30700 23600 0 0 $X=30510 $Y=23360
X141 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=30700 29040 1 0 $X=30510 $Y=26080
X142 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=30700 29040 0 0 $X=30510 $Y=28800
X143 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=30700 34480 1 0 $X=30510 $Y=31520
X144 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=36680 61680 0 0 $X=36490 $Y=61440
X145 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=44040 12720 1 0 $X=43850 $Y=9760
X146 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 34480 0 0 $X=53050 $Y=34240
X147 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 39920 1 0 $X=53050 $Y=36960
X148 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 39920 0 0 $X=53050 $Y=39680
X149 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 45360 1 0 $X=53050 $Y=42400
X150 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 45360 0 0 $X=53050 $Y=45120
X151 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 50800 1 0 $X=53050 $Y=47840
X152 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 50800 0 0 $X=53050 $Y=50560
X153 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 56240 1 0 $X=53050 $Y=53280
X154 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 56240 0 0 $X=53050 $Y=56000
X155 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 61680 1 0 $X=53050 $Y=58720
X156 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=53240 61680 0 0 $X=53050 $Y=61440
X157 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=56460 12720 0 0 $X=56270 $Y=12480
X158 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=56460 18160 1 0 $X=56270 $Y=15200
X159 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=56460 18160 0 0 $X=56270 $Y=17920
X160 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=56460 23600 1 0 $X=56270 $Y=20640
X161 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=56460 23600 0 0 $X=56270 $Y=23360
X162 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=56460 29040 1 0 $X=56270 $Y=26080
X163 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=56460 29040 0 0 $X=56270 $Y=28800
X164 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=56460 34480 1 0 $X=56270 $Y=31520
X165 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=58760 12720 1 0 $X=58570 $Y=9760
X166 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=63360 50800 0 0 $X=63170 $Y=50560
X167 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=63360 61680 1 0 $X=63170 $Y=58720
X168 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=63360 61680 0 0 $X=63170 $Y=61440
X169 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 12720 1 0 $X=73290 $Y=9760
X170 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=73480 61680 0 0 $X=73290 $Y=61440
X171 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 12720 1 0 $X=88010 $Y=9760
X172 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=88200 61680 0 0 $X=88010 $Y=61440
X173 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 12720 0 0 $X=90310 $Y=12480
X174 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 18160 1 0 $X=90310 $Y=15200
X175 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 18160 0 0 $X=90310 $Y=17920
X176 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 23600 1 0 $X=90310 $Y=20640
X177 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 23600 0 0 $X=90310 $Y=23360
X178 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 29040 1 0 $X=90310 $Y=26080
X179 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 29040 0 0 $X=90310 $Y=28800
X180 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 34480 1 0 $X=90310 $Y=31520
X181 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 34480 0 0 $X=90310 $Y=34240
X182 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 39920 1 0 $X=90310 $Y=36960
X183 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 39920 0 0 $X=90310 $Y=39680
X184 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=90500 45360 1 0 $X=90310 $Y=42400
X185 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 23600 0 0 $X=101350 $Y=23360
X186 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 45360 1 0 $X=101350 $Y=42400
X187 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 45360 0 0 $X=101350 $Y=45120
X188 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 50800 1 0 $X=101350 $Y=47840
X189 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 50800 0 0 $X=101350 $Y=50560
X190 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 56240 1 0 $X=101350 $Y=53280
X191 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 56240 0 0 $X=101350 $Y=56000
X192 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 61680 1 0 $X=101350 $Y=58720
X193 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 61680 0 0 $X=101350 $Y=61440
X194 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 67120 1 0 $X=101350 $Y=64160
X195 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 67120 0 0 $X=101350 $Y=66880
X196 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 72560 1 0 $X=101350 $Y=69600
X197 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 72560 0 0 $X=101350 $Y=72320
X198 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 78000 1 0 $X=101350 $Y=75040
X199 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 78000 0 0 $X=101350 $Y=77760
X200 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 83440 1 0 $X=101350 $Y=80480
X201 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 83440 0 0 $X=101350 $Y=83200
X202 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 88880 1 0 $X=101350 $Y=85920
X203 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=101540 88880 0 0 $X=101350 $Y=88640
X204 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=102920 18160 1 0 $X=102730 $Y=15200
X205 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 12720 1 0 $X=117450 $Y=9760
X206 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 12720 0 0 $X=117450 $Y=12480
X207 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=117640 18160 1 0 $X=117450 $Y=15200
X208 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 12720 1 0 $X=132170 $Y=9760
X209 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 12720 0 0 $X=132170 $Y=12480
X210 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=132360 18160 1 0 $X=132170 $Y=15200
X211 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=147080 12720 1 0 $X=146890 $Y=9760
X212 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=161800 18160 1 0 $X=161610 $Y=15200
X213 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=176520 18160 1 0 $X=176330 $Y=15200
X214 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=191240 18160 1 0 $X=191050 $Y=15200
X215 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=205960 12720 1 0 $X=205770 $Y=9760
X216 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=205960 12720 0 0 $X=205770 $Y=12480
X217 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=205960 18160 1 0 $X=205770 $Y=15200
X218 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=220680 12720 1 0 $X=220490 $Y=9760
X219 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=220680 12720 0 0 $X=220490 $Y=12480
X220 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=220680 18160 1 0 $X=220490 $Y=15200
X221 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=235400 18160 1 0 $X=235210 $Y=15200
X222 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=250120 18160 1 0 $X=249930 $Y=15200
X223 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=264840 12720 1 0 $X=264650 $Y=9760
X224 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=264840 12720 0 0 $X=264650 $Y=12480
X225 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=264840 18160 1 0 $X=264650 $Y=15200
X226 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=279560 12720 1 0 $X=279370 $Y=9760
X227 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=279560 12720 0 0 $X=279370 $Y=12480
X228 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=279560 18160 1 0 $X=279370 $Y=15200
X229 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=294280 12720 1 0 $X=294090 $Y=9760
X230 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=294280 12720 0 0 $X=294090 $Y=12480
X231 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=294280 18160 1 0 $X=294090 $Y=15200
X232 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=309000 18160 1 0 $X=308810 $Y=15200
X233 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=309000 18160 0 0 $X=308810 $Y=17920
X234 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=309000 88880 1 0 $X=308810 $Y=85920
X235 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=309000 88880 0 0 $X=308810 $Y=88640
X236 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=321880 12720 0 0 $X=321690 $Y=12480
X237 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=321880 18160 1 0 $X=321690 $Y=15200
X238 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=321880 18160 0 0 $X=321690 $Y=17920
X239 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=321880 50800 1 0 $X=321690 $Y=47840
X240 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=323720 12720 1 0 $X=323530 $Y=9760
X241 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=323720 126960 0 0 $X=323530 $Y=126720
X242 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=338440 12720 1 0 $X=338250 $Y=9760
X243 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=338440 126960 0 0 $X=338250 $Y=126720
X244 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 12720 1 0 $X=352970 $Y=9760
X245 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 12720 0 0 $X=352970 $Y=12480
X246 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 18160 1 0 $X=352970 $Y=15200
X247 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 18160 0 0 $X=352970 $Y=17920
X248 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 23600 1 0 $X=352970 $Y=20640
X249 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 23600 0 0 $X=352970 $Y=23360
X250 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 29040 1 0 $X=352970 $Y=26080
X251 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 29040 0 0 $X=352970 $Y=28800
X252 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 34480 1 0 $X=352970 $Y=31520
X253 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 34480 0 0 $X=352970 $Y=34240
X254 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 39920 1 0 $X=352970 $Y=36960
X255 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 39920 0 0 $X=352970 $Y=39680
X256 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 45360 1 0 $X=352970 $Y=42400
X257 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=353160 45360 0 0 $X=352970 $Y=45120
X258 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=367880 12720 1 0 $X=367690 $Y=9760
X259 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=367880 45360 0 0 $X=367690 $Y=45120
X260 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 12720 1 0 $X=378730 $Y=9760
X261 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 12720 0 0 $X=378730 $Y=12480
X262 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 18160 1 0 $X=378730 $Y=15200
X263 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 18160 0 0 $X=378730 $Y=17920
X264 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 23600 1 0 $X=378730 $Y=20640
X265 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 23600 0 0 $X=378730 $Y=23360
X266 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 29040 1 0 $X=378730 $Y=26080
X267 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 29040 0 0 $X=378730 $Y=28800
X268 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 34480 1 0 $X=378730 $Y=31520
X269 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 34480 0 0 $X=378730 $Y=34240
X270 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 39920 1 0 $X=378730 $Y=36960
X271 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 39920 0 0 $X=378730 $Y=39680
X272 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 45360 1 0 $X=378730 $Y=42400
X273 2 3 sky130_fd_sc_hd__tapvpwrvgnd_1 $T=378920 45360 0 0 $X=378730 $Y=45120
X274 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 12720 1 0 $X=10270 $Y=9760
X275 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 12720 0 0 $X=10270 $Y=12480
X276 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 18160 1 0 $X=10270 $Y=15200
X277 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 18160 0 0 $X=10270 $Y=17920
X278 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 23600 1 0 $X=10270 $Y=20640
X279 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 23600 0 0 $X=10270 $Y=23360
X280 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 29040 1 0 $X=10270 $Y=26080
X281 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 29040 0 0 $X=10270 $Y=28800
X282 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 34480 1 0 $X=10270 $Y=31520
X283 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 34480 0 0 $X=10270 $Y=34240
X284 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 39920 1 0 $X=10270 $Y=36960
X285 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 39920 0 0 $X=10270 $Y=39680
X286 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 45360 1 0 $X=10270 $Y=42400
X287 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 45360 0 0 $X=10270 $Y=45120
X288 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 50800 1 0 $X=10270 $Y=47840
X289 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 50800 0 0 $X=10270 $Y=50560
X290 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 56240 1 0 $X=10270 $Y=53280
X291 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 56240 0 0 $X=10270 $Y=56000
X292 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 61680 1 0 $X=10270 $Y=58720
X293 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 61680 0 0 $X=10270 $Y=61440
X294 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 67120 1 0 $X=10270 $Y=64160
X295 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 67120 0 0 $X=10270 $Y=66880
X296 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 72560 1 0 $X=10270 $Y=69600
X297 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 72560 0 0 $X=10270 $Y=72320
X298 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 78000 1 0 $X=10270 $Y=75040
X299 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 78000 0 0 $X=10270 $Y=77760
X300 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 83440 1 0 $X=10270 $Y=80480
X301 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 83440 0 0 $X=10270 $Y=83200
X302 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 88880 1 0 $X=10270 $Y=85920
X303 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 88880 0 0 $X=10270 $Y=88640
X304 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 94320 1 0 $X=10270 $Y=91360
X305 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 94320 0 0 $X=10270 $Y=94080
X306 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 99760 1 0 $X=10270 $Y=96800
X307 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 99760 0 0 $X=10270 $Y=99520
X308 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 105200 1 0 $X=10270 $Y=102240
X309 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 105200 0 0 $X=10270 $Y=104960
X310 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 110640 1 0 $X=10270 $Y=107680
X311 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 110640 0 0 $X=10270 $Y=110400
X312 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 116080 1 0 $X=10270 $Y=113120
X313 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 116080 0 0 $X=10270 $Y=115840
X314 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 121520 1 0 $X=10270 $Y=118560
X315 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 121520 0 0 $X=10270 $Y=121280
X316 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 126960 1 0 $X=10270 $Y=124000
X317 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=10460 126960 0 0 $X=10270 $Y=126720
X318 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=27940 12720 0 0 $X=27750 $Y=12480
X319 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=27940 34480 1 0 $X=27750 $Y=31520
X320 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=33460 12720 1 0 $X=33270 $Y=9760
X321 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=53700 18160 1 0 $X=53510 $Y=15200
X322 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=53700 18160 0 0 $X=53510 $Y=17920
X323 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=53700 23600 1 0 $X=53510 $Y=20640
X324 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=53700 29040 1 0 $X=53510 $Y=26080
X325 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=53700 29040 0 0 $X=53510 $Y=28800
X326 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=53700 34480 1 0 $X=53510 $Y=31520
X327 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 34480 0 0 $X=59030 $Y=34240
X328 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 39920 1 0 $X=59030 $Y=36960
X329 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 39920 0 0 $X=59030 $Y=39680
X330 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 45360 1 0 $X=59030 $Y=42400
X331 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 45360 0 0 $X=59030 $Y=45120
X332 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 50800 1 0 $X=59030 $Y=47840
X333 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 56240 1 0 $X=59030 $Y=53280
X334 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 56240 0 0 $X=59030 $Y=56000
X335 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 61680 1 0 $X=59030 $Y=58720
X336 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=59220 61680 0 0 $X=59030 $Y=61440
X337 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=60600 50800 0 0 $X=60410 $Y=50560
X338 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 34480 0 0 $X=69150 $Y=34240
X339 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 39920 1 0 $X=69150 $Y=36960
X340 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 39920 0 0 $X=69150 $Y=39680
X341 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 45360 1 0 $X=69150 $Y=42400
X342 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 45360 0 0 $X=69150 $Y=45120
X343 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 50800 1 0 $X=69150 $Y=47840
X344 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 50800 0 0 $X=69150 $Y=50560
X345 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 56240 1 0 $X=69150 $Y=53280
X346 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 56240 0 0 $X=69150 $Y=56000
X347 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 61680 1 0 $X=69150 $Y=58720
X348 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=69340 61680 0 0 $X=69150 $Y=61440
X349 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=73480 34480 1 0 $X=73290 $Y=31520
X350 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=73940 45360 1 0 $X=73750 $Y=42400
X351 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=84520 12720 0 0 $X=84330 $Y=12480
X352 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=87740 45360 1 0 $X=87550 $Y=42400
X353 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=90960 23600 0 0 $X=90770 $Y=23360
X354 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=98780 18160 1 0 $X=98590 $Y=15200
X355 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=100160 12720 0 0 $X=99970 $Y=12480
X356 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=108900 12720 0 0 $X=108710 $Y=12480
X357 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=108900 18160 1 0 $X=108710 $Y=15200
X358 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=132820 12720 0 0 $X=132630 $Y=12480
X359 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=138340 12720 1 0 $X=138150 $Y=9760
X360 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=141100 12720 0 0 $X=140910 $Y=12480
X361 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=147540 18160 1 0 $X=147350 $Y=15200
X362 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=155820 18160 1 0 $X=155630 $Y=15200
X363 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=162260 18160 1 0 $X=162070 $Y=15200
X364 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=167780 12720 1 0 $X=167590 $Y=9760
X365 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=170540 18160 1 0 $X=170350 $Y=15200
X366 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=186640 18160 1 0 $X=186450 $Y=15200
X367 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=195380 12720 0 0 $X=195190 $Y=12480
X368 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=197220 12720 1 0 $X=197030 $Y=9760
X369 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=197220 18160 1 0 $X=197030 $Y=15200
X370 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=211940 18160 1 0 $X=211750 $Y=15200
X371 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=216540 12720 0 0 $X=216350 $Y=12480
X372 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=241380 12720 0 0 $X=241190 $Y=12480
X373 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=256100 12720 1 0 $X=255910 $Y=9760
X374 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=256100 12720 0 0 $X=255910 $Y=12480
X375 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=285540 18160 1 0 $X=285350 $Y=15200
X376 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=289680 12720 0 0 $X=289490 $Y=12480
X377 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=300260 12720 1 0 $X=300070 $Y=9760
X378 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=300260 18160 1 0 $X=300070 $Y=15200
X379 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=306240 18160 0 0 $X=306050 $Y=17920
X380 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=306240 88880 0 0 $X=306050 $Y=88640
X381 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=309460 18160 1 0 $X=309270 $Y=15200
X382 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=327860 12720 1 0 $X=327670 $Y=9760
X383 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=338900 12720 1 0 $X=338710 $Y=9760
X384 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=348100 12720 0 0 $X=347910 $Y=12480
X385 2 3 3 2 sky130_fd_sc_hd__decap_6 $T=348100 50800 1 0 $X=347910 $Y=47840
X386 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=15060 18160 1 0 $X=14870 $Y=15200
X387 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=15060 18160 0 0 $X=14870 $Y=17920
X388 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=15060 23600 1 0 $X=14870 $Y=20640
X389 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=15060 23600 0 0 $X=14870 $Y=23360
X390 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=15060 29040 1 0 $X=14870 $Y=26080
X391 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=15060 29040 0 0 $X=14870 $Y=28800
X392 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=27940 12720 1 0 $X=27750 $Y=9760
X393 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=27940 121520 0 0 $X=27750 $Y=121280
X394 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=27940 126960 1 0 $X=27750 $Y=124000
X395 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=27940 126960 0 0 $X=27750 $Y=126720
X396 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=34840 18160 1 0 $X=34650 $Y=15200
X397 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=34840 18160 0 0 $X=34650 $Y=17920
X398 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=34840 23600 1 0 $X=34650 $Y=20640
X399 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=34840 23600 0 0 $X=34650 $Y=23360
X400 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=34840 29040 1 0 $X=34650 $Y=26080
X401 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=34840 29040 0 0 $X=34650 $Y=28800
X402 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=34840 34480 1 0 $X=34650 $Y=31520
X403 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=35300 61680 0 0 $X=35110 $Y=61440
X404 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=36220 18160 1 0 $X=36030 $Y=15200
X405 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=36220 18160 0 0 $X=36030 $Y=17920
X406 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=36220 23600 1 0 $X=36030 $Y=20640
X407 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=36220 23600 0 0 $X=36030 $Y=23360
X408 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=36220 29040 1 0 $X=36030 $Y=26080
X409 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=36220 29040 0 0 $X=36030 $Y=28800
X410 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=36220 34480 1 0 $X=36030 $Y=31520
X411 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=41740 12720 1 0 $X=41550 $Y=9760
X412 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=51860 61680 0 0 $X=51670 $Y=61440
X413 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=53700 23600 0 0 $X=53510 $Y=23360
X414 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=55080 12720 0 0 $X=54890 $Y=12480
X415 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=57380 12720 1 0 $X=57190 $Y=9760
X416 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=61980 61680 1 0 $X=61790 $Y=58720
X417 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=61980 61680 0 0 $X=61790 $Y=61440
X418 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=72100 12720 1 0 $X=71910 $Y=9760
X419 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=72100 61680 0 0 $X=71910 $Y=61440
X420 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=76240 34480 1 0 $X=76050 $Y=31520
X421 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 12720 1 0 $X=86630 $Y=9760
X422 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 56240 0 0 $X=86630 $Y=56000
X423 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 61680 1 0 $X=86630 $Y=58720
X424 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 61680 0 0 $X=86630 $Y=61440
X425 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 67120 1 0 $X=86630 $Y=64160
X426 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 67120 0 0 $X=86630 $Y=66880
X427 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 72560 1 0 $X=86630 $Y=69600
X428 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 72560 0 0 $X=86630 $Y=72320
X429 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 78000 1 0 $X=86630 $Y=75040
X430 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 78000 0 0 $X=86630 $Y=77760
X431 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 83440 1 0 $X=86630 $Y=80480
X432 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 83440 0 0 $X=86630 $Y=83200
X433 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 88880 1 0 $X=86630 $Y=85920
X434 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 88880 0 0 $X=86630 $Y=88640
X435 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 94320 1 0 $X=86630 $Y=91360
X436 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 94320 0 0 $X=86630 $Y=94080
X437 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 99760 1 0 $X=86630 $Y=96800
X438 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 99760 0 0 $X=86630 $Y=99520
X439 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 105200 1 0 $X=86630 $Y=102240
X440 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 105200 0 0 $X=86630 $Y=104960
X441 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 110640 1 0 $X=86630 $Y=107680
X442 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 110640 0 0 $X=86630 $Y=110400
X443 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 116080 1 0 $X=86630 $Y=113120
X444 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 116080 0 0 $X=86630 $Y=115840
X445 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 121520 1 0 $X=86630 $Y=118560
X446 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 121520 0 0 $X=86630 $Y=121280
X447 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 126960 1 0 $X=86630 $Y=124000
X448 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=86820 126960 0 0 $X=86630 $Y=126720
X449 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=89120 12720 0 0 $X=88930 $Y=12480
X450 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=96940 23600 0 0 $X=96750 $Y=23360
X451 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=100160 45360 1 0 $X=99970 $Y=42400
X452 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=101540 12720 1 0 $X=101350 $Y=9760
X453 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=101540 18160 1 0 $X=101350 $Y=15200
X454 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=116260 12720 1 0 $X=116070 $Y=9760
X455 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=116260 126960 1 0 $X=116070 $Y=124000
X456 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=116260 126960 0 0 $X=116070 $Y=126720
X457 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=130980 12720 1 0 $X=130790 $Y=9760
X458 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=130980 12720 0 0 $X=130790 $Y=12480
X459 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=135580 12720 0 0 $X=135390 $Y=12480
X460 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 94320 1 0 $X=145510 $Y=91360
X461 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 94320 0 0 $X=145510 $Y=94080
X462 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 99760 1 0 $X=145510 $Y=96800
X463 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 99760 0 0 $X=145510 $Y=99520
X464 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 105200 1 0 $X=145510 $Y=102240
X465 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 105200 0 0 $X=145510 $Y=104960
X466 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 110640 1 0 $X=145510 $Y=107680
X467 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 110640 0 0 $X=145510 $Y=110400
X468 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 116080 1 0 $X=145510 $Y=113120
X469 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 116080 0 0 $X=145510 $Y=115840
X470 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 121520 1 0 $X=145510 $Y=118560
X471 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 121520 0 0 $X=145510 $Y=121280
X472 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 126960 1 0 $X=145510 $Y=124000
X473 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=145700 126960 0 0 $X=145510 $Y=126720
X474 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=150300 18160 1 0 $X=150110 $Y=15200
X475 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=160420 12720 1 0 $X=160230 $Y=9760
X476 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=160420 12720 0 0 $X=160230 $Y=12480
X477 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=160420 18160 1 0 $X=160230 $Y=15200
X478 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=165020 18160 1 0 $X=164830 $Y=15200
X479 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=169620 12720 0 0 $X=169430 $Y=12480
X480 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=170540 12720 1 0 $X=170350 $Y=9760
X481 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=175140 12720 0 0 $X=174950 $Y=12480
X482 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=175140 18160 1 0 $X=174950 $Y=15200
X483 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=175140 126960 1 0 $X=174950 $Y=124000
X484 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=175140 126960 0 0 $X=174950 $Y=126720
X485 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=176980 18160 1 0 $X=176790 $Y=15200
X486 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=198140 12720 0 0 $X=197950 $Y=12480
X487 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=203660 12720 0 0 $X=203470 $Y=12480
X488 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 94320 1 0 $X=204390 $Y=91360
X489 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 94320 0 0 $X=204390 $Y=94080
X490 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 99760 1 0 $X=204390 $Y=96800
X491 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 99760 0 0 $X=204390 $Y=99520
X492 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 105200 1 0 $X=204390 $Y=102240
X493 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 105200 0 0 $X=204390 $Y=104960
X494 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 110640 1 0 $X=204390 $Y=107680
X495 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 110640 0 0 $X=204390 $Y=110400
X496 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 116080 1 0 $X=204390 $Y=113120
X497 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 116080 0 0 $X=204390 $Y=115840
X498 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 121520 1 0 $X=204390 $Y=118560
X499 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 121520 0 0 $X=204390 $Y=121280
X500 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 126960 1 0 $X=204390 $Y=124000
X501 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=204580 126960 0 0 $X=204390 $Y=126720
X502 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=219300 12720 1 0 $X=219110 $Y=9760
X503 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=219300 12720 0 0 $X=219110 $Y=12480
X504 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=228500 12720 1 0 $X=228310 $Y=9760
X505 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=234020 126960 1 0 $X=233830 $Y=124000
X506 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=234020 126960 0 0 $X=233830 $Y=126720
X507 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=248740 12720 1 0 $X=248550 $Y=9760
X508 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=248740 18160 1 0 $X=248550 $Y=15200
X509 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 18160 1 0 $X=263270 $Y=15200
X510 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 94320 1 0 $X=263270 $Y=91360
X511 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 94320 0 0 $X=263270 $Y=94080
X512 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 99760 1 0 $X=263270 $Y=96800
X513 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 99760 0 0 $X=263270 $Y=99520
X514 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 105200 1 0 $X=263270 $Y=102240
X515 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 105200 0 0 $X=263270 $Y=104960
X516 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 110640 1 0 $X=263270 $Y=107680
X517 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 110640 0 0 $X=263270 $Y=110400
X518 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 116080 1 0 $X=263270 $Y=113120
X519 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 116080 0 0 $X=263270 $Y=115840
X520 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 121520 1 0 $X=263270 $Y=118560
X521 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 121520 0 0 $X=263270 $Y=121280
X522 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 126960 1 0 $X=263270 $Y=124000
X523 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=263460 126960 0 0 $X=263270 $Y=126720
X524 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=278180 12720 1 0 $X=277990 $Y=9760
X525 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=278180 12720 0 0 $X=277990 $Y=12480
X526 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=278180 18160 1 0 $X=277990 $Y=15200
X527 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=292900 12720 1 0 $X=292710 $Y=9760
X528 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=292900 126960 1 0 $X=292710 $Y=124000
X529 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=292900 126960 0 0 $X=292710 $Y=126720
X530 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=307620 12720 0 0 $X=307430 $Y=12480
X531 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=307620 88880 1 0 $X=307430 $Y=85920
X532 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=320500 12720 0 0 $X=320310 $Y=12480
X533 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=320500 18160 0 0 $X=320310 $Y=17920
X534 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=320500 50800 1 0 $X=320310 $Y=47840
X535 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 12720 1 0 $X=322150 $Y=9760
X536 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 50800 0 0 $X=322150 $Y=50560
X537 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 56240 1 0 $X=322150 $Y=53280
X538 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 56240 0 0 $X=322150 $Y=56000
X539 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 61680 1 0 $X=322150 $Y=58720
X540 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 61680 0 0 $X=322150 $Y=61440
X541 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 67120 1 0 $X=322150 $Y=64160
X542 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 67120 0 0 $X=322150 $Y=66880
X543 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 72560 1 0 $X=322150 $Y=69600
X544 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 72560 0 0 $X=322150 $Y=72320
X545 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 78000 1 0 $X=322150 $Y=75040
X546 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 78000 0 0 $X=322150 $Y=77760
X547 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 83440 1 0 $X=322150 $Y=80480
X548 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 83440 0 0 $X=322150 $Y=83200
X549 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 88880 1 0 $X=322150 $Y=85920
X550 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 88880 0 0 $X=322150 $Y=88640
X551 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 94320 1 0 $X=322150 $Y=91360
X552 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 94320 0 0 $X=322150 $Y=94080
X553 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 99760 1 0 $X=322150 $Y=96800
X554 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 99760 0 0 $X=322150 $Y=99520
X555 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 105200 1 0 $X=322150 $Y=102240
X556 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 105200 0 0 $X=322150 $Y=104960
X557 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 110640 1 0 $X=322150 $Y=107680
X558 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 110640 0 0 $X=322150 $Y=110400
X559 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 116080 1 0 $X=322150 $Y=113120
X560 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 116080 0 0 $X=322150 $Y=115840
X561 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 121520 1 0 $X=322150 $Y=118560
X562 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 121520 0 0 $X=322150 $Y=121280
X563 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 126960 1 0 $X=322150 $Y=124000
X564 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=322340 126960 0 0 $X=322150 $Y=126720
X565 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=337060 126960 0 0 $X=336870 $Y=126720
X566 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=350860 12720 0 0 $X=350670 $Y=12480
X567 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=350860 50800 1 0 $X=350670 $Y=47840
X568 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=351780 12720 1 0 $X=351590 $Y=9760
X569 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=351780 126960 0 0 $X=351590 $Y=126720
X570 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=366500 12720 1 0 $X=366310 $Y=9760
X571 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=366500 45360 0 0 $X=366310 $Y=45120
X572 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 12720 1 0 $X=377350 $Y=9760
X573 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 12720 0 0 $X=377350 $Y=12480
X574 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 18160 1 0 $X=377350 $Y=15200
X575 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 18160 0 0 $X=377350 $Y=17920
X576 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 23600 1 0 $X=377350 $Y=20640
X577 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 23600 0 0 $X=377350 $Y=23360
X578 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 29040 1 0 $X=377350 $Y=26080
X579 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 29040 0 0 $X=377350 $Y=28800
X580 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 34480 1 0 $X=377350 $Y=31520
X581 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 34480 0 0 $X=377350 $Y=34240
X582 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 39920 1 0 $X=377350 $Y=36960
X583 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 39920 0 0 $X=377350 $Y=39680
X584 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 45360 1 0 $X=377350 $Y=42400
X585 2 3 3 2 sky130_fd_sc_hd__decap_3 $T=377540 45360 0 0 $X=377350 $Y=45120
X586 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=15060 12720 1 0 $X=14870 $Y=9760
X587 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=15060 121520 0 0 $X=14870 $Y=121280
X588 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=15060 126960 1 0 $X=14870 $Y=124000
X589 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=15060 126960 0 0 $X=14870 $Y=126720
X590 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=16900 12720 0 0 $X=16710 $Y=12480
X591 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=16900 34480 1 0 $X=16710 $Y=31520
X592 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=20580 12720 1 0 $X=20390 $Y=9760
X593 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=20580 121520 0 0 $X=20390 $Y=121280
X594 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=20580 126960 1 0 $X=20390 $Y=124000
X595 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=20580 126960 0 0 $X=20390 $Y=126720
X596 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=22420 12720 0 0 $X=22230 $Y=12480
X597 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=22420 34480 1 0 $X=22230 $Y=31520
X598 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=29780 126960 0 0 $X=29590 $Y=126720
X599 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=31160 12720 0 0 $X=30970 $Y=12480
X600 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=36680 12720 0 0 $X=36490 $Y=12480
X601 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=37140 61680 0 0 $X=36950 $Y=61440
X602 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=42200 12720 0 0 $X=42010 $Y=12480
X603 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=42660 61680 0 0 $X=42470 $Y=61440
X604 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=44500 12720 1 0 $X=44310 $Y=9760
X605 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=47720 12720 0 0 $X=47530 $Y=12480
X606 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=50020 12720 1 0 $X=49830 $Y=9760
X607 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 34480 0 0 $X=53510 $Y=34240
X608 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 39920 1 0 $X=53510 $Y=36960
X609 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 39920 0 0 $X=53510 $Y=39680
X610 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 45360 1 0 $X=53510 $Y=42400
X611 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 45360 0 0 $X=53510 $Y=45120
X612 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 50800 1 0 $X=53510 $Y=47840
X613 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 56240 1 0 $X=53510 $Y=53280
X614 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 56240 0 0 $X=53510 $Y=56000
X615 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 61680 1 0 $X=53510 $Y=58720
X616 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=53700 61680 0 0 $X=53510 $Y=61440
X617 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=55080 50800 0 0 $X=54890 $Y=50560
X618 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=56920 12720 0 0 $X=56730 $Y=12480
X619 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=56920 34480 1 0 $X=56730 $Y=31520
X620 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=59220 12720 1 0 $X=59030 $Y=9760
X621 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=62440 12720 0 0 $X=62250 $Y=12480
X622 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=62440 34480 1 0 $X=62250 $Y=31520
X623 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 34480 0 0 $X=63630 $Y=34240
X624 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 39920 1 0 $X=63630 $Y=36960
X625 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 39920 0 0 $X=63630 $Y=39680
X626 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 45360 1 0 $X=63630 $Y=42400
X627 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 45360 0 0 $X=63630 $Y=45120
X628 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 50800 1 0 $X=63630 $Y=47840
X629 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 50800 0 0 $X=63630 $Y=50560
X630 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 56240 1 0 $X=63630 $Y=53280
X631 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 56240 0 0 $X=63630 $Y=56000
X632 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 61680 1 0 $X=63630 $Y=58720
X633 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=63820 61680 0 0 $X=63630 $Y=61440
X634 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=64740 12720 1 0 $X=64550 $Y=9760
X635 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=67960 12720 0 0 $X=67770 $Y=12480
X636 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=67960 34480 1 0 $X=67770 $Y=31520
X637 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=73480 12720 0 0 $X=73290 $Y=12480
X638 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=73940 12720 1 0 $X=73750 $Y=9760
X639 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=73940 56240 0 0 $X=73750 $Y=56000
X640 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=73940 61680 1 0 $X=73750 $Y=58720
X641 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=73940 61680 0 0 $X=73750 $Y=61440
X642 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=76700 45360 1 0 $X=76510 $Y=42400
X643 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=79000 12720 0 0 $X=78810 $Y=12480
X644 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=79460 12720 1 0 $X=79270 $Y=9760
X645 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=79460 56240 0 0 $X=79270 $Y=56000
X646 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=79460 61680 1 0 $X=79270 $Y=58720
X647 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=79460 61680 0 0 $X=79270 $Y=61440
X648 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=82220 45360 1 0 $X=82030 $Y=42400
X649 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=88660 12720 1 0 $X=88470 $Y=9760
X650 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=88660 61680 0 0 $X=88470 $Y=61440
X651 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=90960 12720 0 0 $X=90770 $Y=12480
X652 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=90960 18160 0 0 $X=90770 $Y=17920
X653 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=90960 23600 1 0 $X=90770 $Y=20640
X654 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=90960 45360 1 0 $X=90770 $Y=42400
X655 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=94180 12720 1 0 $X=93990 $Y=9760
X656 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=94180 61680 0 0 $X=93990 $Y=61440
X657 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=102000 18160 0 0 $X=101810 $Y=17920
X658 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=102000 88880 0 0 $X=101810 $Y=88640
X659 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=103380 18160 1 0 $X=103190 $Y=15200
X660 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=103380 126960 1 0 $X=103190 $Y=124000
X661 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=103380 126960 0 0 $X=103190 $Y=126720
X662 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=107520 18160 0 0 $X=107330 $Y=17920
X663 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=107520 88880 0 0 $X=107330 $Y=88640
X664 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=108900 12720 1 0 $X=108710 $Y=9760
X665 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=108900 126960 1 0 $X=108710 $Y=124000
X666 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=108900 126960 0 0 $X=108710 $Y=126720
X667 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=113040 18160 0 0 $X=112850 $Y=17920
X668 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=113040 88880 0 0 $X=112850 $Y=88640
X669 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=118100 12720 1 0 $X=117910 $Y=9760
X670 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=118100 12720 0 0 $X=117910 $Y=12480
X671 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=118560 18160 0 0 $X=118370 $Y=17920
X672 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=118560 88880 0 0 $X=118370 $Y=88640
X673 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=123620 12720 1 0 $X=123430 $Y=9760
X674 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=123620 12720 0 0 $X=123430 $Y=12480
X675 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=124080 18160 0 0 $X=123890 $Y=17920
X676 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=124080 88880 0 0 $X=123890 $Y=88640
X677 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=129600 18160 0 0 $X=129410 $Y=17920
X678 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=129600 88880 0 0 $X=129410 $Y=88640
X679 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=132820 12720 1 0 $X=132630 $Y=9760
X680 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=132820 18160 1 0 $X=132630 $Y=15200
X681 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=132820 126960 1 0 $X=132630 $Y=124000
X682 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=132820 126960 0 0 $X=132630 $Y=126720
X683 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=135120 18160 0 0 $X=134930 $Y=17920
X684 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=135120 88880 0 0 $X=134930 $Y=88640
X685 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=138340 18160 1 0 $X=138150 $Y=15200
X686 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=138340 126960 1 0 $X=138150 $Y=124000
X687 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=138340 126960 0 0 $X=138150 $Y=126720
X688 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=140640 18160 0 0 $X=140450 $Y=17920
X689 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=140640 88880 0 0 $X=140450 $Y=88640
X690 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=146160 18160 0 0 $X=145970 $Y=17920
X691 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=146160 88880 0 0 $X=145970 $Y=88640
X692 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=147540 12720 1 0 $X=147350 $Y=9760
X693 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=147540 12720 0 0 $X=147350 $Y=12480
X694 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=151680 18160 0 0 $X=151490 $Y=17920
X695 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=151680 88880 0 0 $X=151490 $Y=88640
X696 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=153060 12720 1 0 $X=152870 $Y=9760
X697 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=153060 12720 0 0 $X=152870 $Y=12480
X698 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=157200 18160 0 0 $X=157010 $Y=17920
X699 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=157200 88880 0 0 $X=157010 $Y=88640
X700 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=162260 126960 1 0 $X=162070 $Y=124000
X701 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=162260 126960 0 0 $X=162070 $Y=126720
X702 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=162720 18160 0 0 $X=162530 $Y=17920
X703 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=162720 88880 0 0 $X=162530 $Y=88640
X704 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=167780 126960 1 0 $X=167590 $Y=124000
X705 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=167780 126960 0 0 $X=167590 $Y=126720
X706 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=168240 18160 0 0 $X=168050 $Y=17920
X707 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=168240 88880 0 0 $X=168050 $Y=88640
X708 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=173760 18160 0 0 $X=173570 $Y=17920
X709 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=173760 88880 0 0 $X=173570 $Y=88640
X710 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=179280 18160 0 0 $X=179090 $Y=17920
X711 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=179280 88880 0 0 $X=179090 $Y=88640
X712 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=184800 18160 0 0 $X=184610 $Y=17920
X713 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=184800 88880 0 0 $X=184610 $Y=88640
X714 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=190320 18160 0 0 $X=190130 $Y=17920
X715 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=190320 88880 0 0 $X=190130 $Y=88640
X716 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=191700 12720 1 0 $X=191510 $Y=9760
X717 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=191700 18160 1 0 $X=191510 $Y=15200
X718 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=191700 126960 1 0 $X=191510 $Y=124000
X719 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=191700 126960 0 0 $X=191510 $Y=126720
X720 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=195840 18160 0 0 $X=195650 $Y=17920
X721 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=195840 88880 0 0 $X=195650 $Y=88640
X722 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=197220 126960 1 0 $X=197030 $Y=124000
X723 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=197220 126960 0 0 $X=197030 $Y=126720
X724 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=201360 18160 0 0 $X=201170 $Y=17920
X725 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=201360 88880 0 0 $X=201170 $Y=88640
X726 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=206420 12720 1 0 $X=206230 $Y=9760
X727 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=206420 18160 1 0 $X=206230 $Y=15200
X728 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=206880 18160 0 0 $X=206690 $Y=17920
X729 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=206880 88880 0 0 $X=206690 $Y=88640
X730 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=211020 12720 0 0 $X=210830 $Y=12480
X731 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=211940 12720 1 0 $X=211750 $Y=9760
X732 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=212400 18160 0 0 $X=212210 $Y=17920
X733 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=212400 88880 0 0 $X=212210 $Y=88640
X734 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=217920 18160 0 0 $X=217730 $Y=17920
X735 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=217920 88880 0 0 $X=217730 $Y=88640
X736 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=221140 12720 1 0 $X=220950 $Y=9760
X737 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=221140 12720 0 0 $X=220950 $Y=12480
X738 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=221140 18160 1 0 $X=220950 $Y=15200
X739 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=221140 126960 1 0 $X=220950 $Y=124000
X740 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=221140 126960 0 0 $X=220950 $Y=126720
X741 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=223440 18160 0 0 $X=223250 $Y=17920
X742 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=223440 88880 0 0 $X=223250 $Y=88640
X743 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=226660 12720 0 0 $X=226470 $Y=12480
X744 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=226660 126960 1 0 $X=226470 $Y=124000
X745 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=226660 126960 0 0 $X=226470 $Y=126720
X746 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=228960 18160 0 0 $X=228770 $Y=17920
X747 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=228960 88880 0 0 $X=228770 $Y=88640
X748 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=234480 18160 0 0 $X=234290 $Y=17920
X749 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=234480 88880 0 0 $X=234290 $Y=88640
X750 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=235860 12720 1 0 $X=235670 $Y=9760
X751 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=235860 12720 0 0 $X=235670 $Y=12480
X752 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=235860 18160 1 0 $X=235670 $Y=15200
X753 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=240000 18160 0 0 $X=239810 $Y=17920
X754 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=240000 88880 0 0 $X=239810 $Y=88640
X755 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=241380 12720 1 0 $X=241190 $Y=9760
X756 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=241380 18160 1 0 $X=241190 $Y=15200
X757 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=245520 18160 0 0 $X=245330 $Y=17920
X758 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=245520 88880 0 0 $X=245330 $Y=88640
X759 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=250580 18160 1 0 $X=250390 $Y=15200
X760 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=250580 126960 1 0 $X=250390 $Y=124000
X761 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=250580 126960 0 0 $X=250390 $Y=126720
X762 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=251040 18160 0 0 $X=250850 $Y=17920
X763 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=251040 88880 0 0 $X=250850 $Y=88640
X764 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=256100 18160 1 0 $X=255910 $Y=15200
X765 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=256100 126960 1 0 $X=255910 $Y=124000
X766 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=256100 126960 0 0 $X=255910 $Y=126720
X767 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=256560 18160 0 0 $X=256370 $Y=17920
X768 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=256560 88880 0 0 $X=256370 $Y=88640
X769 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=262080 18160 0 0 $X=261890 $Y=17920
X770 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=262080 88880 0 0 $X=261890 $Y=88640
X771 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=265300 12720 1 0 $X=265110 $Y=9760
X772 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=265300 12720 0 0 $X=265110 $Y=12480
X773 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=265300 18160 1 0 $X=265110 $Y=15200
X774 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=267600 18160 0 0 $X=267410 $Y=17920
X775 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=267600 88880 0 0 $X=267410 $Y=88640
X776 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=270820 12720 1 0 $X=270630 $Y=9760
X777 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=270820 12720 0 0 $X=270630 $Y=12480
X778 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=270820 18160 1 0 $X=270630 $Y=15200
X779 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=273120 18160 0 0 $X=272930 $Y=17920
X780 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=273120 88880 0 0 $X=272930 $Y=88640
X781 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=278640 18160 0 0 $X=278450 $Y=17920
X782 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=278640 88880 0 0 $X=278450 $Y=88640
X783 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=280020 12720 1 0 $X=279830 $Y=9760
X784 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=280020 18160 1 0 $X=279830 $Y=15200
X785 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=280020 126960 1 0 $X=279830 $Y=124000
X786 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=280020 126960 0 0 $X=279830 $Y=126720
X787 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=284160 12720 0 0 $X=283970 $Y=12480
X788 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=284160 18160 0 0 $X=283970 $Y=17920
X789 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=284160 88880 0 0 $X=283970 $Y=88640
X790 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=285540 12720 1 0 $X=285350 $Y=9760
X791 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=285540 126960 1 0 $X=285350 $Y=124000
X792 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=285540 126960 0 0 $X=285350 $Y=126720
X793 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=289680 18160 0 0 $X=289490 $Y=17920
X794 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=289680 88880 0 0 $X=289490 $Y=88640
X795 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=294740 12720 1 0 $X=294550 $Y=9760
X796 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=294740 12720 0 0 $X=294550 $Y=12480
X797 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=294740 18160 1 0 $X=294550 $Y=15200
X798 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=295200 18160 0 0 $X=295010 $Y=17920
X799 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=295200 88880 0 0 $X=295010 $Y=88640
X800 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=300260 12720 0 0 $X=300070 $Y=12480
X801 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=300720 18160 0 0 $X=300530 $Y=17920
X802 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=300720 88880 0 0 $X=300530 $Y=88640
X803 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=309460 18160 0 0 $X=309270 $Y=17920
X804 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=309460 88880 1 0 $X=309270 $Y=85920
X805 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=309460 88880 0 0 $X=309270 $Y=88640
X806 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=309460 126960 1 0 $X=309270 $Y=124000
X807 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=309460 126960 0 0 $X=309270 $Y=126720
X808 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=314980 12720 1 0 $X=314790 $Y=9760
X809 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=314980 12720 0 0 $X=314790 $Y=12480
X810 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=314980 18160 0 0 $X=314790 $Y=17920
X811 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=314980 88880 1 0 $X=314790 $Y=85920
X812 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=314980 88880 0 0 $X=314790 $Y=88640
X813 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=314980 126960 1 0 $X=314790 $Y=124000
X814 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=314980 126960 0 0 $X=314790 $Y=126720
X815 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=322340 12720 0 0 $X=322150 $Y=12480
X816 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=322340 50800 1 0 $X=322150 $Y=47840
X817 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=324180 126960 0 0 $X=323990 $Y=126720
X818 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=327860 12720 0 0 $X=327670 $Y=12480
X819 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=327860 50800 1 0 $X=327670 $Y=47840
X820 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=329700 126960 0 0 $X=329510 $Y=126720
X821 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=333380 12720 0 0 $X=333190 $Y=12480
X822 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=333380 50800 1 0 $X=333190 $Y=47840
X823 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=338900 12720 0 0 $X=338710 $Y=12480
X824 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=338900 50800 1 0 $X=338710 $Y=47840
X825 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=338900 126960 0 0 $X=338710 $Y=126720
X826 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=344420 126960 0 0 $X=344230 $Y=126720
X827 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=353620 12720 1 0 $X=353430 $Y=9760
X828 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=353620 45360 0 0 $X=353430 $Y=45120
X829 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=359140 12720 1 0 $X=358950 $Y=9760
X830 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=359140 45360 0 0 $X=358950 $Y=45120
X831 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=368340 12720 1 0 $X=368150 $Y=9760
X832 2 3 3 2 sky130_fd_sc_hd__decap_12 $T=368340 45360 0 0 $X=368150 $Y=45120
X833 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=15060 12720 0 0 $X=14870 $Y=12480
X834 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=15060 34480 1 0 $X=14870 $Y=31520
X835 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=26100 12720 1 0 $X=25910 $Y=9760
X836 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=26100 121520 0 0 $X=25910 $Y=121280
X837 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=26100 126960 1 0 $X=25910 $Y=124000
X838 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=26100 126960 0 0 $X=25910 $Y=126720
X839 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=53240 12720 0 0 $X=53050 $Y=12480
X840 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=55540 12720 1 0 $X=55350 $Y=9760
X841 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=70260 12720 1 0 $X=70070 $Y=9760
X842 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=73940 34480 0 0 $X=73750 $Y=34240
X843 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=73940 39920 1 0 $X=73750 $Y=36960
X844 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=73940 39920 0 0 $X=73750 $Y=39680
X845 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=75780 34480 0 0 $X=75590 $Y=34240
X846 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=75780 39920 1 0 $X=75590 $Y=36960
X847 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=75780 39920 0 0 $X=75590 $Y=39680
X848 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 12720 1 0 $X=84790 $Y=9760
X849 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 56240 0 0 $X=84790 $Y=56000
X850 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 61680 1 0 $X=84790 $Y=58720
X851 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 61680 0 0 $X=84790 $Y=61440
X852 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 67120 1 0 $X=84790 $Y=64160
X853 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 67120 0 0 $X=84790 $Y=66880
X854 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 72560 1 0 $X=84790 $Y=69600
X855 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 72560 0 0 $X=84790 $Y=72320
X856 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 78000 1 0 $X=84790 $Y=75040
X857 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 78000 0 0 $X=84790 $Y=77760
X858 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 83440 1 0 $X=84790 $Y=80480
X859 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 83440 0 0 $X=84790 $Y=83200
X860 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 88880 1 0 $X=84790 $Y=85920
X861 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 88880 0 0 $X=84790 $Y=88640
X862 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 94320 1 0 $X=84790 $Y=91360
X863 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 94320 0 0 $X=84790 $Y=94080
X864 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 99760 1 0 $X=84790 $Y=96800
X865 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 99760 0 0 $X=84790 $Y=99520
X866 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 105200 1 0 $X=84790 $Y=102240
X867 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 105200 0 0 $X=84790 $Y=104960
X868 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 110640 1 0 $X=84790 $Y=107680
X869 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 110640 0 0 $X=84790 $Y=110400
X870 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 116080 1 0 $X=84790 $Y=113120
X871 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 116080 0 0 $X=84790 $Y=115840
X872 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 121520 1 0 $X=84790 $Y=118560
X873 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 121520 0 0 $X=84790 $Y=121280
X874 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 126960 1 0 $X=84790 $Y=124000
X875 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=84980 126960 0 0 $X=84790 $Y=126720
X876 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=87280 12720 0 0 $X=87090 $Y=12480
X877 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=93720 23600 0 0 $X=93530 $Y=23360
X878 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=99700 12720 1 0 $X=99510 $Y=9760
X879 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=99700 61680 0 0 $X=99510 $Y=61440
X880 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=111660 12720 0 0 $X=111470 $Y=12480
X881 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=111660 18160 1 0 $X=111470 $Y=15200
X882 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=114420 12720 1 0 $X=114230 $Y=9760
X883 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=114420 126960 1 0 $X=114230 $Y=124000
X884 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=114420 126960 0 0 $X=114230 $Y=126720
X885 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=122240 18160 1 0 $X=122050 $Y=15200
X886 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=129140 12720 1 0 $X=128950 $Y=9760
X887 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=129140 12720 0 0 $X=128950 $Y=12480
X888 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 12720 0 0 $X=143670 $Y=12480
X889 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 18160 1 0 $X=143670 $Y=15200
X890 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 94320 1 0 $X=143670 $Y=91360
X891 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 94320 0 0 $X=143670 $Y=94080
X892 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 99760 1 0 $X=143670 $Y=96800
X893 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 99760 0 0 $X=143670 $Y=99520
X894 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 105200 1 0 $X=143670 $Y=102240
X895 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 105200 0 0 $X=143670 $Y=104960
X896 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 110640 1 0 $X=143670 $Y=107680
X897 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 110640 0 0 $X=143670 $Y=110400
X898 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 116080 1 0 $X=143670 $Y=113120
X899 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 116080 0 0 $X=143670 $Y=115840
X900 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 121520 1 0 $X=143670 $Y=118560
X901 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 121520 0 0 $X=143670 $Y=121280
X902 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 126960 1 0 $X=143670 $Y=124000
X903 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=143860 126960 0 0 $X=143670 $Y=126720
X904 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=145240 12720 1 0 $X=145050 $Y=9760
X905 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=158580 12720 1 0 $X=158390 $Y=9760
X906 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=158580 12720 0 0 $X=158390 $Y=12480
X907 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=158580 18160 1 0 $X=158390 $Y=15200
X908 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=167780 12720 0 0 $X=167590 $Y=12480
X909 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=173300 18160 1 0 $X=173110 $Y=15200
X910 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=173300 126960 1 0 $X=173110 $Y=124000
X911 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=173300 126960 0 0 $X=173110 $Y=126720
X912 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=189400 18160 1 0 $X=189210 $Y=15200
X913 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=199980 12720 1 0 $X=199790 $Y=9760
X914 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=199980 18160 1 0 $X=199790 $Y=15200
X915 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 94320 1 0 $X=202550 $Y=91360
X916 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 94320 0 0 $X=202550 $Y=94080
X917 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 99760 1 0 $X=202550 $Y=96800
X918 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 99760 0 0 $X=202550 $Y=99520
X919 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 105200 1 0 $X=202550 $Y=102240
X920 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 105200 0 0 $X=202550 $Y=104960
X921 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 110640 1 0 $X=202550 $Y=107680
X922 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 110640 0 0 $X=202550 $Y=110400
X923 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 116080 1 0 $X=202550 $Y=113120
X924 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 116080 0 0 $X=202550 $Y=115840
X925 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 121520 1 0 $X=202550 $Y=118560
X926 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 121520 0 0 $X=202550 $Y=121280
X927 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 126960 1 0 $X=202550 $Y=124000
X928 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=202740 126960 0 0 $X=202550 $Y=126720
X929 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=214700 18160 1 0 $X=214510 $Y=15200
X930 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=217460 12720 1 0 $X=217270 $Y=9760
X931 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=226660 12720 1 0 $X=226470 $Y=9760
X932 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=232180 12720 0 0 $X=231990 $Y=12480
X933 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=232180 126960 1 0 $X=231990 $Y=124000
X934 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=232180 126960 0 0 $X=231990 $Y=126720
X935 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=246900 12720 1 0 $X=246710 $Y=9760
X936 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=246900 18160 1 0 $X=246710 $Y=15200
X937 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=248280 12720 0 0 $X=248090 $Y=12480
X938 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 18160 1 0 $X=261430 $Y=15200
X939 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 94320 1 0 $X=261430 $Y=91360
X940 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 94320 0 0 $X=261430 $Y=94080
X941 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 99760 1 0 $X=261430 $Y=96800
X942 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 99760 0 0 $X=261430 $Y=99520
X943 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 105200 1 0 $X=261430 $Y=102240
X944 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 105200 0 0 $X=261430 $Y=104960
X945 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 110640 1 0 $X=261430 $Y=107680
X946 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 110640 0 0 $X=261430 $Y=110400
X947 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 116080 1 0 $X=261430 $Y=113120
X948 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 116080 0 0 $X=261430 $Y=115840
X949 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 121520 1 0 $X=261430 $Y=118560
X950 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 121520 0 0 $X=261430 $Y=121280
X951 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 126960 1 0 $X=261430 $Y=124000
X952 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=261620 126960 0 0 $X=261430 $Y=126720
X953 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=263000 12720 1 0 $X=262810 $Y=9760
X954 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=263000 12720 0 0 $X=262810 $Y=12480
X955 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=276340 12720 1 0 $X=276150 $Y=9760
X956 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=276340 12720 0 0 $X=276150 $Y=12480
X957 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=276340 18160 1 0 $X=276150 $Y=15200
X958 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=288300 18160 1 0 $X=288110 $Y=15200
X959 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=291060 12720 1 0 $X=290870 $Y=9760
X960 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=291060 126960 1 0 $X=290870 $Y=124000
X961 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=291060 126960 0 0 $X=290870 $Y=126720
X962 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=292440 12720 0 0 $X=292250 $Y=12480
X963 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=305780 12720 0 0 $X=305590 $Y=12480
X964 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=307160 12720 1 0 $X=306970 $Y=9760
X965 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=307160 18160 1 0 $X=306970 $Y=15200
X966 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=312220 18160 1 0 $X=312030 $Y=15200
X967 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 12720 1 0 $X=320310 $Y=9760
X968 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 50800 0 0 $X=320310 $Y=50560
X969 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 56240 1 0 $X=320310 $Y=53280
X970 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 56240 0 0 $X=320310 $Y=56000
X971 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 61680 1 0 $X=320310 $Y=58720
X972 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 61680 0 0 $X=320310 $Y=61440
X973 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 67120 1 0 $X=320310 $Y=64160
X974 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 67120 0 0 $X=320310 $Y=66880
X975 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 72560 1 0 $X=320310 $Y=69600
X976 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 72560 0 0 $X=320310 $Y=72320
X977 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 78000 1 0 $X=320310 $Y=75040
X978 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 78000 0 0 $X=320310 $Y=77760
X979 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 83440 1 0 $X=320310 $Y=80480
X980 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 83440 0 0 $X=320310 $Y=83200
X981 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 88880 1 0 $X=320310 $Y=85920
X982 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 88880 0 0 $X=320310 $Y=88640
X983 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 94320 1 0 $X=320310 $Y=91360
X984 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 94320 0 0 $X=320310 $Y=94080
X985 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 99760 1 0 $X=320310 $Y=96800
X986 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 99760 0 0 $X=320310 $Y=99520
X987 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 105200 1 0 $X=320310 $Y=102240
X988 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 105200 0 0 $X=320310 $Y=104960
X989 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 110640 1 0 $X=320310 $Y=107680
X990 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 110640 0 0 $X=320310 $Y=110400
X991 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 116080 1 0 $X=320310 $Y=113120
X992 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 116080 0 0 $X=320310 $Y=115840
X993 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 121520 1 0 $X=320310 $Y=118560
X994 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 121520 0 0 $X=320310 $Y=121280
X995 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 126960 1 0 $X=320310 $Y=124000
X996 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=320500 126960 0 0 $X=320310 $Y=126720
X997 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=335220 126960 0 0 $X=335030 $Y=126720
X998 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=349940 12720 1 0 $X=349750 $Y=9760
X999 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=349940 126960 0 0 $X=349750 $Y=126720
X1000 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 18160 1 0 $X=351130 $Y=15200
X1001 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 18160 0 0 $X=351130 $Y=17920
X1002 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 23600 1 0 $X=351130 $Y=20640
X1003 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 23600 0 0 $X=351130 $Y=23360
X1004 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 29040 1 0 $X=351130 $Y=26080
X1005 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 29040 0 0 $X=351130 $Y=28800
X1006 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 34480 1 0 $X=351130 $Y=31520
X1007 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 34480 0 0 $X=351130 $Y=34240
X1008 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 39920 1 0 $X=351130 $Y=36960
X1009 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 39920 0 0 $X=351130 $Y=39680
X1010 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 45360 1 0 $X=351130 $Y=42400
X1011 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=351320 45360 0 0 $X=351130 $Y=45120
X1012 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=364660 12720 1 0 $X=364470 $Y=9760
X1013 2 3 3 2 sky130_fd_sc_hd__decap_4 $T=364660 45360 0 0 $X=364470 $Y=45120
X1014 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=29780 12720 1 0 $X=29590 $Y=9760
X1015 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=31160 18160 1 0 $X=30970 $Y=15200
X1016 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=31160 18160 0 0 $X=30970 $Y=17920
X1017 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=31160 23600 1 0 $X=30970 $Y=20640
X1018 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=31160 23600 0 0 $X=30970 $Y=23360
X1019 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=31160 29040 1 0 $X=30970 $Y=26080
X1020 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=31160 29040 0 0 $X=30970 $Y=28800
X1021 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=31160 34480 1 0 $X=30970 $Y=31520
X1022 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=48180 61680 0 0 $X=47990 $Y=61440
X1023 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=95100 18160 1 0 $X=94910 $Y=15200
X1024 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=96480 12720 0 0 $X=96290 $Y=12480
X1025 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=96480 18160 0 0 $X=96290 $Y=17920
X1026 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=96480 23600 1 0 $X=96290 $Y=20640
X1027 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=96480 45360 1 0 $X=96290 $Y=42400
X1028 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=191700 12720 0 0 $X=191510 $Y=12480
X1029 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=226660 18160 1 0 $X=226470 $Y=15200
X1030 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=318200 18160 1 0 $X=318010 $Y=15200
X1031 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=324180 12720 1 0 $X=323990 $Y=9760
X1032 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=334760 12720 1 0 $X=334570 $Y=9760
X1033 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=344420 12720 0 0 $X=344230 $Y=12480
X1034 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=344420 50800 1 0 $X=344230 $Y=47840
X1035 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 12720 1 0 $X=373670 $Y=9760
X1036 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 12720 0 0 $X=373670 $Y=12480
X1037 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 18160 1 0 $X=373670 $Y=15200
X1038 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 18160 0 0 $X=373670 $Y=17920
X1039 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 23600 1 0 $X=373670 $Y=20640
X1040 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 23600 0 0 $X=373670 $Y=23360
X1041 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 29040 1 0 $X=373670 $Y=26080
X1042 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 29040 0 0 $X=373670 $Y=28800
X1043 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 34480 1 0 $X=373670 $Y=31520
X1044 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 34480 0 0 $X=373670 $Y=34240
X1045 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 39920 1 0 $X=373670 $Y=36960
X1046 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 39920 0 0 $X=373670 $Y=39680
X1047 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 45360 1 0 $X=373670 $Y=42400
X1048 2 3 3 2 sky130_fd_sc_hd__decap_8 $T=373860 45360 0 0 $X=373670 $Y=45120
X1049 2 3 3 2 sky130_fd_sc_hd__fill_2 $T=43120 12720 1 0 $X=42930 $Y=9760
X1050 2 3 3 2 sky130_fd_sc_hd__fill_2 $T=205040 12720 0 0 $X=204850 $Y=12480
X1051 2 3 3 2 sky130_fd_sc_hd__fill_2 $T=234480 18160 1 0 $X=234290 $Y=15200
X1052 2 3 3 2 sky130_fd_sc_hd__fill_2 $T=352240 50800 1 0 $X=352050 $Y=47840
X1053 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16440 18160 1 0 $X=16250 $Y=15200
X1054 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16440 18160 0 0 $X=16250 $Y=17920
X1055 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16440 23600 1 0 $X=16250 $Y=20640
X1056 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16440 23600 0 0 $X=16250 $Y=23360
X1057 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16440 29040 1 0 $X=16250 $Y=26080
X1058 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16440 29040 0 0 $X=16250 $Y=28800
X1059 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16900 18160 1 0 $X=16710 $Y=15200
X1060 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16900 18160 0 0 $X=16710 $Y=17920
X1061 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16900 23600 1 0 $X=16710 $Y=20640
X1062 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16900 23600 0 0 $X=16710 $Y=23360
X1063 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16900 29040 1 0 $X=16710 $Y=26080
X1064 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=16900 29040 0 0 $X=16710 $Y=28800
X1065 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=30240 18160 1 0 $X=30050 $Y=15200
X1066 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=30240 18160 0 0 $X=30050 $Y=17920
X1067 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=30240 23600 1 0 $X=30050 $Y=20640
X1068 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=30240 23600 0 0 $X=30050 $Y=23360
X1069 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=30240 29040 1 0 $X=30050 $Y=26080
X1070 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=30240 29040 0 0 $X=30050 $Y=28800
X1071 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 34480 0 0 $X=36950 $Y=34240
X1072 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 39920 1 0 $X=36950 $Y=36960
X1073 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 39920 0 0 $X=36950 $Y=39680
X1074 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 45360 1 0 $X=36950 $Y=42400
X1075 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 45360 0 0 $X=36950 $Y=45120
X1076 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 50800 1 0 $X=36950 $Y=47840
X1077 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 50800 0 0 $X=36950 $Y=50560
X1078 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 56240 1 0 $X=36950 $Y=53280
X1079 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 56240 0 0 $X=36950 $Y=56000
X1080 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=37140 61680 1 0 $X=36950 $Y=58720
X1081 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 18160 1 0 $X=52590 $Y=15200
X1082 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 18160 0 0 $X=52590 $Y=17920
X1083 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 23600 1 0 $X=52590 $Y=20640
X1084 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 23600 0 0 $X=52590 $Y=23360
X1085 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 29040 1 0 $X=52590 $Y=26080
X1086 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 29040 0 0 $X=52590 $Y=28800
X1087 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 34480 1 0 $X=52590 $Y=31520
X1088 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 34480 0 0 $X=52590 $Y=34240
X1089 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 39920 1 0 $X=52590 $Y=36960
X1090 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 39920 0 0 $X=52590 $Y=39680
X1091 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 45360 1 0 $X=52590 $Y=42400
X1092 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 45360 0 0 $X=52590 $Y=45120
X1093 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 50800 1 0 $X=52590 $Y=47840
X1094 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 50800 0 0 $X=52590 $Y=50560
X1095 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 56240 1 0 $X=52590 $Y=53280
X1096 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 56240 0 0 $X=52590 $Y=56000
X1097 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=52780 61680 1 0 $X=52590 $Y=58720
X1098 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=53240 18160 1 0 $X=53050 $Y=15200
X1099 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=53240 18160 0 0 $X=53050 $Y=17920
X1100 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=53240 23600 1 0 $X=53050 $Y=20640
X1101 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=53240 23600 0 0 $X=53050 $Y=23360
X1102 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=53240 29040 1 0 $X=53050 $Y=26080
X1103 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=53240 29040 0 0 $X=53050 $Y=28800
X1104 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=53240 34480 1 0 $X=53050 $Y=31520
X1105 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=56920 18160 1 0 $X=56730 $Y=15200
X1106 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=56920 18160 0 0 $X=56730 $Y=17920
X1107 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=56920 23600 1 0 $X=56730 $Y=20640
X1108 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=56920 23600 0 0 $X=56730 $Y=23360
X1109 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=56920 29040 1 0 $X=56730 $Y=26080
X1110 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=56920 29040 0 0 $X=56730 $Y=28800
X1111 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 18160 1 0 $X=89850 $Y=15200
X1112 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 18160 0 0 $X=89850 $Y=17920
X1113 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 23600 1 0 $X=89850 $Y=20640
X1114 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 23600 0 0 $X=89850 $Y=23360
X1115 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 29040 1 0 $X=89850 $Y=26080
X1116 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 29040 0 0 $X=89850 $Y=28800
X1117 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 34480 1 0 $X=89850 $Y=31520
X1118 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 34480 0 0 $X=89850 $Y=34240
X1119 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 39920 1 0 $X=89850 $Y=36960
X1120 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=90040 39920 0 0 $X=89850 $Y=39680
X1121 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=99700 23600 0 0 $X=99510 $Y=23360
X1122 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 23600 1 0 $X=101810 $Y=20640
X1123 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 23600 0 0 $X=101810 $Y=23360
X1124 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 29040 1 0 $X=101810 $Y=26080
X1125 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 29040 0 0 $X=101810 $Y=28800
X1126 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 34480 1 0 $X=101810 $Y=31520
X1127 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 34480 0 0 $X=101810 $Y=34240
X1128 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 39920 1 0 $X=101810 $Y=36960
X1129 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 39920 0 0 $X=101810 $Y=39680
X1130 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 45360 1 0 $X=101810 $Y=42400
X1131 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 45360 0 0 $X=101810 $Y=45120
X1132 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 50800 1 0 $X=101810 $Y=47840
X1133 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 50800 0 0 $X=101810 $Y=50560
X1134 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 56240 1 0 $X=101810 $Y=53280
X1135 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 56240 0 0 $X=101810 $Y=56000
X1136 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 61680 1 0 $X=101810 $Y=58720
X1137 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 61680 0 0 $X=101810 $Y=61440
X1138 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 67120 1 0 $X=101810 $Y=64160
X1139 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 67120 0 0 $X=101810 $Y=66880
X1140 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 72560 1 0 $X=101810 $Y=69600
X1141 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 72560 0 0 $X=101810 $Y=72320
X1142 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 78000 1 0 $X=101810 $Y=75040
X1143 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 78000 0 0 $X=101810 $Y=77760
X1144 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 83440 1 0 $X=101810 $Y=80480
X1145 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 83440 0 0 $X=101810 $Y=83200
X1146 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=102000 88880 1 0 $X=101810 $Y=85920
X1147 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=176060 12720 1 0 $X=175870 $Y=9760
X1148 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=206420 12720 0 0 $X=206230 $Y=12480
X1149 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 18160 1 0 $X=322150 $Y=15200
X1150 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 18160 0 0 $X=322150 $Y=17920
X1151 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 23600 1 0 $X=322150 $Y=20640
X1152 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 23600 0 0 $X=322150 $Y=23360
X1153 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 29040 1 0 $X=322150 $Y=26080
X1154 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 29040 0 0 $X=322150 $Y=28800
X1155 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 34480 1 0 $X=322150 $Y=31520
X1156 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 34480 0 0 $X=322150 $Y=34240
X1157 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 39920 1 0 $X=322150 $Y=36960
X1158 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 39920 0 0 $X=322150 $Y=39680
X1159 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 45360 1 0 $X=322150 $Y=42400
X1160 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=322340 45360 0 0 $X=322150 $Y=45120
X1161 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 18160 1 0 $X=350210 $Y=15200
X1162 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 18160 0 0 $X=350210 $Y=17920
X1163 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 23600 1 0 $X=350210 $Y=20640
X1164 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 23600 0 0 $X=350210 $Y=23360
X1165 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 29040 1 0 $X=350210 $Y=26080
X1166 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 29040 0 0 $X=350210 $Y=28800
X1167 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 34480 1 0 $X=350210 $Y=31520
X1168 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 34480 0 0 $X=350210 $Y=34240
X1169 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 39920 1 0 $X=350210 $Y=36960
X1170 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 39920 0 0 $X=350210 $Y=39680
X1171 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 45360 1 0 $X=350210 $Y=42400
X1172 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350400 45360 0 0 $X=350210 $Y=45120
X1173 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 18160 1 0 $X=350670 $Y=15200
X1174 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 18160 0 0 $X=350670 $Y=17920
X1175 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 23600 1 0 $X=350670 $Y=20640
X1176 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 23600 0 0 $X=350670 $Y=23360
X1177 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 29040 1 0 $X=350670 $Y=26080
X1178 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 29040 0 0 $X=350670 $Y=28800
X1179 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 34480 1 0 $X=350670 $Y=31520
X1180 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 34480 0 0 $X=350670 $Y=34240
X1181 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 39920 1 0 $X=350670 $Y=36960
X1182 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 39920 0 0 $X=350670 $Y=39680
X1183 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 45360 1 0 $X=350670 $Y=42400
X1184 2 3 3 2 sky130_fd_sc_hd__fill_1 $T=350860 45360 0 0 $X=350670 $Y=45120
X1185 6 M2M3_PR $T=23110 22980 0 0 $X=22945 $Y=22795
X1186 10 M2M3_PR $T=35990 2240 0 0 $X=35825 $Y=2055
X1187 6 M2M3_PR $T=54390 22980 0 0 $X=54225 $Y=22795
X1188 5 M2M3_PR $T=54390 51650 0 0 $X=54225 $Y=51465
X1189 7 M2M3_PR $T=57610 22980 0 0 $X=57445 $Y=22795
X1190 150 M2M3_PR $T=88890 8950 0 0 $X=88725 $Y=8765
X1191 123 M2M3_PR $T=90730 1020 0 0 $X=90565 $Y=835
X1192 119 M2M3_PR $T=94410 14440 0 0 $X=94245 $Y=14255
X1193 7 M2M3_PR $T=94870 22980 0 0 $X=94705 $Y=22795
X1194 5 M2M3_PR $T=98550 51650 0 0 $X=98385 $Y=51465
X1195 8 M2M3_PR $T=101770 1020 0 0 $X=101605 $Y=835
X1196 9 M2M3_PR $T=105450 43720 0 0 $X=105285 $Y=43535
X1197 149 M2M3_PR $T=109590 2240 0 0 $X=109425 $Y=2055
X1198 151 M2M3_PR $T=113270 4680 0 0 $X=113105 $Y=4495
X1199 151 M2M3_PR $T=113270 18100 0 0 $X=113105 $Y=17915
X1200 13 M2M3_PR $T=116490 26630 0 0 $X=116325 $Y=26445
X1201 151 M2M3_PR $T=116950 18100 0 0 $X=116785 $Y=17915
X1202 119 M2M3_PR $T=124310 14440 0 0 $X=124145 $Y=14255
X1203 37 M2M3_PR $T=148690 60190 0 0 $X=148525 $Y=60005
X1204 155 M2M3_PR $T=153290 2850 0 0 $X=153125 $Y=2665
X1205 22 M2M3_PR $T=153750 18710 0 0 $X=153585 $Y=18525
X1206 37 M2M3_PR $T=164790 60190 0 0 $X=164625 $Y=60005
X1207 125 M2M3_PR $T=167550 2240 0 0 $X=167385 $Y=2055
X1208 132 M2M3_PR $T=178130 9560 0 0 $X=177965 $Y=9375
X1209 129 M2M3_PR $T=183190 4680 0 0 $X=183025 $Y=4495
X1210 26 M2M3_PR $T=186870 28470 0 0 $X=186705 $Y=28285
X1211 30 M2M3_PR $T=201130 13830 0 0 $X=200965 $Y=13645
X1212 132 M2M3_PR $T=204350 9560 0 0 $X=204185 $Y=9375
X1213 131 M2M3_PR $T=204810 2240 0 0 $X=204645 $Y=2055
X1214 119 M2M3_PR $T=216310 18100 0 0 $X=216145 $Y=17915
X1215 32 M2M3_PR $T=231030 27860 0 0 $X=230865 $Y=27675
X1216 136 M2M3_PR $T=234250 8950 0 0 $X=234085 $Y=8765
X1217 34 M2M3_PR $T=253110 22370 0 0 $X=252945 $Y=22185
X1218 1 M2M3_PR $T=255410 7730 0 0 $X=255245 $Y=7545
X1219 112 M2M3_PR $T=256790 14440 0 0 $X=256625 $Y=14255
X1220 42 M2M3_PR $T=258630 22370 0 0 $X=258465 $Y=22185
X1221 138 M2M3_PR $T=259550 2240 0 0 $X=259385 $Y=2055
X1222 43 M2M3_PR $T=272890 34570 0 0 $X=272725 $Y=34385
X1223 42 M2M3_PR $T=282090 22370 0 0 $X=281925 $Y=22185
X1224 1 M2M3_PR $T=292670 8340 0 0 $X=292505 $Y=8155
X1225 112 M2M3_PR $T=293130 13830 0 0 $X=292965 $Y=13645
X1226 142 M2M3_PR $T=300950 2850 0 0 $X=300785 $Y=2665
X1227 1 M2M3_PR $T=304170 8340 0 0 $X=304005 $Y=8155
X1228 43 M2M3_PR $T=307850 34570 0 0 $X=307685 $Y=34385
X1229 144 M2M3_PR $T=315670 2240 0 0 $X=315505 $Y=2055
X1230 39 M2M3_PR $T=315670 27250 0 0 $X=315505 $Y=27065
X1231 108 M2M3_PR $T=322570 26640 0 0 $X=322405 $Y=26455
X1232 104 M2M3_PR $T=323490 35180 0 0 $X=323325 $Y=34995
X1233 41 M2M3_PR $T=326250 9560 0 0 $X=326085 $Y=9375
X1234 119 M2M3_PR $T=329010 18100 0 0 $X=328845 $Y=17915
X1235 145 M2M3_PR $T=330390 10780 0 0 $X=330225 $Y=10595
X1236 104 M2M3_PR $T=336370 35180 0 0 $X=336205 $Y=34995
X1237 108 M2M3_PR $T=338210 26640 0 0 $X=338045 $Y=26455
X1238 8 M2M3_PR $T=346030 1020 0 0 $X=345865 $Y=835
X1239 146 M2M3_PR $T=348330 1020 0 0 $X=348165 $Y=835
X1240 147 M2M3_PR $T=352010 2850 0 0 $X=351845 $Y=2665
X1241 141 M1M2_PR $T=10230 650 0 0 $X=10070 $Y=490
X1242 6 M1M2_PR $T=23110 23770 0 0 $X=22950 $Y=23610
X1243 148 M1M2_PR $T=27710 16970 0 0 $X=27550 $Y=16810
X1244 10 M1M2_PR $T=35990 11190 0 0 $X=35830 $Y=11030
X1245 152 M1M2_PR $T=43350 14250 0 0 $X=43190 $Y=14090
X1246 11 M1M2_PR $T=45650 30230 0 0 $X=45490 $Y=30070
X1247 11 M1M2_PR $T=46570 6770 0 0 $X=46410 $Y=6610
X1248 11 M1M2_PR $T=46570 11530 0 0 $X=46410 $Y=11370
X1249 121 M1M2_PR $T=47030 25470 0 0 $X=46870 $Y=25310
X1250 4 M1M2_PR $T=50710 50630 0 0 $X=50550 $Y=50470
X1251 4 M1M2_PR $T=50710 52670 0 0 $X=50550 $Y=52510
X1252 6 M1M2_PR $T=54390 24110 0 0 $X=54230 $Y=23950
X1253 5 M1M2_PR $T=54390 51990 0 0 $X=54230 $Y=51830
X1254 7 M1M2_PR $T=57610 24790 0 0 $X=57450 $Y=24630
X1255 120 M1M2_PR $T=57610 34990 0 0 $X=57450 $Y=34830
X1256 120 M1M2_PR $T=58530 23770 0 0 $X=58370 $Y=23610
X1257 153 M1M2_PR $T=60830 3030 0 0 $X=60670 $Y=2870
X1258 122 M1M2_PR $T=70950 1670 0 0 $X=70790 $Y=1510
X1259 122 M1M2_PR $T=70950 30910 0 0 $X=70790 $Y=30750
X1260 86 M1M2_PR $T=72790 25130 0 0 $X=72630 $Y=24970
X1261 86 M1M2_PR $T=72790 33290 0 0 $X=72630 $Y=33130
X1262 154 M1M2_PR $T=79690 11530 0 0 $X=79530 $Y=11370
X1263 37 M1M2_PR $T=83830 60150 0 0 $X=83670 $Y=59990
X1264 37 M1M2_PR $T=84290 23090 0 0 $X=84130 $Y=22930
X1265 150 M1M2_PR $T=88890 17650 0 0 $X=88730 $Y=17490
X1266 123 M1M2_PR $T=90730 16290 0 0 $X=90570 $Y=16130
X1267 124 M1M2_PR $T=94410 8470 0 0 $X=94250 $Y=8310
X1268 119 M1M2_PR $T=94410 15950 0 0 $X=94250 $Y=15790
X1269 7 M1M2_PR $T=94870 24110 0 0 $X=94710 $Y=23950
X1270 5 M1M2_PR $T=98550 24110 0 0 $X=98390 $Y=23950
X1271 5 M1M2_PR $T=98550 24790 0 0 $X=98390 $Y=24630
X1272 8 M1M2_PR $T=101770 25130 0 0 $X=101610 $Y=24970
X1273 9 M1M2_PR $T=105450 25810 0 0 $X=105290 $Y=25650
X1274 149 M1M2_PR $T=109590 13230 0 0 $X=109430 $Y=13070
X1275 126 M1M2_PR $T=112810 13570 0 0 $X=112650 $Y=13410
X1276 123 M1M2_PR $T=112810 14250 0 0 $X=112650 $Y=14090
X1277 123 M1M2_PR $T=112810 16290 0 0 $X=112650 $Y=16130
X1278 14 M1M2_PR $T=116490 16970 0 0 $X=116330 $Y=16810
X1279 13 M1M2_PR $T=116490 17650 0 0 $X=116330 $Y=17490
X1280 16 M1M2_PR $T=116950 12210 0 0 $X=116790 $Y=12050
X1281 16 M1M2_PR $T=116950 14250 0 0 $X=116790 $Y=14090
X1282 151 M1M2_PR $T=116950 17650 0 0 $X=116790 $Y=17490
X1283 123 M1M2_PR $T=120170 13910 0 0 $X=120010 $Y=13750
X1284 123 M1M2_PR $T=120170 16630 0 0 $X=120010 $Y=16470
X1285 18 M1M2_PR $T=120170 17310 0 0 $X=120010 $Y=17150
X1286 18 M1M2_PR $T=120170 19690 0 0 $X=120010 $Y=19530
X1287 91 M1M2_PR $T=120170 27170 0 0 $X=120010 $Y=27010
X1288 91 M1M2_PR $T=120630 14930 0 0 $X=120470 $Y=14770
X1289 89 M1M2_PR $T=123850 5410 0 0 $X=123690 $Y=5250
X1290 89 M1M2_PR $T=123850 15950 0 0 $X=123690 $Y=15790
X1291 93 M1M2_PR $T=123850 16970 0 0 $X=123690 $Y=16810
X1292 93 M1M2_PR $T=123850 24790 0 0 $X=123690 $Y=24630
X1293 93 M1M2_PR $T=123850 26150 0 0 $X=123690 $Y=25990
X1294 93 M1M2_PR $T=123850 30570 0 0 $X=123690 $Y=30410
X1295 119 M1M2_PR $T=124310 15950 0 0 $X=124150 $Y=15790
X1296 15 M1M2_PR $T=124310 17650 0 0 $X=124150 $Y=17490
X1297 123 M1M2_PR $T=127530 13910 0 0 $X=127370 $Y=13750
X1298 88 M1M2_PR $T=127530 17650 0 0 $X=127370 $Y=17490
X1299 88 M1M2_PR $T=127530 28190 0 0 $X=127370 $Y=28030
X1300 127 M1M2_PR $T=127990 7790 0 0 $X=127830 $Y=7630
X1301 152 M1M2_PR $T=127990 14590 0 0 $X=127830 $Y=14430
X1302 123 M1M2_PR $T=127990 16630 0 0 $X=127830 $Y=16470
X1303 152 M1M2_PR $T=127990 17310 0 0 $X=127830 $Y=17150
X1304 153 M1M2_PR $T=130750 4050 0 0 $X=130590 $Y=3890
X1305 16 M1M2_PR $T=131210 12210 0 0 $X=131050 $Y=12050
X1306 153 M1M2_PR $T=131210 17310 0 0 $X=131050 $Y=17150
X1307 17 M1M2_PR $T=134890 17650 0 0 $X=134730 $Y=17490
X1308 123 M1M2_PR $T=135350 10850 0 0 $X=135190 $Y=10690
X1309 123 M1M2_PR $T=135350 14250 0 0 $X=135190 $Y=14090
X1310 123 M1M2_PR $T=135350 16290 0 0 $X=135190 $Y=16130
X1311 154 M1M2_PR $T=138570 12210 0 0 $X=138410 $Y=12050
X1312 154 M1M2_PR $T=138570 13230 0 0 $X=138410 $Y=13070
X1313 90 M1M2_PR $T=138570 15950 0 0 $X=138410 $Y=15790
X1314 90 M1M2_PR $T=138570 32610 0 0 $X=138410 $Y=32450
X1315 18 M1M2_PR $T=139490 20030 0 0 $X=139330 $Y=19870
X1316 124 M1M2_PR $T=142710 9150 0 0 $X=142550 $Y=8990
X1317 124 M1M2_PR $T=142710 11530 0 0 $X=142550 $Y=11370
X1318 19 M1M2_PR $T=142710 14250 0 0 $X=142550 $Y=14090
X1319 128 M1M2_PR $T=144550 9490 0 0 $X=144390 $Y=9330
X1320 21 M1M2_PR $T=145930 11870 0 0 $X=145770 $Y=11710
X1321 37 M1M2_PR $T=148690 60490 0 0 $X=148530 $Y=60330
X1322 155 M1M2_PR $T=153290 17650 0 0 $X=153130 $Y=17490
X1323 22 M1M2_PR $T=153750 16630 0 0 $X=153590 $Y=16470
X1324 92 M1M2_PR $T=156970 14930 0 0 $X=156810 $Y=14770
X1325 92 M1M2_PR $T=156970 25810 0 0 $X=156810 $Y=25650
X1326 23 M1M2_PR $T=161110 14250 0 0 $X=160950 $Y=14090
X1327 130 M1M2_PR $T=161570 8470 0 0 $X=161410 $Y=8310
X1328 95 M1M2_PR $T=164790 15950 0 0 $X=164630 $Y=15790
X1329 95 M1M2_PR $T=164790 31250 0 0 $X=164630 $Y=31090
X1330 37 M1M2_PR $T=164790 60490 0 0 $X=164630 $Y=60330
X1331 125 M1M2_PR $T=168010 17310 0 0 $X=167850 $Y=17150
X1332 123 M1M2_PR $T=168470 14930 0 0 $X=168310 $Y=14770
X1333 123 M1M2_PR $T=168470 16290 0 0 $X=168310 $Y=16130
X1334 24 M1M2_PR $T=168470 17650 0 0 $X=168310 $Y=17490
X1335 97 M1M2_PR $T=169850 3710 0 0 $X=169690 $Y=3550
X1336 97 M1M2_PR $T=170220 15950 0 0 $X=170060 $Y=15790
X1337 128 M1M2_PR $T=171230 9490 0 0 $X=171070 $Y=9330
X1338 127 M1M2_PR $T=171690 7790 0 0 $X=171530 $Y=7630
X1339 127 M1M2_PR $T=171690 11870 0 0 $X=171530 $Y=11710
X1340 128 M1M2_PR $T=171690 17310 0 0 $X=171530 $Y=17150
X1341 25 M1M2_PR $T=172150 12210 0 0 $X=171990 $Y=12050
X1342 123 M1M2_PR $T=175370 11530 0 0 $X=175210 $Y=11370
X1343 123 M1M2_PR $T=175370 14590 0 0 $X=175210 $Y=14430
X1344 123 M1M2_PR $T=175370 15950 0 0 $X=175210 $Y=15790
X1345 100 M1M2_PR $T=179050 17650 0 0 $X=178890 $Y=17490
X1346 100 M1M2_PR $T=179050 28870 0 0 $X=178890 $Y=28710
X1347 28 M1M2_PR $T=182730 17650 0 0 $X=182570 $Y=17490
X1348 129 M1M2_PR $T=183190 17310 0 0 $X=183030 $Y=17150
X1349 26 M1M2_PR $T=186870 17310 0 0 $X=186710 $Y=17150
X1350 130 M1M2_PR $T=190550 9150 0 0 $X=190390 $Y=8990
X1351 130 M1M2_PR $T=190550 13230 0 0 $X=190390 $Y=13070
X1352 96 M1M2_PR $T=190550 14930 0 0 $X=190390 $Y=14770
X1353 96 M1M2_PR $T=190550 32270 0 0 $X=190390 $Y=32110
X1354 94 M1M2_PR $T=194230 11190 0 0 $X=194070 $Y=11030
X1355 94 M1M2_PR $T=194230 33630 0 0 $X=194070 $Y=33470
X1356 133 M1M2_PR $T=197450 13910 0 0 $X=197290 $Y=13750
X1357 99 M1M2_PR $T=197450 17650 0 0 $X=197290 $Y=17490
X1358 99 M1M2_PR $T=197450 27850 0 0 $X=197290 $Y=27690
X1359 30 M1M2_PR $T=201130 12210 0 0 $X=200970 $Y=12050
X1360 123 M1M2_PR $T=201130 14930 0 0 $X=200970 $Y=14770
X1361 123 M1M2_PR $T=201130 15950 0 0 $X=200970 $Y=15790
X1362 31 M1M2_PR $T=201130 17310 0 0 $X=200970 $Y=17150
X1363 98 M1M2_PR $T=201590 2690 0 0 $X=201430 $Y=2530
X1364 98 M1M2_PR $T=201590 10510 0 0 $X=201430 $Y=10350
X1365 29 M1M2_PR $T=201590 13570 0 0 $X=201430 $Y=13410
X1366 29 M1M2_PR $T=201590 25130 0 0 $X=201430 $Y=24970
X1367 131 M1M2_PR $T=204810 11190 0 0 $X=204650 $Y=11030
X1368 123 M1M2_PR $T=204810 14590 0 0 $X=204650 $Y=14430
X1369 123 M1M2_PR $T=204810 15950 0 0 $X=204650 $Y=15790
X1370 132 M1M2_PR $T=204810 17310 0 0 $X=204650 $Y=17150
X1371 123 M1M2_PR $T=205270 11190 0 0 $X=205110 $Y=11030
X1372 102 M1M2_PR $T=205270 14930 0 0 $X=205110 $Y=14770
X1373 102 M1M2_PR $T=205270 29890 0 0 $X=205110 $Y=29730
X1374 33 M1M2_PR $T=208950 13230 0 0 $X=208790 $Y=13070
X1375 104 M1M2_PR $T=212170 17650 0 0 $X=212010 $Y=17490
X1376 104 M1M2_PR $T=212170 25130 0 0 $X=212010 $Y=24970
X1377 134 M1M2_PR $T=212630 17310 0 0 $X=212470 $Y=17150
X1378 119 M1M2_PR $T=216310 16630 0 0 $X=216150 $Y=16470
X1379 35 M1M2_PR $T=219530 17650 0 0 $X=219370 $Y=17490
X1380 123 M1M2_PR $T=219990 14590 0 0 $X=219830 $Y=14430
X1381 123 M1M2_PR $T=219990 16630 0 0 $X=219830 $Y=16470
X1382 108 M1M2_PR $T=223210 15950 0 0 $X=223050 $Y=15790
X1383 108 M1M2_PR $T=223210 22070 0 0 $X=223050 $Y=21910
X1384 37 M1M2_PR $T=225970 58450 0 0 $X=225810 $Y=58290
X1385 37 M1M2_PR $T=225970 60490 0 0 $X=225810 $Y=60330
X1386 36 M1M2_PR $T=227350 12210 0 0 $X=227190 $Y=12050
X1387 123 M1M2_PR $T=230570 11190 0 0 $X=230410 $Y=11030
X1388 123 M1M2_PR $T=230570 14250 0 0 $X=230410 $Y=14090
X1389 123 M1M2_PR $T=230570 16630 0 0 $X=230410 $Y=16470
X1390 135 M1M2_PR $T=231030 11530 0 0 $X=230870 $Y=11370
X1391 32 M1M2_PR $T=231030 17310 0 0 $X=230870 $Y=17150
X1392 136 M1M2_PR $T=234250 16970 0 0 $X=234090 $Y=16810
X1393 110 M1M2_PR $T=237930 6090 0 0 $X=237770 $Y=5930
X1394 110 M1M2_PR $T=237930 10510 0 0 $X=237770 $Y=10350
X1395 38 M1M2_PR $T=239310 19010 0 0 $X=239150 $Y=18850
X1396 137 M1M2_PR $T=245290 14250 0 0 $X=245130 $Y=14090
X1397 123 M1M2_PR $T=245290 14930 0 0 $X=245130 $Y=14770
X1398 123 M1M2_PR $T=245290 15950 0 0 $X=245130 $Y=15790
X1399 38 M1M2_PR $T=245750 14930 0 0 $X=245590 $Y=14770
X1400 38 M1M2_PR $T=245750 19010 0 0 $X=245590 $Y=18850
X1401 11 M1M2_PR $T=248970 6770 0 0 $X=248810 $Y=6610
X1402 11 M1M2_PR $T=248970 7450 0 0 $X=248810 $Y=7290
X1403 40 M1M2_PR $T=248970 14930 0 0 $X=248810 $Y=14770
X1404 34 M1M2_PR $T=253110 12210 0 0 $X=252950 $Y=12050
X1405 1 M1M2_PR $T=255410 7450 0 0 $X=255250 $Y=7290
X1406 112 M1M2_PR $T=256790 14250 0 0 $X=256630 $Y=14090
X1407 138 M1M2_PR $T=260010 11870 0 0 $X=259850 $Y=11710
X1408 123 M1M2_PR $T=260010 14590 0 0 $X=259850 $Y=14430
X1409 123 M1M2_PR $T=260010 15950 0 0 $X=259850 $Y=15790
X1410 139 M1M2_PR $T=260470 13230 0 0 $X=260310 $Y=13070
X1411 40 M1M2_PR $T=260470 13910 0 0 $X=260310 $Y=13750
X1412 40 M1M2_PR $T=260470 14930 0 0 $X=260310 $Y=14770
X1413 114 M1M2_PR $T=263690 4730 0 0 $X=263530 $Y=4570
X1414 114 M1M2_PR $T=263690 13230 0 0 $X=263530 $Y=13070
X1415 123 M1M2_PR $T=264150 11530 0 0 $X=263990 $Y=11370
X1416 123 M1M2_PR $T=264150 14590 0 0 $X=263990 $Y=14430
X1417 44 M1M2_PR $T=269670 8470 0 0 $X=269510 $Y=8310
X1418 43 M1M2_PR $T=272890 35670 0 0 $X=272730 $Y=35510
X1419 140 M1M2_PR $T=278870 13230 0 0 $X=278710 $Y=13070
X1420 42 M1M2_PR $T=282090 13910 0 0 $X=281930 $Y=13750
X1421 46 M1M2_PR $T=283930 9150 0 0 $X=283770 $Y=8990
X1422 45 M1M2_PR $T=286690 650 0 0 $X=286530 $Y=490
X1423 141 M1M2_PR $T=289450 990 0 0 $X=289290 $Y=830
X1424 141 M1M2_PR $T=289450 16630 0 0 $X=289290 $Y=16470
X1425 1 M1M2_PR $T=292670 7450 0 0 $X=292510 $Y=7290
X1426 112 M1M2_PR $T=293130 13910 0 0 $X=292970 $Y=13750
X1427 123 M1M2_PR $T=293130 14590 0 0 $X=292970 $Y=14430
X1428 123 M1M2_PR $T=293130 16630 0 0 $X=292970 $Y=16470
X1429 47 M1M2_PR $T=293130 17650 0 0 $X=292970 $Y=17490
X1430 116 M1M2_PR $T=293590 7790 0 0 $X=293430 $Y=7630
X1431 116 M1M2_PR $T=293590 14930 0 0 $X=293430 $Y=14770
X1432 110 M1M2_PR $T=296350 6090 0 0 $X=296190 $Y=5930
X1433 110 M1M2_PR $T=296810 34990 0 0 $X=296650 $Y=34830
X1434 143 M1M2_PR $T=297270 17650 0 0 $X=297110 $Y=17490
X1435 94 M1M2_PR $T=297270 33630 0 0 $X=297110 $Y=33470
X1436 94 M1M2_PR $T=297270 46550 0 0 $X=297110 $Y=46390
X1437 101 M1M2_PR $T=300490 11190 0 0 $X=300330 $Y=11030
X1438 101 M1M2_PR $T=300490 22750 0 0 $X=300330 $Y=22590
X1439 92 M1M2_PR $T=300490 26490 0 0 $X=300330 $Y=26330
X1440 92 M1M2_PR $T=300490 45870 0 0 $X=300330 $Y=45710
X1441 142 M1M2_PR $T=300950 12210 0 0 $X=300790 $Y=12050
X1442 102 M1M2_PR $T=300950 29890 0 0 $X=300790 $Y=29730
X1443 102 M1M2_PR $T=300950 33630 0 0 $X=300790 $Y=33470
X1444 1 M1M2_PR $T=304170 11530 0 0 $X=304010 $Y=11370
X1445 123 M1M2_PR $T=304170 14590 0 0 $X=304010 $Y=14430
X1446 123 M1M2_PR $T=304170 16630 0 0 $X=304010 $Y=16470
X1447 123 M1M2_PR $T=304630 10850 0 0 $X=304470 $Y=10690
X1448 43 M1M2_PR $T=307850 17310 0 0 $X=307690 $Y=17150
X1449 106 M1M2_PR $T=311530 13570 0 0 $X=311370 $Y=13410
X1450 106 M1M2_PR $T=311530 35670 0 0 $X=311370 $Y=35510
X1451 122 M1M2_PR $T=312450 1670 0 0 $X=312290 $Y=1510
X1452 123 M1M2_PR $T=315210 14930 0 0 $X=315050 $Y=14770
X1453 123 M1M2_PR $T=315210 16630 0 0 $X=315050 $Y=16470
X1454 118 M1M2_PR $T=315210 17650 0 0 $X=315050 $Y=17490
X1455 118 M1M2_PR $T=315210 18670 0 0 $X=315050 $Y=18510
X1456 90 M1M2_PR $T=315210 32950 0 0 $X=315050 $Y=32790
X1457 90 M1M2_PR $T=315210 44510 0 0 $X=315050 $Y=44350
X1458 144 M1M2_PR $T=315670 16630 0 0 $X=315510 $Y=16470
X1459 39 M1M2_PR $T=315670 17650 0 0 $X=315510 $Y=17490
X1460 89 M1M2_PR $T=318890 5410 0 0 $X=318730 $Y=5250
X1461 89 M1M2_PR $T=319350 27510 0 0 $X=319190 $Y=27350
X1462 96 M1M2_PR $T=319350 32270 0 0 $X=319190 $Y=32110
X1463 96 M1M2_PR $T=319350 38050 0 0 $X=319190 $Y=37890
X1464 1 M1M2_PR $T=322570 12210 0 0 $X=322410 $Y=12050
X1465 1 M1M2_PR $T=322570 13230 0 0 $X=322410 $Y=13070
X1466 108 M1M2_PR $T=322570 22070 0 0 $X=322410 $Y=21910
X1467 100 M1M2_PR $T=322570 29550 0 0 $X=322410 $Y=29390
X1468 100 M1M2_PR $T=322570 36690 0 0 $X=322410 $Y=36530
X1469 105 M1M2_PR $T=323030 11870 0 0 $X=322870 $Y=11710
X1470 105 M1M2_PR $T=323490 23770 0 0 $X=323330 $Y=23610
X1471 104 M1M2_PR $T=323490 25470 0 0 $X=323330 $Y=25310
X1472 109 M1M2_PR $T=324410 17650 0 0 $X=324250 $Y=17490
X1473 109 M1M2_PR $T=324410 22750 0 0 $X=324250 $Y=22590
X1474 88 M1M2_PR $T=324410 28530 0 0 $X=324250 $Y=28370
X1475 88 M1M2_PR $T=324410 39410 0 0 $X=324250 $Y=39250
X1476 41 M1M2_PR $T=326250 12210 0 0 $X=326090 $Y=12050
X1477 95 M1M2_PR $T=327170 26150 0 0 $X=327010 $Y=25990
X1478 95 M1M2_PR $T=327170 30910 0 0 $X=327010 $Y=30750
X1479 118 M1M2_PR $T=328090 18670 0 0 $X=327930 $Y=18510
X1480 118 M1M2_PR $T=328090 32610 0 0 $X=327930 $Y=32450
X1481 102 M1M2_PR $T=328090 33630 0 0 $X=327930 $Y=33470
X1482 102 M1M2_PR $T=328090 36690 0 0 $X=327930 $Y=36530
X1483 90 M1M2_PR $T=328090 39920 0 0 $X=327930 $Y=39760
X1484 90 M1M2_PR $T=328090 44510 0 0 $X=327930 $Y=44350
X1485 119 M1M2_PR $T=329010 20030 0 0 $X=328850 $Y=19870
X1486 45 M1M2_PR $T=329470 650 0 0 $X=329310 $Y=490
X1487 117 M1M2_PR $T=329470 16290 0 0 $X=329310 $Y=16130
X1488 117 M1M2_PR $T=329470 20710 0 0 $X=329310 $Y=20550
X1489 92 M1M2_PR $T=329470 40090 0 0 $X=329310 $Y=39930
X1490 92 M1M2_PR $T=329470 45870 0 0 $X=329310 $Y=45710
X1491 123 M1M2_PR $T=329930 10850 0 0 $X=329770 $Y=10690
X1492 123 M1M2_PR $T=329930 14930 0 0 $X=329770 $Y=14770
X1493 93 M1M2_PR $T=329930 27850 0 0 $X=329770 $Y=27690
X1494 93 M1M2_PR $T=329930 28870 0 0 $X=329770 $Y=28710
X1495 145 M1M2_PR $T=330390 11530 0 0 $X=330230 $Y=11370
X1496 94 M1M2_PR $T=330390 40090 0 0 $X=330230 $Y=39930
X1497 94 M1M2_PR $T=330390 46550 0 0 $X=330230 $Y=46390
X1498 98 M1M2_PR $T=331770 2690 0 0 $X=331610 $Y=2530
X1499 98 M1M2_PR $T=332230 37710 0 0 $X=332070 $Y=37550
X1500 107 M1M2_PR $T=332690 27170 0 0 $X=332530 $Y=27010
X1501 107 M1M2_PR $T=333610 10510 0 0 $X=333450 $Y=10350
X1502 112 M1M2_PR $T=333610 14250 0 0 $X=333450 $Y=14090
X1503 112 M1M2_PR $T=333610 33970 0 0 $X=333450 $Y=33810
X1504 97 M1M2_PR $T=334530 3710 0 0 $X=334370 $Y=3550
X1505 97 M1M2_PR $T=334530 25810 0 0 $X=334370 $Y=25650
X1506 114 M1M2_PR $T=335450 4730 0 0 $X=335290 $Y=4570
X1507 114 M1M2_PR $T=335450 33630 0 0 $X=335290 $Y=33470
X1508 103 M1M2_PR $T=335910 24450 0 0 $X=335750 $Y=24290
X1509 103 M1M2_PR $T=336370 16970 0 0 $X=336210 $Y=16810
X1510 104 M1M2_PR $T=336370 36350 0 0 $X=336210 $Y=36190
X1511 46 M1M2_PR $T=337290 9150 0 0 $X=337130 $Y=8990
X1512 46 M1M2_PR $T=337290 11530 0 0 $X=337130 $Y=11370
X1513 108 M1M2_PR $T=338670 40090 0 0 $X=338510 $Y=39930
X1514 11 M1M2_PR $T=339130 6770 0 0 $X=338970 $Y=6610
X1515 11 M1M2_PR $T=339130 28190 0 0 $X=338970 $Y=28030
X1516 111 M1M2_PR $T=340050 22410 0 0 $X=339890 $Y=22250
X1517 111 M1M2_PR $T=340970 10510 0 0 $X=340810 $Y=10350
X1518 115 M1M2_PR $T=341430 12210 0 0 $X=341270 $Y=12050
X1519 115 M1M2_PR $T=341890 21050 0 0 $X=341730 $Y=20890
X1520 116 M1M2_PR $T=342810 7790 0 0 $X=342650 $Y=7630
X1521 113 M1M2_PR $T=343270 22070 0 0 $X=343110 $Y=21910
X1522 116 M1M2_PR $T=343270 33290 0 0 $X=343110 $Y=33130
X1523 113 M1M2_PR $T=344650 12210 0 0 $X=344490 $Y=12050
X1524 146 M1M2_PR $T=348330 12210 0 0 $X=348170 $Y=12050
X1525 44 M1M2_PR $T=348790 11870 0 0 $X=348630 $Y=11710
X1526 44 M1M2_PR $T=349250 8470 0 0 $X=349090 $Y=8310
X1527 147 M1M2_PR $T=352010 11530 0 0 $X=351850 $Y=11370
X1528 2 M1M2_PR $T=379610 9490 0 0 $X=379450 $Y=9330
X1529 11 L1M1_PR $T=37370 11530 0 0 $X=37225 $Y=11415
X1530 10 L1M1_PR $T=38290 11190 0 0 $X=38145 $Y=11075
X1531 11 L1M1_PR $T=45650 30400 0 0 $X=45505 $Y=30285
X1532 4 L1M1_PR $T=53930 52670 0 0 $X=53785 $Y=52555
X1533 5 L1M1_PR $T=54850 51990 0 0 $X=54705 $Y=51875
X1534 6 L1M1_PR $T=55310 24110 0 0 $X=55165 $Y=23995
X1535 7 L1M1_PR $T=56230 24790 0 0 $X=56085 $Y=24675
X1536 85 L1M1_PR $T=65890 23430 0 0 $X=65745 $Y=23315
X1537 123 L1M1_PR $T=91650 16630 0 0 $X=91505 $Y=16515
X1538 148 L1M1_PR $T=92110 17310 0 0 $X=91965 $Y=17195
X1539 14 L1M1_PR $T=93030 16970 0 0 $X=92885 $Y=16855
X1540 119 L1M1_PR $T=94410 15950 0 0 $X=94265 $Y=15835
X1541 7 L1M1_PR $T=95790 24110 0 0 $X=95645 $Y=23995
X1542 5 L1M1_PR $T=96710 24790 0 0 $X=96565 $Y=24675
X1543 5 L1M1_PR $T=98550 24110 0 0 $X=98405 $Y=23995
X1544 8 L1M1_PR $T=99470 24790 0 0 $X=99325 $Y=24675
X1545 9 L1M1_PR $T=100390 25810 0 0 $X=100245 $Y=25695
X1546 7 L1M1_PR $T=101310 24790 0 0 $X=101165 $Y=24675
X1547 123 L1M1_PR $T=114190 14250 0 0 $X=114045 $Y=14135
X1548 123 L1M1_PR $T=114190 16630 0 0 $X=114045 $Y=16515
X1549 149 L1M1_PR $T=114650 13230 0 0 $X=114505 $Y=13115
X1550 150 L1M1_PR $T=114650 17650 0 0 $X=114505 $Y=17535
X1551 16 L1M1_PR $T=115230 14250 0 0 $X=115085 $Y=14135
X1552 13 L1M1_PR $T=115570 17310 0 0 $X=115425 $Y=17195
X1553 91 L1M1_PR $T=116950 14930 0 0 $X=116805 $Y=14815
X1554 89 L1M1_PR $T=116950 15950 0 0 $X=116805 $Y=15835
X1555 123 L1M1_PR $T=118790 16630 0 0 $X=118645 $Y=16515
X1556 151 L1M1_PR $T=119250 17650 0 0 $X=119105 $Y=17535
X1557 18 L1M1_PR $T=120170 17310 0 0 $X=120025 $Y=17195
X1558 93 L1M1_PR $T=121550 16290 0 0 $X=121405 $Y=16175
X1559 88 L1M1_PR $T=124770 16290 0 0 $X=124625 $Y=16175
X1560 15 L1M1_PR $T=126140 17310 0 0 $X=125995 $Y=17195
X1561 152 L1M1_PR $T=127070 17310 0 0 $X=126925 $Y=17195
X1562 123 L1M1_PR $T=127530 16630 0 0 $X=127385 $Y=16515
X1563 90 L1M1_PR $T=128910 15950 0 0 $X=128765 $Y=15835
X1564 17 L1M1_PR $T=130290 17310 0 0 $X=130145 $Y=17195
X1565 153 L1M1_PR $T=131210 17310 0 0 $X=131065 $Y=17195
X1566 123 L1M1_PR $T=131670 16630 0 0 $X=131525 $Y=16515
X1567 123 L1M1_PR $T=137650 14250 0 0 $X=137505 $Y=14135
X1568 154 L1M1_PR $T=138110 13230 0 0 $X=137965 $Y=13115
X1569 19 L1M1_PR $T=139030 13910 0 0 $X=138885 $Y=13795
X1570 92 L1M1_PR $T=140410 14930 0 0 $X=140265 $Y=14815
X1571 123 L1M1_PR $T=141790 11190 0 0 $X=141645 $Y=11075
X1572 124 L1M1_PR $T=142710 11530 0 0 $X=142565 $Y=11415
X1573 21 L1M1_PR $T=143170 11870 0 0 $X=143025 $Y=11755
X1574 94 L1M1_PR $T=145010 10850 0 0 $X=144865 $Y=10735
X1575 123 L1M1_PR $T=152370 16630 0 0 $X=152225 $Y=16515
X1576 155 L1M1_PR $T=152830 17650 0 0 $X=152685 $Y=17535
X1577 22 L1M1_PR $T=153290 16630 0 0 $X=153145 $Y=16515
X1578 95 L1M1_PR $T=155130 15950 0 0 $X=154985 $Y=15835
X1579 123 L1M1_PR $T=167090 16630 0 0 $X=166945 $Y=16515
X1580 125 L1M1_PR $T=168010 17310 0 0 $X=167865 $Y=17195
X1581 24 L1M1_PR $T=168470 17650 0 0 $X=168325 $Y=17535
X1582 97 L1M1_PR $T=170220 15950 0 0 $X=170075 $Y=15835
X1583 123 L1M1_PR $T=171690 14250 0 0 $X=171545 $Y=14135
X1584 126 L1M1_PR $T=172600 13570 0 0 $X=172455 $Y=13455
X1585 23 L1M1_PR $T=173070 13910 0 0 $X=172925 $Y=13795
X1586 127 L1M1_PR $T=173530 11870 0 0 $X=173385 $Y=11755
X1587 25 L1M1_PR $T=173990 12210 0 0 $X=173845 $Y=12095
X1588 96 L1M1_PR $T=174910 14930 0 0 $X=174765 $Y=14815
X1589 123 L1M1_PR $T=175120 11530 0 0 $X=174975 $Y=11415
X1590 98 L1M1_PR $T=175830 10510 0 0 $X=175685 $Y=10395
X1591 100 L1M1_PR $T=178590 17650 0 0 $X=178445 $Y=17535
X1592 28 L1M1_PR $T=180430 17650 0 0 $X=180285 $Y=17535
X1593 128 L1M1_PR $T=180880 17310 0 0 $X=180735 $Y=17195
X1594 123 L1M1_PR $T=181810 16630 0 0 $X=181665 $Y=16515
X1595 123 L1M1_PR $T=183775 15950 0 0 $X=183630 $Y=15835
X1596 129 L1M1_PR $T=184110 17310 0 0 $X=183965 $Y=17195
X1597 26 L1M1_PR $T=184570 17310 0 0 $X=184425 $Y=17195
X1598 99 L1M1_PR $T=186410 17650 0 0 $X=186265 $Y=17535
X1599 123 L1M1_PR $T=200835 14930 0 0 $X=200690 $Y=14815
X1600 130 L1M1_PR $T=201130 13230 0 0 $X=200985 $Y=13115
X1601 29 L1M1_PR $T=201590 13570 0 0 $X=201445 $Y=13455
X1602 101 L1M1_PR $T=202050 10850 0 0 $X=201905 $Y=10735
X1603 104 L1M1_PR $T=202050 17650 0 0 $X=201905 $Y=17535
X1604 102 L1M1_PR $T=203430 14930 0 0 $X=203285 $Y=14815
X1605 30 L1M1_PR $T=203890 12210 0 0 $X=203745 $Y=12095
X1606 31 L1M1_PR $T=203890 17310 0 0 $X=203745 $Y=17195
X1607 131 L1M1_PR $T=204350 11190 0 0 $X=204205 $Y=11075
X1608 132 L1M1_PR $T=204350 17310 0 0 $X=204205 $Y=17195
X1609 123 L1M1_PR $T=204810 16630 0 0 $X=204665 $Y=16515
X1610 123 L1M1_PR $T=205270 11190 0 0 $X=205125 $Y=11075
X1611 123 L1M1_PR $T=207570 14250 0 0 $X=207425 $Y=14135
X1612 133 L1M1_PR $T=208490 13910 0 0 $X=208345 $Y=13795
X1613 33 L1M1_PR $T=208950 13230 0 0 $X=208805 $Y=13115
X1614 106 L1M1_PR $T=210790 13230 0 0 $X=210645 $Y=13115
X1615 108 L1M1_PR $T=216770 15950 0 0 $X=216625 $Y=15835
X1616 35 L1M1_PR $T=218610 17650 0 0 $X=218465 $Y=17535
X1617 134 L1M1_PR $T=219070 16970 0 0 $X=218925 $Y=16855
X1618 123 L1M1_PR $T=219990 16630 0 0 $X=219845 $Y=16515
X1619 123 L1M1_PR $T=230570 11190 0 0 $X=230425 $Y=11075
X1620 103 L1M1_PR $T=230570 17650 0 0 $X=230425 $Y=17535
X1621 135 L1M1_PR $T=231490 11530 0 0 $X=231345 $Y=11415
X1622 36 L1M1_PR $T=231950 12210 0 0 $X=231805 $Y=12095
X1623 32 L1M1_PR $T=232410 17310 0 0 $X=232265 $Y=17195
X1624 136 L1M1_PR $T=232870 16970 0 0 $X=232725 $Y=16855
X1625 123 L1M1_PR $T=233330 16630 0 0 $X=233185 $Y=16515
X1626 110 L1M1_PR $T=233790 10510 0 0 $X=233645 $Y=10395
X1627 123 L1M1_PR $T=244830 14250 0 0 $X=244685 $Y=14135
X1628 137 L1M1_PR $T=245750 14250 0 0 $X=245605 $Y=14135
X1629 38 L1M1_PR $T=246160 13910 0 0 $X=246015 $Y=13795
X1630 112 L1M1_PR $T=248050 14590 0 0 $X=247905 $Y=14475
X1631 123 L1M1_PR $T=259550 14250 0 0 $X=259405 $Y=14135
X1632 123 L1M1_PR $T=260010 11190 0 0 $X=259865 $Y=11075
X1633 138 L1M1_PR $T=260470 11870 0 0 $X=260325 $Y=11755
X1634 139 L1M1_PR $T=260470 13230 0 0 $X=260325 $Y=13115
X1635 34 L1M1_PR $T=260930 12210 0 0 $X=260785 $Y=12095
X1636 40 L1M1_PR $T=260930 13910 0 0 $X=260785 $Y=13795
X1637 105 L1M1_PR $T=262770 12210 0 0 $X=262625 $Y=12095
X1638 114 L1M1_PR $T=262770 13230 0 0 $X=262625 $Y=13115
X1639 43 L1M1_PR $T=272640 35670 0 0 $X=272495 $Y=35555
X1640 123 L1M1_PR $T=281170 14250 0 0 $X=281025 $Y=14135
X1641 140 L1M1_PR $T=281630 13230 0 0 $X=281485 $Y=13115
X1642 42 L1M1_PR $T=282090 13910 0 0 $X=281945 $Y=13795
X1643 116 L1M1_PR $T=283930 14930 0 0 $X=283785 $Y=14815
X1644 117 L1M1_PR $T=290370 16290 0 0 $X=290225 $Y=16175
X1645 47 L1M1_PR $T=292210 17650 0 0 $X=292065 $Y=17535
X1646 141 L1M1_PR $T=292670 16630 0 0 $X=292525 $Y=16515
X1647 123 L1M1_PR $T=293130 16630 0 0 $X=292985 $Y=16515
X1648 123 L1M1_PR $T=303710 11190 0 0 $X=303565 $Y=11075
X1649 123 L1M1_PR $T=304170 16630 0 0 $X=304025 $Y=16515
X1650 142 L1M1_PR $T=304630 12210 0 0 $X=304485 $Y=12095
X1651 143 L1M1_PR $T=304630 17650 0 0 $X=304485 $Y=17535
X1652 1 L1M1_PR $T=305090 11530 0 0 $X=304945 $Y=11415
X1653 43 L1M1_PR $T=305090 17310 0 0 $X=304945 $Y=17195
X1654 107 L1M1_PR $T=306930 10510 0 0 $X=306785 $Y=10395
X1655 118 L1M1_PR $T=306930 17650 0 0 $X=306785 $Y=17535
X1656 123 L1M1_PR $T=314750 16630 0 0 $X=314605 $Y=16515
X1657 144 L1M1_PR $T=315670 16630 0 0 $X=315525 $Y=16515
X1658 39 L1M1_PR $T=316130 17650 0 0 $X=315985 $Y=17535
X1659 109 L1M1_PR $T=317970 17650 0 0 $X=317825 $Y=17535
X1660 123 L1M1_PR $T=331310 11190 0 0 $X=331165 $Y=11075
X1661 145 L1M1_PR $T=332230 11530 0 0 $X=332085 $Y=11415
X1662 41 L1M1_PR $T=332690 12210 0 0 $X=332545 $Y=12095
X1663 111 L1M1_PR $T=334530 10510 0 0 $X=334385 $Y=10395
X1664 11 L1M1_PR $T=338210 28190 0 0 $X=338065 $Y=28075
X1665 115 L1M1_PR $T=341890 12210 0 0 $X=341745 $Y=12095
X1666 46 L1M1_PR $T=343730 11530 0 0 $X=343585 $Y=11415
X1667 146 L1M1_PR $T=344190 11870 0 0 $X=344045 $Y=11755
X1668 123 L1M1_PR $T=344650 11190 0 0 $X=344505 $Y=11075
X1669 113 L1M1_PR $T=346030 12210 0 0 $X=345885 $Y=12095
X1670 44 L1M1_PR $T=347870 11870 0 0 $X=347725 $Y=11755
X1671 147 L1M1_PR $T=348330 11530 0 0 $X=348185 $Y=11415
X1672 123 L1M1_PR $T=348790 11190 0 0 $X=348645 $Y=11075
X1673 1 L1M1_PR $T=352470 13570 0 0 $X=352325 $Y=13455
X1674 10 M3M4_PR $T=10230 2240 0 0 $X=10040 $Y=2075
X1675 123 M3M4_PR $T=35070 1020 0 0 $X=34880 $Y=855
X1676 150 M3M4_PR $T=59910 8950 0 0 $X=59720 $Y=8785
X1677 149 M3M4_PR $T=84060 2240 0 0 $X=83870 $Y=2075
X1678 8 M3M4_PR $T=105450 1020 0 0 $X=105260 $Y=855
X1679 8 M3M4_PR $T=106140 1020 0 0 $X=105950 $Y=855
X1680 151 M3M4_PR $T=108900 4680 0 0 $X=108710 $Y=4515
X1681 8 M3M4_PR $T=116490 1020 0 0 $X=116300 $Y=855
X1682 8 M3M4_PR $T=117180 1020 0 0 $X=116990 $Y=855
X1683 155 M3M4_PR $T=133740 2850 0 0 $X=133550 $Y=2685
X1684 22 M3M4_PR $T=153750 18710 0 0 $X=153560 $Y=18545
X1685 125 M3M4_PR $T=157890 2240 0 0 $X=157700 $Y=2075
X1686 9 M3M4_PR $T=170310 43720 0 0 $X=170120 $Y=43555
X1687 9 M3M4_PR $T=170310 47380 0 0 $X=170120 $Y=47215
X1688 129 M3M4_PR $T=182730 4680 0 0 $X=182540 $Y=4515
X1689 30 M3M4_PR $T=193080 14440 0 0 $X=192890 $Y=14275
X1690 131 M3M4_PR $T=207570 2240 0 0 $X=207380 $Y=2075
X1691 34 M3M4_PR $T=219990 22370 0 0 $X=219800 $Y=22205
X1692 1 M3M4_PR $T=230340 7730 0 0 $X=230150 $Y=7565
X1693 136 M3M4_PR $T=232410 8950 0 0 $X=232220 $Y=8785
X1694 1 M3M4_PR $T=235170 7730 0 0 $X=234980 $Y=7565
X1695 1 M3M4_PR $T=235860 7730 0 0 $X=235670 $Y=7565
X1696 34 M3M4_PR $T=236550 22370 0 0 $X=236360 $Y=22205
X1697 34 M3M4_PR $T=237240 22370 0 0 $X=237050 $Y=22205
X1698 1 M3M4_PR $T=247590 7730 0 0 $X=247400 $Y=7565
X1699 34 M3M4_PR $T=247590 22370 0 0 $X=247400 $Y=22205
X1700 1 M3M4_PR $T=248280 7730 0 0 $X=248090 $Y=7565
X1701 34 M3M4_PR $T=248280 22370 0 0 $X=248090 $Y=22205
X1702 138 M3M4_PR $T=256560 2240 0 0 $X=256370 $Y=2075
X1703 41 M3M4_PR $T=257940 9560 0 0 $X=257750 $Y=9395
X1704 142 M3M4_PR $T=281400 2850 0 0 $X=281210 $Y=2685
X1705 43 M3M4_PR $T=291750 34570 0 0 $X=291560 $Y=34405
X1706 43 M3M4_PR $T=292440 34570 0 0 $X=292250 $Y=34405
X1707 39 M3M4_PR $T=297270 27250 0 0 $X=297080 $Y=27085
X1708 39 M3M4_PR $T=297960 27250 0 0 $X=297770 $Y=27085
X1709 43 M3M4_PR $T=302790 34570 0 0 $X=302600 $Y=34405
X1710 43 M3M4_PR $T=303480 34570 0 0 $X=303290 $Y=34405
X1711 144 M3M4_PR $T=305550 2240 0 0 $X=305360 $Y=2075
X1712 39 M3M4_PR $T=308310 27250 0 0 $X=308120 $Y=27085
X1713 39 M3M4_PR $T=309000 27250 0 0 $X=308810 $Y=27085
X1714 41 M3M4_PR $T=311070 8950 0 0 $X=310880 $Y=8785
X1715 41 M3M4_PR $T=311760 8950 0 0 $X=311570 $Y=8785
X1716 41 M3M4_PR $T=324180 9560 0 0 $X=323990 $Y=9395
X1717 41 M3M4_PR $T=324870 9560 0 0 $X=324680 $Y=9395
X1718 145 M3M4_PR $T=330390 10780 0 0 $X=330200 $Y=10615
X1719 146 M3M4_PR $T=352470 1020 0 0 $X=352280 $Y=855
X1720 146 M3M4_PR $T=353160 1020 0 0 $X=352970 $Y=855
X1721 147 M3M4_PR $T=355230 2850 0 0 $X=355040 $Y=2685
X1722 146 M3M4_PR $T=364890 1020 0 0 $X=364700 $Y=855
X1723 146 M3M4_PR $T=365580 1020 0 0 $X=365390 $Y=855
X1724 146 M3M4_PR $T=379380 1020 0 0 $X=379190 $Y=855
X1725 2 digital_ldo_top_VIA0 $T=12530 10110 0 0 $X=12280 $Y=9980
X1726 2 digital_ldo_top_VIA0 $T=16210 10110 0 0 $X=15960 $Y=9980
X1727 2 digital_ldo_top_VIA0 $T=19890 10110 0 0 $X=19640 $Y=9980
X1728 2 digital_ldo_top_VIA0 $T=23570 10110 0 0 $X=23320 $Y=9980
X1729 2 digital_ldo_top_VIA0 $T=27250 10110 0 0 $X=27000 $Y=9980
X1730 2 digital_ldo_top_VIA0 $T=30930 10110 0 0 $X=30680 $Y=9980
X1731 2 digital_ldo_top_VIA0 $T=34610 10110 0 0 $X=34360 $Y=9980
X1732 2 digital_ldo_top_VIA0 $T=38290 10110 0 0 $X=38040 $Y=9980
X1733 2 digital_ldo_top_VIA0 $T=41970 10110 0 0 $X=41720 $Y=9980
X1734 2 digital_ldo_top_VIA0 $T=45650 10110 0 0 $X=45400 $Y=9980
X1735 2 digital_ldo_top_VIA0 $T=49330 10110 0 0 $X=49080 $Y=9980
X1736 2 digital_ldo_top_VIA0 $T=53010 10110 0 0 $X=52760 $Y=9980
X1737 2 digital_ldo_top_VIA0 $T=56690 10110 0 0 $X=56440 $Y=9980
X1738 2 digital_ldo_top_VIA0 $T=60370 10110 0 0 $X=60120 $Y=9980
X1739 2 digital_ldo_top_VIA0 $T=64050 10110 0 0 $X=63800 $Y=9980
X1740 2 digital_ldo_top_VIA0 $T=67730 10110 0 0 $X=67480 $Y=9980
X1741 2 digital_ldo_top_VIA0 $T=71410 10110 0 0 $X=71160 $Y=9980
X1742 2 digital_ldo_top_VIA0 $T=75090 10110 0 0 $X=74840 $Y=9980
X1743 2 digital_ldo_top_VIA0 $T=78770 10110 0 0 $X=78520 $Y=9980
X1744 2 digital_ldo_top_VIA0 $T=82450 10110 0 0 $X=82200 $Y=9980
X1745 2 digital_ldo_top_VIA0 $T=86130 10110 0 0 $X=85880 $Y=9980
X1746 2 digital_ldo_top_VIA0 $T=89810 10110 0 0 $X=89560 $Y=9980
X1747 2 digital_ldo_top_VIA0 $T=93490 10110 0 0 $X=93240 $Y=9980
X1748 2 digital_ldo_top_VIA0 $T=97170 10110 0 0 $X=96920 $Y=9980
X1749 2 digital_ldo_top_VIA0 $T=100850 10110 0 0 $X=100600 $Y=9980
X1750 2 digital_ldo_top_VIA0 $T=104530 10110 0 0 $X=104280 $Y=9980
X1751 2 digital_ldo_top_VIA0 $T=108210 10110 0 0 $X=107960 $Y=9980
X1752 2 digital_ldo_top_VIA0 $T=111890 10110 0 0 $X=111640 $Y=9980
X1753 2 digital_ldo_top_VIA0 $T=115570 10110 0 0 $X=115320 $Y=9980
X1754 2 digital_ldo_top_VIA0 $T=119250 10110 0 0 $X=119000 $Y=9980
X1755 2 digital_ldo_top_VIA0 $T=122930 10110 0 0 $X=122680 $Y=9980
X1756 2 digital_ldo_top_VIA0 $T=126610 10110 0 0 $X=126360 $Y=9980
X1757 2 digital_ldo_top_VIA0 $T=130290 10110 0 0 $X=130040 $Y=9980
X1758 2 digital_ldo_top_VIA0 $T=133970 10110 0 0 $X=133720 $Y=9980
X1759 2 digital_ldo_top_VIA0 $T=137650 10110 0 0 $X=137400 $Y=9980
X1760 2 digital_ldo_top_VIA0 $T=141330 10110 0 0 $X=141080 $Y=9980
X1761 2 digital_ldo_top_VIA0 $T=145010 10110 0 0 $X=144760 $Y=9980
X1762 2 digital_ldo_top_VIA0 $T=148690 10110 0 0 $X=148440 $Y=9980
X1763 2 digital_ldo_top_VIA0 $T=152370 10110 0 0 $X=152120 $Y=9980
X1764 2 digital_ldo_top_VIA0 $T=156050 10110 0 0 $X=155800 $Y=9980
X1765 2 digital_ldo_top_VIA0 $T=159730 10110 0 0 $X=159480 $Y=9980
X1766 2 digital_ldo_top_VIA0 $T=163410 10110 0 0 $X=163160 $Y=9980
X1767 2 digital_ldo_top_VIA0 $T=167090 10110 0 0 $X=166840 $Y=9980
X1768 2 digital_ldo_top_VIA0 $T=170770 10110 0 0 $X=170520 $Y=9980
X1769 2 digital_ldo_top_VIA0 $T=174450 10110 0 0 $X=174200 $Y=9980
X1770 2 digital_ldo_top_VIA0 $T=178130 10110 0 0 $X=177880 $Y=9980
X1771 2 digital_ldo_top_VIA0 $T=181810 10110 0 0 $X=181560 $Y=9980
X1772 2 digital_ldo_top_VIA0 $T=185490 10110 0 0 $X=185240 $Y=9980
X1773 2 digital_ldo_top_VIA0 $T=189170 10110 0 0 $X=188920 $Y=9980
X1774 2 digital_ldo_top_VIA0 $T=192850 10110 0 0 $X=192600 $Y=9980
X1775 2 digital_ldo_top_VIA0 $T=196530 10110 0 0 $X=196280 $Y=9980
X1776 2 digital_ldo_top_VIA0 $T=200210 10110 0 0 $X=199960 $Y=9980
X1777 2 digital_ldo_top_VIA0 $T=203890 10110 0 0 $X=203640 $Y=9980
X1778 2 digital_ldo_top_VIA0 $T=207570 10110 0 0 $X=207320 $Y=9980
X1779 2 digital_ldo_top_VIA0 $T=211250 10110 0 0 $X=211000 $Y=9980
X1780 2 digital_ldo_top_VIA0 $T=214930 10110 0 0 $X=214680 $Y=9980
X1781 2 digital_ldo_top_VIA0 $T=218610 10110 0 0 $X=218360 $Y=9980
X1782 2 digital_ldo_top_VIA0 $T=222290 10110 0 0 $X=222040 $Y=9980
X1783 2 digital_ldo_top_VIA0 $T=225970 10110 0 0 $X=225720 $Y=9980
X1784 2 digital_ldo_top_VIA0 $T=229650 10110 0 0 $X=229400 $Y=9980
X1785 2 digital_ldo_top_VIA0 $T=233330 10110 0 0 $X=233080 $Y=9980
X1786 2 digital_ldo_top_VIA0 $T=237010 10110 0 0 $X=236760 $Y=9980
X1787 2 digital_ldo_top_VIA0 $T=240690 10110 0 0 $X=240440 $Y=9980
X1788 2 digital_ldo_top_VIA0 $T=244370 10110 0 0 $X=244120 $Y=9980
X1789 2 digital_ldo_top_VIA0 $T=248050 10110 0 0 $X=247800 $Y=9980
X1790 2 digital_ldo_top_VIA0 $T=251730 10110 0 0 $X=251480 $Y=9980
X1791 2 digital_ldo_top_VIA0 $T=255410 10110 0 0 $X=255160 $Y=9980
X1792 2 digital_ldo_top_VIA0 $T=259090 10110 0 0 $X=258840 $Y=9980
X1793 2 digital_ldo_top_VIA0 $T=262770 10110 0 0 $X=262520 $Y=9980
X1794 2 digital_ldo_top_VIA0 $T=266450 10110 0 0 $X=266200 $Y=9980
X1795 2 digital_ldo_top_VIA0 $T=270130 10110 0 0 $X=269880 $Y=9980
X1796 2 digital_ldo_top_VIA0 $T=273810 10110 0 0 $X=273560 $Y=9980
X1797 2 digital_ldo_top_VIA0 $T=277490 10110 0 0 $X=277240 $Y=9980
X1798 2 digital_ldo_top_VIA0 $T=281170 10110 0 0 $X=280920 $Y=9980
X1799 2 digital_ldo_top_VIA0 $T=284850 10110 0 0 $X=284600 $Y=9980
X1800 2 digital_ldo_top_VIA0 $T=288530 10110 0 0 $X=288280 $Y=9980
X1801 2 digital_ldo_top_VIA0 $T=292210 10110 0 0 $X=291960 $Y=9980
X1802 2 digital_ldo_top_VIA0 $T=295890 10110 0 0 $X=295640 $Y=9980
X1803 2 digital_ldo_top_VIA0 $T=299570 10110 0 0 $X=299320 $Y=9980
X1804 2 digital_ldo_top_VIA0 $T=303250 10110 0 0 $X=303000 $Y=9980
X1805 2 digital_ldo_top_VIA0 $T=306930 10110 0 0 $X=306680 $Y=9980
X1806 2 digital_ldo_top_VIA0 $T=310610 10110 0 0 $X=310360 $Y=9980
X1807 2 digital_ldo_top_VIA0 $T=314290 10110 0 0 $X=314040 $Y=9980
X1808 2 digital_ldo_top_VIA0 $T=317970 10110 0 0 $X=317720 $Y=9980
X1809 2 digital_ldo_top_VIA0 $T=321650 10110 0 0 $X=321400 $Y=9980
X1810 2 digital_ldo_top_VIA0 $T=325330 10110 0 0 $X=325080 $Y=9980
X1811 2 digital_ldo_top_VIA0 $T=329010 10110 0 0 $X=328760 $Y=9980
X1812 2 digital_ldo_top_VIA0 $T=332690 10110 0 0 $X=332440 $Y=9980
X1813 2 digital_ldo_top_VIA0 $T=336370 10110 0 0 $X=336120 $Y=9980
X1814 2 digital_ldo_top_VIA0 $T=340050 10110 0 0 $X=339800 $Y=9980
X1815 2 digital_ldo_top_VIA0 $T=343730 10110 0 0 $X=343480 $Y=9980
X1816 2 digital_ldo_top_VIA0 $T=347410 10110 0 0 $X=347160 $Y=9980
X1817 2 digital_ldo_top_VIA0 $T=351090 10110 0 0 $X=350840 $Y=9980
X1818 2 digital_ldo_top_VIA0 $T=354770 10110 0 0 $X=354520 $Y=9980
X1819 2 digital_ldo_top_VIA0 $T=358450 10110 0 0 $X=358200 $Y=9980
X1820 2 digital_ldo_top_VIA0 $T=362130 10110 0 0 $X=361880 $Y=9980
X1821 2 digital_ldo_top_VIA0 $T=365810 10110 0 0 $X=365560 $Y=9980
X1822 2 digital_ldo_top_VIA0 $T=369490 10110 0 0 $X=369240 $Y=9980
X1823 2 digital_ldo_top_VIA0 $T=373170 10110 0 0 $X=372920 $Y=9980
X1824 2 digital_ldo_top_VIA0 $T=376850 10110 0 0 $X=376600 $Y=9980
X1825 3 digital_ldo_top_VIA1 $T=11150 12720 0 0 $X=10900 $Y=12480
X1826 3 digital_ldo_top_VIA1 $T=11150 18160 0 0 $X=10900 $Y=17920
X1827 3 digital_ldo_top_VIA1 $T=11150 23600 0 0 $X=10900 $Y=23360
X1828 3 digital_ldo_top_VIA1 $T=11150 29040 0 0 $X=10900 $Y=28800
X1829 3 digital_ldo_top_VIA1 $T=11150 34480 0 0 $X=10900 $Y=34240
X1830 3 digital_ldo_top_VIA1 $T=11150 39920 0 0 $X=10900 $Y=39680
X1831 3 digital_ldo_top_VIA1 $T=11150 45360 0 0 $X=10900 $Y=45120
X1832 3 digital_ldo_top_VIA1 $T=11150 50800 0 0 $X=10900 $Y=50560
X1833 3 digital_ldo_top_VIA1 $T=11150 56240 0 0 $X=10900 $Y=56000
X1834 3 digital_ldo_top_VIA1 $T=11150 61680 0 0 $X=10900 $Y=61440
X1835 3 digital_ldo_top_VIA1 $T=11150 67120 0 0 $X=10900 $Y=66880
X1836 3 digital_ldo_top_VIA1 $T=11150 72560 0 0 $X=10900 $Y=72320
X1837 3 digital_ldo_top_VIA1 $T=11150 78000 0 0 $X=10900 $Y=77760
X1838 3 digital_ldo_top_VIA1 $T=11150 83440 0 0 $X=10900 $Y=83200
X1839 3 digital_ldo_top_VIA1 $T=11150 88880 0 0 $X=10900 $Y=88640
X1840 3 digital_ldo_top_VIA1 $T=11150 94320 0 0 $X=10900 $Y=94080
X1841 3 digital_ldo_top_VIA1 $T=11150 99760 0 0 $X=10900 $Y=99520
X1842 3 digital_ldo_top_VIA1 $T=11150 105200 0 0 $X=10900 $Y=104960
X1843 3 digital_ldo_top_VIA1 $T=11150 110640 0 0 $X=10900 $Y=110400
X1844 3 digital_ldo_top_VIA1 $T=11150 116080 0 0 $X=10900 $Y=115840
X1845 3 digital_ldo_top_VIA1 $T=11150 121520 0 0 $X=10900 $Y=121280
X1846 3 digital_ldo_top_VIA1 $T=11150 126960 0 0 $X=10900 $Y=126720
X1847 2 digital_ldo_top_VIA1 $T=12530 15440 0 0 $X=12280 $Y=15200
X1848 2 digital_ldo_top_VIA1 $T=12530 20880 0 0 $X=12280 $Y=20640
X1849 2 digital_ldo_top_VIA1 $T=12530 26320 0 0 $X=12280 $Y=26080
X1850 2 digital_ldo_top_VIA1 $T=12530 31760 0 0 $X=12280 $Y=31520
X1851 2 digital_ldo_top_VIA1 $T=12530 37200 0 0 $X=12280 $Y=36960
X1852 2 digital_ldo_top_VIA1 $T=12530 42640 0 0 $X=12280 $Y=42400
X1853 2 digital_ldo_top_VIA1 $T=12530 48080 0 0 $X=12280 $Y=47840
X1854 2 digital_ldo_top_VIA1 $T=12530 53520 0 0 $X=12280 $Y=53280
X1855 2 digital_ldo_top_VIA1 $T=12530 58960 0 0 $X=12280 $Y=58720
X1856 2 digital_ldo_top_VIA1 $T=12530 64400 0 0 $X=12280 $Y=64160
X1857 2 digital_ldo_top_VIA1 $T=12530 69840 0 0 $X=12280 $Y=69600
X1858 2 digital_ldo_top_VIA1 $T=12530 75280 0 0 $X=12280 $Y=75040
X1859 2 digital_ldo_top_VIA1 $T=12530 80720 0 0 $X=12280 $Y=80480
X1860 2 digital_ldo_top_VIA1 $T=12530 86160 0 0 $X=12280 $Y=85920
X1861 2 digital_ldo_top_VIA1 $T=12530 91600 0 0 $X=12280 $Y=91360
X1862 2 digital_ldo_top_VIA1 $T=12530 97040 0 0 $X=12280 $Y=96800
X1863 2 digital_ldo_top_VIA1 $T=12530 102480 0 0 $X=12280 $Y=102240
X1864 2 digital_ldo_top_VIA1 $T=12530 107920 0 0 $X=12280 $Y=107680
X1865 2 digital_ldo_top_VIA1 $T=12530 113360 0 0 $X=12280 $Y=113120
X1866 2 digital_ldo_top_VIA1 $T=12530 118800 0 0 $X=12280 $Y=118560
X1867 2 digital_ldo_top_VIA1 $T=12530 124240 0 0 $X=12280 $Y=124000
X1868 2 digital_ldo_top_VIA1 $T=12530 129680 0 0 $X=12280 $Y=129440
X1869 3 digital_ldo_top_VIA1 $T=14830 12720 0 0 $X=14580 $Y=12480
X1870 3 digital_ldo_top_VIA1 $T=14830 18160 0 0 $X=14580 $Y=17920
X1871 3 digital_ldo_top_VIA1 $T=14830 23600 0 0 $X=14580 $Y=23360
X1872 3 digital_ldo_top_VIA1 $T=14830 29040 0 0 $X=14580 $Y=28800
X1873 3 digital_ldo_top_VIA1 $T=14830 34480 0 0 $X=14580 $Y=34240
X1874 3 digital_ldo_top_VIA1 $T=14830 39920 0 0 $X=14580 $Y=39680
X1875 3 digital_ldo_top_VIA1 $T=14830 45360 0 0 $X=14580 $Y=45120
X1876 3 digital_ldo_top_VIA1 $T=14830 50800 0 0 $X=14580 $Y=50560
X1877 3 digital_ldo_top_VIA1 $T=14830 56240 0 0 $X=14580 $Y=56000
X1878 3 digital_ldo_top_VIA1 $T=14830 61680 0 0 $X=14580 $Y=61440
X1879 3 digital_ldo_top_VIA1 $T=14830 67120 0 0 $X=14580 $Y=66880
X1880 3 digital_ldo_top_VIA1 $T=14830 72560 0 0 $X=14580 $Y=72320
X1881 3 digital_ldo_top_VIA1 $T=14830 78000 0 0 $X=14580 $Y=77760
X1882 3 digital_ldo_top_VIA1 $T=14830 83440 0 0 $X=14580 $Y=83200
X1883 3 digital_ldo_top_VIA1 $T=14830 88880 0 0 $X=14580 $Y=88640
X1884 3 digital_ldo_top_VIA1 $T=14830 94320 0 0 $X=14580 $Y=94080
X1885 3 digital_ldo_top_VIA1 $T=14830 99760 0 0 $X=14580 $Y=99520
X1886 3 digital_ldo_top_VIA1 $T=14830 105200 0 0 $X=14580 $Y=104960
X1887 3 digital_ldo_top_VIA1 $T=14830 110640 0 0 $X=14580 $Y=110400
X1888 3 digital_ldo_top_VIA1 $T=14830 116080 0 0 $X=14580 $Y=115840
X1889 3 digital_ldo_top_VIA1 $T=14830 121520 0 0 $X=14580 $Y=121280
X1890 3 digital_ldo_top_VIA1 $T=14830 126960 0 0 $X=14580 $Y=126720
X1891 2 digital_ldo_top_VIA1 $T=16210 15440 0 0 $X=15960 $Y=15200
X1892 2 digital_ldo_top_VIA1 $T=16210 20880 0 0 $X=15960 $Y=20640
X1893 2 digital_ldo_top_VIA1 $T=16210 26320 0 0 $X=15960 $Y=26080
X1894 2 digital_ldo_top_VIA1 $T=16210 31760 0 0 $X=15960 $Y=31520
X1895 2 digital_ldo_top_VIA1 $T=16210 37200 0 0 $X=15960 $Y=36960
X1896 2 digital_ldo_top_VIA1 $T=16210 42640 0 0 $X=15960 $Y=42400
X1897 2 digital_ldo_top_VIA1 $T=16210 48080 0 0 $X=15960 $Y=47840
X1898 2 digital_ldo_top_VIA1 $T=16210 53520 0 0 $X=15960 $Y=53280
X1899 2 digital_ldo_top_VIA1 $T=16210 58960 0 0 $X=15960 $Y=58720
X1900 2 digital_ldo_top_VIA1 $T=16210 64400 0 0 $X=15960 $Y=64160
X1901 2 digital_ldo_top_VIA1 $T=16210 69840 0 0 $X=15960 $Y=69600
X1902 2 digital_ldo_top_VIA1 $T=16210 75280 0 0 $X=15960 $Y=75040
X1903 2 digital_ldo_top_VIA1 $T=16210 80720 0 0 $X=15960 $Y=80480
X1904 2 digital_ldo_top_VIA1 $T=16210 86160 0 0 $X=15960 $Y=85920
X1905 2 digital_ldo_top_VIA1 $T=16210 91600 0 0 $X=15960 $Y=91360
X1906 2 digital_ldo_top_VIA1 $T=16210 97040 0 0 $X=15960 $Y=96800
X1907 2 digital_ldo_top_VIA1 $T=16210 102480 0 0 $X=15960 $Y=102240
X1908 2 digital_ldo_top_VIA1 $T=16210 107920 0 0 $X=15960 $Y=107680
X1909 2 digital_ldo_top_VIA1 $T=16210 113360 0 0 $X=15960 $Y=113120
X1910 2 digital_ldo_top_VIA1 $T=16210 118800 0 0 $X=15960 $Y=118560
X1911 2 digital_ldo_top_VIA1 $T=16210 124240 0 0 $X=15960 $Y=124000
X1912 2 digital_ldo_top_VIA1 $T=16210 129680 0 0 $X=15960 $Y=129440
X1913 3 digital_ldo_top_VIA1 $T=18510 12720 0 0 $X=18260 $Y=12480
X1914 3 digital_ldo_top_VIA1 $T=18510 34480 0 0 $X=18260 $Y=34240
X1915 3 digital_ldo_top_VIA1 $T=18510 39920 0 0 $X=18260 $Y=39680
X1916 3 digital_ldo_top_VIA1 $T=18510 45360 0 0 $X=18260 $Y=45120
X1917 3 digital_ldo_top_VIA1 $T=18510 50800 0 0 $X=18260 $Y=50560
X1918 3 digital_ldo_top_VIA1 $T=18510 56240 0 0 $X=18260 $Y=56000
X1919 3 digital_ldo_top_VIA1 $T=18510 61680 0 0 $X=18260 $Y=61440
X1920 3 digital_ldo_top_VIA1 $T=18510 67120 0 0 $X=18260 $Y=66880
X1921 3 digital_ldo_top_VIA1 $T=18510 72560 0 0 $X=18260 $Y=72320
X1922 3 digital_ldo_top_VIA1 $T=18510 78000 0 0 $X=18260 $Y=77760
X1923 3 digital_ldo_top_VIA1 $T=18510 83440 0 0 $X=18260 $Y=83200
X1924 3 digital_ldo_top_VIA1 $T=18510 88880 0 0 $X=18260 $Y=88640
X1925 3 digital_ldo_top_VIA1 $T=18510 94320 0 0 $X=18260 $Y=94080
X1926 3 digital_ldo_top_VIA1 $T=18510 99760 0 0 $X=18260 $Y=99520
X1927 3 digital_ldo_top_VIA1 $T=18510 105200 0 0 $X=18260 $Y=104960
X1928 3 digital_ldo_top_VIA1 $T=18510 110640 0 0 $X=18260 $Y=110400
X1929 3 digital_ldo_top_VIA1 $T=18510 116080 0 0 $X=18260 $Y=115840
X1930 3 digital_ldo_top_VIA1 $T=18510 121520 0 0 $X=18260 $Y=121280
X1931 3 digital_ldo_top_VIA1 $T=18510 126960 0 0 $X=18260 $Y=126720
X1932 2 digital_ldo_top_VIA1 $T=19890 37200 0 0 $X=19640 $Y=36960
X1933 2 digital_ldo_top_VIA1 $T=19890 42640 0 0 $X=19640 $Y=42400
X1934 2 digital_ldo_top_VIA1 $T=19890 48080 0 0 $X=19640 $Y=47840
X1935 2 digital_ldo_top_VIA1 $T=19890 53520 0 0 $X=19640 $Y=53280
X1936 2 digital_ldo_top_VIA1 $T=19890 58960 0 0 $X=19640 $Y=58720
X1937 2 digital_ldo_top_VIA1 $T=19890 64400 0 0 $X=19640 $Y=64160
X1938 2 digital_ldo_top_VIA1 $T=19890 69840 0 0 $X=19640 $Y=69600
X1939 2 digital_ldo_top_VIA1 $T=19890 75280 0 0 $X=19640 $Y=75040
X1940 2 digital_ldo_top_VIA1 $T=19890 80720 0 0 $X=19640 $Y=80480
X1941 2 digital_ldo_top_VIA1 $T=19890 86160 0 0 $X=19640 $Y=85920
X1942 2 digital_ldo_top_VIA1 $T=19890 91600 0 0 $X=19640 $Y=91360
X1943 2 digital_ldo_top_VIA1 $T=19890 97040 0 0 $X=19640 $Y=96800
X1944 2 digital_ldo_top_VIA1 $T=19890 102480 0 0 $X=19640 $Y=102240
X1945 2 digital_ldo_top_VIA1 $T=19890 107920 0 0 $X=19640 $Y=107680
X1946 2 digital_ldo_top_VIA1 $T=19890 113360 0 0 $X=19640 $Y=113120
X1947 2 digital_ldo_top_VIA1 $T=19890 118800 0 0 $X=19640 $Y=118560
X1948 2 digital_ldo_top_VIA1 $T=19890 124240 0 0 $X=19640 $Y=124000
X1949 2 digital_ldo_top_VIA1 $T=19890 129680 0 0 $X=19640 $Y=129440
X1950 3 digital_ldo_top_VIA1 $T=22190 12720 0 0 $X=21940 $Y=12480
X1951 3 digital_ldo_top_VIA1 $T=22190 34480 0 0 $X=21940 $Y=34240
X1952 3 digital_ldo_top_VIA1 $T=22190 39920 0 0 $X=21940 $Y=39680
X1953 3 digital_ldo_top_VIA1 $T=22190 45360 0 0 $X=21940 $Y=45120
X1954 3 digital_ldo_top_VIA1 $T=22190 50800 0 0 $X=21940 $Y=50560
X1955 3 digital_ldo_top_VIA1 $T=22190 56240 0 0 $X=21940 $Y=56000
X1956 3 digital_ldo_top_VIA1 $T=22190 61680 0 0 $X=21940 $Y=61440
X1957 3 digital_ldo_top_VIA1 $T=22190 67120 0 0 $X=21940 $Y=66880
X1958 3 digital_ldo_top_VIA1 $T=22190 72560 0 0 $X=21940 $Y=72320
X1959 3 digital_ldo_top_VIA1 $T=22190 78000 0 0 $X=21940 $Y=77760
X1960 3 digital_ldo_top_VIA1 $T=22190 83440 0 0 $X=21940 $Y=83200
X1961 3 digital_ldo_top_VIA1 $T=22190 88880 0 0 $X=21940 $Y=88640
X1962 3 digital_ldo_top_VIA1 $T=22190 94320 0 0 $X=21940 $Y=94080
X1963 3 digital_ldo_top_VIA1 $T=22190 99760 0 0 $X=21940 $Y=99520
X1964 3 digital_ldo_top_VIA1 $T=22190 105200 0 0 $X=21940 $Y=104960
X1965 3 digital_ldo_top_VIA1 $T=22190 110640 0 0 $X=21940 $Y=110400
X1966 3 digital_ldo_top_VIA1 $T=22190 116080 0 0 $X=21940 $Y=115840
X1967 3 digital_ldo_top_VIA1 $T=22190 121520 0 0 $X=21940 $Y=121280
X1968 3 digital_ldo_top_VIA1 $T=22190 126960 0 0 $X=21940 $Y=126720
X1969 2 digital_ldo_top_VIA1 $T=23570 37200 0 0 $X=23320 $Y=36960
X1970 2 digital_ldo_top_VIA1 $T=23570 42640 0 0 $X=23320 $Y=42400
X1971 2 digital_ldo_top_VIA1 $T=23570 48080 0 0 $X=23320 $Y=47840
X1972 2 digital_ldo_top_VIA1 $T=23570 53520 0 0 $X=23320 $Y=53280
X1973 2 digital_ldo_top_VIA1 $T=23570 58960 0 0 $X=23320 $Y=58720
X1974 2 digital_ldo_top_VIA1 $T=23570 64400 0 0 $X=23320 $Y=64160
X1975 2 digital_ldo_top_VIA1 $T=23570 69840 0 0 $X=23320 $Y=69600
X1976 2 digital_ldo_top_VIA1 $T=23570 75280 0 0 $X=23320 $Y=75040
X1977 2 digital_ldo_top_VIA1 $T=23570 80720 0 0 $X=23320 $Y=80480
X1978 2 digital_ldo_top_VIA1 $T=23570 86160 0 0 $X=23320 $Y=85920
X1979 2 digital_ldo_top_VIA1 $T=23570 91600 0 0 $X=23320 $Y=91360
X1980 2 digital_ldo_top_VIA1 $T=23570 97040 0 0 $X=23320 $Y=96800
X1981 2 digital_ldo_top_VIA1 $T=23570 102480 0 0 $X=23320 $Y=102240
X1982 2 digital_ldo_top_VIA1 $T=23570 107920 0 0 $X=23320 $Y=107680
X1983 2 digital_ldo_top_VIA1 $T=23570 113360 0 0 $X=23320 $Y=113120
X1984 2 digital_ldo_top_VIA1 $T=23570 118800 0 0 $X=23320 $Y=118560
X1985 2 digital_ldo_top_VIA1 $T=23570 124240 0 0 $X=23320 $Y=124000
X1986 2 digital_ldo_top_VIA1 $T=23570 129680 0 0 $X=23320 $Y=129440
X1987 3 digital_ldo_top_VIA1 $T=25870 12720 0 0 $X=25620 $Y=12480
X1988 3 digital_ldo_top_VIA1 $T=25870 34480 0 0 $X=25620 $Y=34240
X1989 3 digital_ldo_top_VIA1 $T=25870 39920 0 0 $X=25620 $Y=39680
X1990 3 digital_ldo_top_VIA1 $T=25870 45360 0 0 $X=25620 $Y=45120
X1991 3 digital_ldo_top_VIA1 $T=25870 50800 0 0 $X=25620 $Y=50560
X1992 3 digital_ldo_top_VIA1 $T=25870 56240 0 0 $X=25620 $Y=56000
X1993 3 digital_ldo_top_VIA1 $T=25870 61680 0 0 $X=25620 $Y=61440
X1994 3 digital_ldo_top_VIA1 $T=25870 67120 0 0 $X=25620 $Y=66880
X1995 3 digital_ldo_top_VIA1 $T=25870 72560 0 0 $X=25620 $Y=72320
X1996 3 digital_ldo_top_VIA1 $T=25870 78000 0 0 $X=25620 $Y=77760
X1997 3 digital_ldo_top_VIA1 $T=25870 83440 0 0 $X=25620 $Y=83200
X1998 3 digital_ldo_top_VIA1 $T=25870 88880 0 0 $X=25620 $Y=88640
X1999 3 digital_ldo_top_VIA1 $T=25870 94320 0 0 $X=25620 $Y=94080
X2000 3 digital_ldo_top_VIA1 $T=25870 99760 0 0 $X=25620 $Y=99520
X2001 3 digital_ldo_top_VIA1 $T=25870 105200 0 0 $X=25620 $Y=104960
X2002 3 digital_ldo_top_VIA1 $T=25870 110640 0 0 $X=25620 $Y=110400
X2003 3 digital_ldo_top_VIA1 $T=25870 116080 0 0 $X=25620 $Y=115840
X2004 3 digital_ldo_top_VIA1 $T=25870 121520 0 0 $X=25620 $Y=121280
X2005 3 digital_ldo_top_VIA1 $T=25870 126960 0 0 $X=25620 $Y=126720
X2006 2 digital_ldo_top_VIA1 $T=27250 37200 0 0 $X=27000 $Y=36960
X2007 2 digital_ldo_top_VIA1 $T=27250 42640 0 0 $X=27000 $Y=42400
X2008 2 digital_ldo_top_VIA1 $T=27250 48080 0 0 $X=27000 $Y=47840
X2009 2 digital_ldo_top_VIA1 $T=27250 53520 0 0 $X=27000 $Y=53280
X2010 2 digital_ldo_top_VIA1 $T=27250 58960 0 0 $X=27000 $Y=58720
X2011 2 digital_ldo_top_VIA1 $T=27250 64400 0 0 $X=27000 $Y=64160
X2012 2 digital_ldo_top_VIA1 $T=27250 69840 0 0 $X=27000 $Y=69600
X2013 2 digital_ldo_top_VIA1 $T=27250 75280 0 0 $X=27000 $Y=75040
X2014 2 digital_ldo_top_VIA1 $T=27250 80720 0 0 $X=27000 $Y=80480
X2015 2 digital_ldo_top_VIA1 $T=27250 86160 0 0 $X=27000 $Y=85920
X2016 2 digital_ldo_top_VIA1 $T=27250 91600 0 0 $X=27000 $Y=91360
X2017 2 digital_ldo_top_VIA1 $T=27250 97040 0 0 $X=27000 $Y=96800
X2018 2 digital_ldo_top_VIA1 $T=27250 102480 0 0 $X=27000 $Y=102240
X2019 2 digital_ldo_top_VIA1 $T=27250 107920 0 0 $X=27000 $Y=107680
X2020 2 digital_ldo_top_VIA1 $T=27250 113360 0 0 $X=27000 $Y=113120
X2021 2 digital_ldo_top_VIA1 $T=27250 118800 0 0 $X=27000 $Y=118560
X2022 2 digital_ldo_top_VIA1 $T=27250 124240 0 0 $X=27000 $Y=124000
X2023 2 digital_ldo_top_VIA1 $T=27250 129680 0 0 $X=27000 $Y=129440
X2024 3 digital_ldo_top_VIA1 $T=29550 12720 0 0 $X=29300 $Y=12480
X2025 3 digital_ldo_top_VIA1 $T=29550 34480 0 0 $X=29300 $Y=34240
X2026 3 digital_ldo_top_VIA1 $T=29550 39920 0 0 $X=29300 $Y=39680
X2027 3 digital_ldo_top_VIA1 $T=29550 45360 0 0 $X=29300 $Y=45120
X2028 3 digital_ldo_top_VIA1 $T=29550 50800 0 0 $X=29300 $Y=50560
X2029 3 digital_ldo_top_VIA1 $T=29550 56240 0 0 $X=29300 $Y=56000
X2030 3 digital_ldo_top_VIA1 $T=29550 61680 0 0 $X=29300 $Y=61440
X2031 3 digital_ldo_top_VIA1 $T=29550 67120 0 0 $X=29300 $Y=66880
X2032 3 digital_ldo_top_VIA1 $T=29550 72560 0 0 $X=29300 $Y=72320
X2033 3 digital_ldo_top_VIA1 $T=29550 78000 0 0 $X=29300 $Y=77760
X2034 3 digital_ldo_top_VIA1 $T=29550 83440 0 0 $X=29300 $Y=83200
X2035 3 digital_ldo_top_VIA1 $T=29550 88880 0 0 $X=29300 $Y=88640
X2036 3 digital_ldo_top_VIA1 $T=29550 94320 0 0 $X=29300 $Y=94080
X2037 3 digital_ldo_top_VIA1 $T=29550 99760 0 0 $X=29300 $Y=99520
X2038 3 digital_ldo_top_VIA1 $T=29550 105200 0 0 $X=29300 $Y=104960
X2039 3 digital_ldo_top_VIA1 $T=29550 110640 0 0 $X=29300 $Y=110400
X2040 3 digital_ldo_top_VIA1 $T=29550 116080 0 0 $X=29300 $Y=115840
X2041 3 digital_ldo_top_VIA1 $T=29550 121520 0 0 $X=29300 $Y=121280
X2042 3 digital_ldo_top_VIA1 $T=29550 126960 0 0 $X=29300 $Y=126720
X2043 2 digital_ldo_top_VIA1 $T=30930 15440 0 0 $X=30680 $Y=15200
X2044 2 digital_ldo_top_VIA1 $T=30930 20880 0 0 $X=30680 $Y=20640
X2045 2 digital_ldo_top_VIA1 $T=30930 26320 0 0 $X=30680 $Y=26080
X2046 2 digital_ldo_top_VIA1 $T=30930 31760 0 0 $X=30680 $Y=31520
X2047 2 digital_ldo_top_VIA1 $T=30930 37200 0 0 $X=30680 $Y=36960
X2048 2 digital_ldo_top_VIA1 $T=30930 42640 0 0 $X=30680 $Y=42400
X2049 2 digital_ldo_top_VIA1 $T=30930 48080 0 0 $X=30680 $Y=47840
X2050 2 digital_ldo_top_VIA1 $T=30930 53520 0 0 $X=30680 $Y=53280
X2051 2 digital_ldo_top_VIA1 $T=30930 58960 0 0 $X=30680 $Y=58720
X2052 2 digital_ldo_top_VIA1 $T=30930 64400 0 0 $X=30680 $Y=64160
X2053 2 digital_ldo_top_VIA1 $T=30930 69840 0 0 $X=30680 $Y=69600
X2054 2 digital_ldo_top_VIA1 $T=30930 75280 0 0 $X=30680 $Y=75040
X2055 2 digital_ldo_top_VIA1 $T=30930 80720 0 0 $X=30680 $Y=80480
X2056 2 digital_ldo_top_VIA1 $T=30930 86160 0 0 $X=30680 $Y=85920
X2057 2 digital_ldo_top_VIA1 $T=30930 91600 0 0 $X=30680 $Y=91360
X2058 2 digital_ldo_top_VIA1 $T=30930 97040 0 0 $X=30680 $Y=96800
X2059 2 digital_ldo_top_VIA1 $T=30930 102480 0 0 $X=30680 $Y=102240
X2060 2 digital_ldo_top_VIA1 $T=30930 107920 0 0 $X=30680 $Y=107680
X2061 2 digital_ldo_top_VIA1 $T=30930 113360 0 0 $X=30680 $Y=113120
X2062 2 digital_ldo_top_VIA1 $T=30930 118800 0 0 $X=30680 $Y=118560
X2063 2 digital_ldo_top_VIA1 $T=30930 124240 0 0 $X=30680 $Y=124000
X2064 2 digital_ldo_top_VIA1 $T=30930 129680 0 0 $X=30680 $Y=129440
X2065 3 digital_ldo_top_VIA1 $T=33230 12720 0 0 $X=32980 $Y=12480
X2066 3 digital_ldo_top_VIA1 $T=33230 18160 0 0 $X=32980 $Y=17920
X2067 3 digital_ldo_top_VIA1 $T=33230 23600 0 0 $X=32980 $Y=23360
X2068 3 digital_ldo_top_VIA1 $T=33230 29040 0 0 $X=32980 $Y=28800
X2069 3 digital_ldo_top_VIA1 $T=33230 34480 0 0 $X=32980 $Y=34240
X2070 3 digital_ldo_top_VIA1 $T=33230 39920 0 0 $X=32980 $Y=39680
X2071 3 digital_ldo_top_VIA1 $T=33230 45360 0 0 $X=32980 $Y=45120
X2072 3 digital_ldo_top_VIA1 $T=33230 50800 0 0 $X=32980 $Y=50560
X2073 3 digital_ldo_top_VIA1 $T=33230 56240 0 0 $X=32980 $Y=56000
X2074 3 digital_ldo_top_VIA1 $T=33230 61680 0 0 $X=32980 $Y=61440
X2075 3 digital_ldo_top_VIA1 $T=33230 67120 0 0 $X=32980 $Y=66880
X2076 3 digital_ldo_top_VIA1 $T=33230 72560 0 0 $X=32980 $Y=72320
X2077 3 digital_ldo_top_VIA1 $T=33230 78000 0 0 $X=32980 $Y=77760
X2078 3 digital_ldo_top_VIA1 $T=33230 83440 0 0 $X=32980 $Y=83200
X2079 3 digital_ldo_top_VIA1 $T=33230 88880 0 0 $X=32980 $Y=88640
X2080 3 digital_ldo_top_VIA1 $T=33230 94320 0 0 $X=32980 $Y=94080
X2081 3 digital_ldo_top_VIA1 $T=33230 99760 0 0 $X=32980 $Y=99520
X2082 3 digital_ldo_top_VIA1 $T=33230 105200 0 0 $X=32980 $Y=104960
X2083 3 digital_ldo_top_VIA1 $T=33230 110640 0 0 $X=32980 $Y=110400
X2084 3 digital_ldo_top_VIA1 $T=33230 116080 0 0 $X=32980 $Y=115840
X2085 3 digital_ldo_top_VIA1 $T=33230 121520 0 0 $X=32980 $Y=121280
X2086 3 digital_ldo_top_VIA1 $T=33230 126960 0 0 $X=32980 $Y=126720
X2087 2 digital_ldo_top_VIA1 $T=34610 15440 0 0 $X=34360 $Y=15200
X2088 2 digital_ldo_top_VIA1 $T=34610 20880 0 0 $X=34360 $Y=20640
X2089 2 digital_ldo_top_VIA1 $T=34610 26320 0 0 $X=34360 $Y=26080
X2090 2 digital_ldo_top_VIA1 $T=34610 31760 0 0 $X=34360 $Y=31520
X2091 2 digital_ldo_top_VIA1 $T=34610 37200 0 0 $X=34360 $Y=36960
X2092 2 digital_ldo_top_VIA1 $T=34610 42640 0 0 $X=34360 $Y=42400
X2093 2 digital_ldo_top_VIA1 $T=34610 48080 0 0 $X=34360 $Y=47840
X2094 2 digital_ldo_top_VIA1 $T=34610 53520 0 0 $X=34360 $Y=53280
X2095 2 digital_ldo_top_VIA1 $T=34610 58960 0 0 $X=34360 $Y=58720
X2096 2 digital_ldo_top_VIA1 $T=34610 64400 0 0 $X=34360 $Y=64160
X2097 2 digital_ldo_top_VIA1 $T=34610 69840 0 0 $X=34360 $Y=69600
X2098 2 digital_ldo_top_VIA1 $T=34610 75280 0 0 $X=34360 $Y=75040
X2099 2 digital_ldo_top_VIA1 $T=34610 80720 0 0 $X=34360 $Y=80480
X2100 2 digital_ldo_top_VIA1 $T=34610 86160 0 0 $X=34360 $Y=85920
X2101 2 digital_ldo_top_VIA1 $T=34610 91600 0 0 $X=34360 $Y=91360
X2102 2 digital_ldo_top_VIA1 $T=34610 97040 0 0 $X=34360 $Y=96800
X2103 2 digital_ldo_top_VIA1 $T=34610 102480 0 0 $X=34360 $Y=102240
X2104 2 digital_ldo_top_VIA1 $T=34610 107920 0 0 $X=34360 $Y=107680
X2105 2 digital_ldo_top_VIA1 $T=34610 113360 0 0 $X=34360 $Y=113120
X2106 2 digital_ldo_top_VIA1 $T=34610 118800 0 0 $X=34360 $Y=118560
X2107 2 digital_ldo_top_VIA1 $T=34610 124240 0 0 $X=34360 $Y=124000
X2108 2 digital_ldo_top_VIA1 $T=34610 129680 0 0 $X=34360 $Y=129440
X2109 3 digital_ldo_top_VIA1 $T=36910 12720 0 0 $X=36660 $Y=12480
X2110 3 digital_ldo_top_VIA1 $T=36910 18160 0 0 $X=36660 $Y=17920
X2111 3 digital_ldo_top_VIA1 $T=36910 23600 0 0 $X=36660 $Y=23360
X2112 3 digital_ldo_top_VIA1 $T=36910 29040 0 0 $X=36660 $Y=28800
X2113 3 digital_ldo_top_VIA1 $T=36910 34480 0 0 $X=36660 $Y=34240
X2114 3 digital_ldo_top_VIA1 $T=36910 39920 0 0 $X=36660 $Y=39680
X2115 3 digital_ldo_top_VIA1 $T=36910 45360 0 0 $X=36660 $Y=45120
X2116 3 digital_ldo_top_VIA1 $T=36910 50800 0 0 $X=36660 $Y=50560
X2117 3 digital_ldo_top_VIA1 $T=36910 56240 0 0 $X=36660 $Y=56000
X2118 3 digital_ldo_top_VIA1 $T=36910 61680 0 0 $X=36660 $Y=61440
X2119 3 digital_ldo_top_VIA1 $T=36910 67120 0 0 $X=36660 $Y=66880
X2120 3 digital_ldo_top_VIA1 $T=36910 72560 0 0 $X=36660 $Y=72320
X2121 3 digital_ldo_top_VIA1 $T=36910 78000 0 0 $X=36660 $Y=77760
X2122 3 digital_ldo_top_VIA1 $T=36910 83440 0 0 $X=36660 $Y=83200
X2123 3 digital_ldo_top_VIA1 $T=36910 88880 0 0 $X=36660 $Y=88640
X2124 3 digital_ldo_top_VIA1 $T=36910 94320 0 0 $X=36660 $Y=94080
X2125 3 digital_ldo_top_VIA1 $T=36910 99760 0 0 $X=36660 $Y=99520
X2126 3 digital_ldo_top_VIA1 $T=36910 105200 0 0 $X=36660 $Y=104960
X2127 3 digital_ldo_top_VIA1 $T=36910 110640 0 0 $X=36660 $Y=110400
X2128 3 digital_ldo_top_VIA1 $T=36910 116080 0 0 $X=36660 $Y=115840
X2129 3 digital_ldo_top_VIA1 $T=36910 121520 0 0 $X=36660 $Y=121280
X2130 3 digital_ldo_top_VIA1 $T=36910 126960 0 0 $X=36660 $Y=126720
X2131 2 digital_ldo_top_VIA1 $T=38290 64400 0 0 $X=38040 $Y=64160
X2132 2 digital_ldo_top_VIA1 $T=38290 69840 0 0 $X=38040 $Y=69600
X2133 2 digital_ldo_top_VIA1 $T=38290 75280 0 0 $X=38040 $Y=75040
X2134 2 digital_ldo_top_VIA1 $T=38290 80720 0 0 $X=38040 $Y=80480
X2135 2 digital_ldo_top_VIA1 $T=38290 86160 0 0 $X=38040 $Y=85920
X2136 2 digital_ldo_top_VIA1 $T=38290 91600 0 0 $X=38040 $Y=91360
X2137 2 digital_ldo_top_VIA1 $T=38290 97040 0 0 $X=38040 $Y=96800
X2138 2 digital_ldo_top_VIA1 $T=38290 102480 0 0 $X=38040 $Y=102240
X2139 2 digital_ldo_top_VIA1 $T=38290 107920 0 0 $X=38040 $Y=107680
X2140 2 digital_ldo_top_VIA1 $T=38290 113360 0 0 $X=38040 $Y=113120
X2141 2 digital_ldo_top_VIA1 $T=38290 118800 0 0 $X=38040 $Y=118560
X2142 2 digital_ldo_top_VIA1 $T=38290 124240 0 0 $X=38040 $Y=124000
X2143 2 digital_ldo_top_VIA1 $T=38290 129680 0 0 $X=38040 $Y=129440
X2144 3 digital_ldo_top_VIA1 $T=40590 12720 0 0 $X=40340 $Y=12480
X2145 3 digital_ldo_top_VIA1 $T=40590 67120 0 0 $X=40340 $Y=66880
X2146 3 digital_ldo_top_VIA1 $T=40590 72560 0 0 $X=40340 $Y=72320
X2147 3 digital_ldo_top_VIA1 $T=40590 78000 0 0 $X=40340 $Y=77760
X2148 3 digital_ldo_top_VIA1 $T=40590 83440 0 0 $X=40340 $Y=83200
X2149 3 digital_ldo_top_VIA1 $T=40590 88880 0 0 $X=40340 $Y=88640
X2150 3 digital_ldo_top_VIA1 $T=40590 94320 0 0 $X=40340 $Y=94080
X2151 3 digital_ldo_top_VIA1 $T=40590 99760 0 0 $X=40340 $Y=99520
X2152 3 digital_ldo_top_VIA1 $T=40590 105200 0 0 $X=40340 $Y=104960
X2153 3 digital_ldo_top_VIA1 $T=40590 110640 0 0 $X=40340 $Y=110400
X2154 3 digital_ldo_top_VIA1 $T=40590 116080 0 0 $X=40340 $Y=115840
X2155 3 digital_ldo_top_VIA1 $T=40590 121520 0 0 $X=40340 $Y=121280
X2156 3 digital_ldo_top_VIA1 $T=40590 126960 0 0 $X=40340 $Y=126720
X2157 2 digital_ldo_top_VIA1 $T=41970 64400 0 0 $X=41720 $Y=64160
X2158 2 digital_ldo_top_VIA1 $T=41970 69840 0 0 $X=41720 $Y=69600
X2159 2 digital_ldo_top_VIA1 $T=41970 75280 0 0 $X=41720 $Y=75040
X2160 2 digital_ldo_top_VIA1 $T=41970 80720 0 0 $X=41720 $Y=80480
X2161 2 digital_ldo_top_VIA1 $T=41970 86160 0 0 $X=41720 $Y=85920
X2162 2 digital_ldo_top_VIA1 $T=41970 91600 0 0 $X=41720 $Y=91360
X2163 2 digital_ldo_top_VIA1 $T=41970 97040 0 0 $X=41720 $Y=96800
X2164 2 digital_ldo_top_VIA1 $T=41970 102480 0 0 $X=41720 $Y=102240
X2165 2 digital_ldo_top_VIA1 $T=41970 107920 0 0 $X=41720 $Y=107680
X2166 2 digital_ldo_top_VIA1 $T=41970 113360 0 0 $X=41720 $Y=113120
X2167 2 digital_ldo_top_VIA1 $T=41970 118800 0 0 $X=41720 $Y=118560
X2168 2 digital_ldo_top_VIA1 $T=41970 124240 0 0 $X=41720 $Y=124000
X2169 2 digital_ldo_top_VIA1 $T=41970 129680 0 0 $X=41720 $Y=129440
X2170 3 digital_ldo_top_VIA1 $T=44270 12720 0 0 $X=44020 $Y=12480
X2171 3 digital_ldo_top_VIA1 $T=44270 67120 0 0 $X=44020 $Y=66880
X2172 3 digital_ldo_top_VIA1 $T=44270 72560 0 0 $X=44020 $Y=72320
X2173 3 digital_ldo_top_VIA1 $T=44270 78000 0 0 $X=44020 $Y=77760
X2174 3 digital_ldo_top_VIA1 $T=44270 83440 0 0 $X=44020 $Y=83200
X2175 3 digital_ldo_top_VIA1 $T=44270 88880 0 0 $X=44020 $Y=88640
X2176 3 digital_ldo_top_VIA1 $T=44270 94320 0 0 $X=44020 $Y=94080
X2177 3 digital_ldo_top_VIA1 $T=44270 99760 0 0 $X=44020 $Y=99520
X2178 3 digital_ldo_top_VIA1 $T=44270 105200 0 0 $X=44020 $Y=104960
X2179 3 digital_ldo_top_VIA1 $T=44270 110640 0 0 $X=44020 $Y=110400
X2180 3 digital_ldo_top_VIA1 $T=44270 116080 0 0 $X=44020 $Y=115840
X2181 3 digital_ldo_top_VIA1 $T=44270 121520 0 0 $X=44020 $Y=121280
X2182 3 digital_ldo_top_VIA1 $T=44270 126960 0 0 $X=44020 $Y=126720
X2183 2 digital_ldo_top_VIA1 $T=45650 64400 0 0 $X=45400 $Y=64160
X2184 2 digital_ldo_top_VIA1 $T=45650 69840 0 0 $X=45400 $Y=69600
X2185 2 digital_ldo_top_VIA1 $T=45650 75280 0 0 $X=45400 $Y=75040
X2186 2 digital_ldo_top_VIA1 $T=45650 80720 0 0 $X=45400 $Y=80480
X2187 2 digital_ldo_top_VIA1 $T=45650 86160 0 0 $X=45400 $Y=85920
X2188 2 digital_ldo_top_VIA1 $T=45650 91600 0 0 $X=45400 $Y=91360
X2189 2 digital_ldo_top_VIA1 $T=45650 97040 0 0 $X=45400 $Y=96800
X2190 2 digital_ldo_top_VIA1 $T=45650 102480 0 0 $X=45400 $Y=102240
X2191 2 digital_ldo_top_VIA1 $T=45650 107920 0 0 $X=45400 $Y=107680
X2192 2 digital_ldo_top_VIA1 $T=45650 113360 0 0 $X=45400 $Y=113120
X2193 2 digital_ldo_top_VIA1 $T=45650 118800 0 0 $X=45400 $Y=118560
X2194 2 digital_ldo_top_VIA1 $T=45650 124240 0 0 $X=45400 $Y=124000
X2195 2 digital_ldo_top_VIA1 $T=45650 129680 0 0 $X=45400 $Y=129440
X2196 3 digital_ldo_top_VIA1 $T=47950 12720 0 0 $X=47700 $Y=12480
X2197 3 digital_ldo_top_VIA1 $T=47950 67120 0 0 $X=47700 $Y=66880
X2198 3 digital_ldo_top_VIA1 $T=47950 72560 0 0 $X=47700 $Y=72320
X2199 3 digital_ldo_top_VIA1 $T=47950 78000 0 0 $X=47700 $Y=77760
X2200 3 digital_ldo_top_VIA1 $T=47950 83440 0 0 $X=47700 $Y=83200
X2201 3 digital_ldo_top_VIA1 $T=47950 88880 0 0 $X=47700 $Y=88640
X2202 3 digital_ldo_top_VIA1 $T=47950 94320 0 0 $X=47700 $Y=94080
X2203 3 digital_ldo_top_VIA1 $T=47950 99760 0 0 $X=47700 $Y=99520
X2204 3 digital_ldo_top_VIA1 $T=47950 105200 0 0 $X=47700 $Y=104960
X2205 3 digital_ldo_top_VIA1 $T=47950 110640 0 0 $X=47700 $Y=110400
X2206 3 digital_ldo_top_VIA1 $T=47950 116080 0 0 $X=47700 $Y=115840
X2207 3 digital_ldo_top_VIA1 $T=47950 121520 0 0 $X=47700 $Y=121280
X2208 3 digital_ldo_top_VIA1 $T=47950 126960 0 0 $X=47700 $Y=126720
X2209 2 digital_ldo_top_VIA1 $T=49330 64400 0 0 $X=49080 $Y=64160
X2210 2 digital_ldo_top_VIA1 $T=49330 69840 0 0 $X=49080 $Y=69600
X2211 2 digital_ldo_top_VIA1 $T=49330 75280 0 0 $X=49080 $Y=75040
X2212 2 digital_ldo_top_VIA1 $T=49330 80720 0 0 $X=49080 $Y=80480
X2213 2 digital_ldo_top_VIA1 $T=49330 86160 0 0 $X=49080 $Y=85920
X2214 2 digital_ldo_top_VIA1 $T=49330 91600 0 0 $X=49080 $Y=91360
X2215 2 digital_ldo_top_VIA1 $T=49330 97040 0 0 $X=49080 $Y=96800
X2216 2 digital_ldo_top_VIA1 $T=49330 102480 0 0 $X=49080 $Y=102240
X2217 2 digital_ldo_top_VIA1 $T=49330 107920 0 0 $X=49080 $Y=107680
X2218 2 digital_ldo_top_VIA1 $T=49330 113360 0 0 $X=49080 $Y=113120
X2219 2 digital_ldo_top_VIA1 $T=49330 118800 0 0 $X=49080 $Y=118560
X2220 2 digital_ldo_top_VIA1 $T=49330 124240 0 0 $X=49080 $Y=124000
X2221 2 digital_ldo_top_VIA1 $T=49330 129680 0 0 $X=49080 $Y=129440
X2222 3 digital_ldo_top_VIA1 $T=51630 12720 0 0 $X=51380 $Y=12480
X2223 3 digital_ldo_top_VIA1 $T=51630 67120 0 0 $X=51380 $Y=66880
X2224 3 digital_ldo_top_VIA1 $T=51630 72560 0 0 $X=51380 $Y=72320
X2225 3 digital_ldo_top_VIA1 $T=51630 78000 0 0 $X=51380 $Y=77760
X2226 3 digital_ldo_top_VIA1 $T=51630 83440 0 0 $X=51380 $Y=83200
X2227 3 digital_ldo_top_VIA1 $T=51630 88880 0 0 $X=51380 $Y=88640
X2228 3 digital_ldo_top_VIA1 $T=51630 94320 0 0 $X=51380 $Y=94080
X2229 3 digital_ldo_top_VIA1 $T=51630 99760 0 0 $X=51380 $Y=99520
X2230 3 digital_ldo_top_VIA1 $T=51630 105200 0 0 $X=51380 $Y=104960
X2231 3 digital_ldo_top_VIA1 $T=51630 110640 0 0 $X=51380 $Y=110400
X2232 3 digital_ldo_top_VIA1 $T=51630 116080 0 0 $X=51380 $Y=115840
X2233 3 digital_ldo_top_VIA1 $T=51630 121520 0 0 $X=51380 $Y=121280
X2234 3 digital_ldo_top_VIA1 $T=51630 126960 0 0 $X=51380 $Y=126720
X2235 2 digital_ldo_top_VIA1 $T=53010 64400 0 0 $X=52760 $Y=64160
X2236 2 digital_ldo_top_VIA1 $T=53010 69840 0 0 $X=52760 $Y=69600
X2237 2 digital_ldo_top_VIA1 $T=53010 75280 0 0 $X=52760 $Y=75040
X2238 2 digital_ldo_top_VIA1 $T=53010 80720 0 0 $X=52760 $Y=80480
X2239 2 digital_ldo_top_VIA1 $T=53010 86160 0 0 $X=52760 $Y=85920
X2240 2 digital_ldo_top_VIA1 $T=53010 91600 0 0 $X=52760 $Y=91360
X2241 2 digital_ldo_top_VIA1 $T=53010 97040 0 0 $X=52760 $Y=96800
X2242 2 digital_ldo_top_VIA1 $T=53010 102480 0 0 $X=52760 $Y=102240
X2243 2 digital_ldo_top_VIA1 $T=53010 107920 0 0 $X=52760 $Y=107680
X2244 2 digital_ldo_top_VIA1 $T=53010 113360 0 0 $X=52760 $Y=113120
X2245 2 digital_ldo_top_VIA1 $T=53010 118800 0 0 $X=52760 $Y=118560
X2246 2 digital_ldo_top_VIA1 $T=53010 124240 0 0 $X=52760 $Y=124000
X2247 2 digital_ldo_top_VIA1 $T=53010 129680 0 0 $X=52760 $Y=129440
X2248 3 digital_ldo_top_VIA1 $T=55310 12720 0 0 $X=55060 $Y=12480
X2249 3 digital_ldo_top_VIA1 $T=55310 18160 0 0 $X=55060 $Y=17920
X2250 3 digital_ldo_top_VIA1 $T=55310 23600 0 0 $X=55060 $Y=23360
X2251 3 digital_ldo_top_VIA1 $T=55310 29040 0 0 $X=55060 $Y=28800
X2252 3 digital_ldo_top_VIA1 $T=55310 34480 0 0 $X=55060 $Y=34240
X2253 3 digital_ldo_top_VIA1 $T=55310 39920 0 0 $X=55060 $Y=39680
X2254 3 digital_ldo_top_VIA1 $T=55310 45360 0 0 $X=55060 $Y=45120
X2255 3 digital_ldo_top_VIA1 $T=55310 50800 0 0 $X=55060 $Y=50560
X2256 3 digital_ldo_top_VIA1 $T=55310 56240 0 0 $X=55060 $Y=56000
X2257 3 digital_ldo_top_VIA1 $T=55310 61680 0 0 $X=55060 $Y=61440
X2258 3 digital_ldo_top_VIA1 $T=55310 67120 0 0 $X=55060 $Y=66880
X2259 3 digital_ldo_top_VIA1 $T=55310 72560 0 0 $X=55060 $Y=72320
X2260 3 digital_ldo_top_VIA1 $T=55310 78000 0 0 $X=55060 $Y=77760
X2261 3 digital_ldo_top_VIA1 $T=55310 83440 0 0 $X=55060 $Y=83200
X2262 3 digital_ldo_top_VIA1 $T=55310 88880 0 0 $X=55060 $Y=88640
X2263 3 digital_ldo_top_VIA1 $T=55310 94320 0 0 $X=55060 $Y=94080
X2264 3 digital_ldo_top_VIA1 $T=55310 99760 0 0 $X=55060 $Y=99520
X2265 3 digital_ldo_top_VIA1 $T=55310 105200 0 0 $X=55060 $Y=104960
X2266 3 digital_ldo_top_VIA1 $T=55310 110640 0 0 $X=55060 $Y=110400
X2267 3 digital_ldo_top_VIA1 $T=55310 116080 0 0 $X=55060 $Y=115840
X2268 3 digital_ldo_top_VIA1 $T=55310 121520 0 0 $X=55060 $Y=121280
X2269 3 digital_ldo_top_VIA1 $T=55310 126960 0 0 $X=55060 $Y=126720
X2270 2 digital_ldo_top_VIA1 $T=56690 15440 0 0 $X=56440 $Y=15200
X2271 2 digital_ldo_top_VIA1 $T=56690 20880 0 0 $X=56440 $Y=20640
X2272 2 digital_ldo_top_VIA1 $T=56690 26320 0 0 $X=56440 $Y=26080
X2273 2 digital_ldo_top_VIA1 $T=56690 31760 0 0 $X=56440 $Y=31520
X2274 2 digital_ldo_top_VIA1 $T=56690 37200 0 0 $X=56440 $Y=36960
X2275 2 digital_ldo_top_VIA1 $T=56690 42640 0 0 $X=56440 $Y=42400
X2276 2 digital_ldo_top_VIA1 $T=56690 48080 0 0 $X=56440 $Y=47840
X2277 2 digital_ldo_top_VIA1 $T=56690 53520 0 0 $X=56440 $Y=53280
X2278 2 digital_ldo_top_VIA1 $T=56690 58960 0 0 $X=56440 $Y=58720
X2279 2 digital_ldo_top_VIA1 $T=56690 64400 0 0 $X=56440 $Y=64160
X2280 2 digital_ldo_top_VIA1 $T=56690 69840 0 0 $X=56440 $Y=69600
X2281 2 digital_ldo_top_VIA1 $T=56690 75280 0 0 $X=56440 $Y=75040
X2282 2 digital_ldo_top_VIA1 $T=56690 80720 0 0 $X=56440 $Y=80480
X2283 2 digital_ldo_top_VIA1 $T=56690 86160 0 0 $X=56440 $Y=85920
X2284 2 digital_ldo_top_VIA1 $T=56690 91600 0 0 $X=56440 $Y=91360
X2285 2 digital_ldo_top_VIA1 $T=56690 97040 0 0 $X=56440 $Y=96800
X2286 2 digital_ldo_top_VIA1 $T=56690 102480 0 0 $X=56440 $Y=102240
X2287 2 digital_ldo_top_VIA1 $T=56690 107920 0 0 $X=56440 $Y=107680
X2288 2 digital_ldo_top_VIA1 $T=56690 113360 0 0 $X=56440 $Y=113120
X2289 2 digital_ldo_top_VIA1 $T=56690 118800 0 0 $X=56440 $Y=118560
X2290 2 digital_ldo_top_VIA1 $T=56690 124240 0 0 $X=56440 $Y=124000
X2291 2 digital_ldo_top_VIA1 $T=56690 129680 0 0 $X=56440 $Y=129440
X2292 3 digital_ldo_top_VIA1 $T=58990 12720 0 0 $X=58740 $Y=12480
X2293 3 digital_ldo_top_VIA1 $T=58990 34480 0 0 $X=58740 $Y=34240
X2294 3 digital_ldo_top_VIA1 $T=58990 39920 0 0 $X=58740 $Y=39680
X2295 3 digital_ldo_top_VIA1 $T=58990 45360 0 0 $X=58740 $Y=45120
X2296 3 digital_ldo_top_VIA1 $T=58990 50800 0 0 $X=58740 $Y=50560
X2297 3 digital_ldo_top_VIA1 $T=58990 56240 0 0 $X=58740 $Y=56000
X2298 3 digital_ldo_top_VIA1 $T=58990 61680 0 0 $X=58740 $Y=61440
X2299 3 digital_ldo_top_VIA1 $T=58990 67120 0 0 $X=58740 $Y=66880
X2300 3 digital_ldo_top_VIA1 $T=58990 72560 0 0 $X=58740 $Y=72320
X2301 3 digital_ldo_top_VIA1 $T=58990 78000 0 0 $X=58740 $Y=77760
X2302 3 digital_ldo_top_VIA1 $T=58990 83440 0 0 $X=58740 $Y=83200
X2303 3 digital_ldo_top_VIA1 $T=58990 88880 0 0 $X=58740 $Y=88640
X2304 3 digital_ldo_top_VIA1 $T=58990 94320 0 0 $X=58740 $Y=94080
X2305 3 digital_ldo_top_VIA1 $T=58990 99760 0 0 $X=58740 $Y=99520
X2306 3 digital_ldo_top_VIA1 $T=58990 105200 0 0 $X=58740 $Y=104960
X2307 3 digital_ldo_top_VIA1 $T=58990 110640 0 0 $X=58740 $Y=110400
X2308 3 digital_ldo_top_VIA1 $T=58990 116080 0 0 $X=58740 $Y=115840
X2309 3 digital_ldo_top_VIA1 $T=58990 121520 0 0 $X=58740 $Y=121280
X2310 3 digital_ldo_top_VIA1 $T=58990 126960 0 0 $X=58740 $Y=126720
X2311 2 digital_ldo_top_VIA1 $T=60370 37200 0 0 $X=60120 $Y=36960
X2312 2 digital_ldo_top_VIA1 $T=60370 42640 0 0 $X=60120 $Y=42400
X2313 2 digital_ldo_top_VIA1 $T=60370 48080 0 0 $X=60120 $Y=47840
X2314 2 digital_ldo_top_VIA1 $T=60370 53520 0 0 $X=60120 $Y=53280
X2315 2 digital_ldo_top_VIA1 $T=60370 58960 0 0 $X=60120 $Y=58720
X2316 2 digital_ldo_top_VIA1 $T=60370 64400 0 0 $X=60120 $Y=64160
X2317 2 digital_ldo_top_VIA1 $T=60370 69840 0 0 $X=60120 $Y=69600
X2318 2 digital_ldo_top_VIA1 $T=60370 75280 0 0 $X=60120 $Y=75040
X2319 2 digital_ldo_top_VIA1 $T=60370 80720 0 0 $X=60120 $Y=80480
X2320 2 digital_ldo_top_VIA1 $T=60370 86160 0 0 $X=60120 $Y=85920
X2321 2 digital_ldo_top_VIA1 $T=60370 91600 0 0 $X=60120 $Y=91360
X2322 2 digital_ldo_top_VIA1 $T=60370 97040 0 0 $X=60120 $Y=96800
X2323 2 digital_ldo_top_VIA1 $T=60370 102480 0 0 $X=60120 $Y=102240
X2324 2 digital_ldo_top_VIA1 $T=60370 107920 0 0 $X=60120 $Y=107680
X2325 2 digital_ldo_top_VIA1 $T=60370 113360 0 0 $X=60120 $Y=113120
X2326 2 digital_ldo_top_VIA1 $T=60370 118800 0 0 $X=60120 $Y=118560
X2327 2 digital_ldo_top_VIA1 $T=60370 124240 0 0 $X=60120 $Y=124000
X2328 2 digital_ldo_top_VIA1 $T=60370 129680 0 0 $X=60120 $Y=129440
X2329 3 digital_ldo_top_VIA1 $T=62670 12720 0 0 $X=62420 $Y=12480
X2330 3 digital_ldo_top_VIA1 $T=62670 34480 0 0 $X=62420 $Y=34240
X2331 3 digital_ldo_top_VIA1 $T=62670 39920 0 0 $X=62420 $Y=39680
X2332 3 digital_ldo_top_VIA1 $T=62670 45360 0 0 $X=62420 $Y=45120
X2333 3 digital_ldo_top_VIA1 $T=62670 50800 0 0 $X=62420 $Y=50560
X2334 3 digital_ldo_top_VIA1 $T=62670 56240 0 0 $X=62420 $Y=56000
X2335 3 digital_ldo_top_VIA1 $T=62670 61680 0 0 $X=62420 $Y=61440
X2336 3 digital_ldo_top_VIA1 $T=62670 67120 0 0 $X=62420 $Y=66880
X2337 3 digital_ldo_top_VIA1 $T=62670 72560 0 0 $X=62420 $Y=72320
X2338 3 digital_ldo_top_VIA1 $T=62670 78000 0 0 $X=62420 $Y=77760
X2339 3 digital_ldo_top_VIA1 $T=62670 83440 0 0 $X=62420 $Y=83200
X2340 3 digital_ldo_top_VIA1 $T=62670 88880 0 0 $X=62420 $Y=88640
X2341 3 digital_ldo_top_VIA1 $T=62670 94320 0 0 $X=62420 $Y=94080
X2342 3 digital_ldo_top_VIA1 $T=62670 99760 0 0 $X=62420 $Y=99520
X2343 3 digital_ldo_top_VIA1 $T=62670 105200 0 0 $X=62420 $Y=104960
X2344 3 digital_ldo_top_VIA1 $T=62670 110640 0 0 $X=62420 $Y=110400
X2345 3 digital_ldo_top_VIA1 $T=62670 116080 0 0 $X=62420 $Y=115840
X2346 3 digital_ldo_top_VIA1 $T=62670 121520 0 0 $X=62420 $Y=121280
X2347 3 digital_ldo_top_VIA1 $T=62670 126960 0 0 $X=62420 $Y=126720
X2348 2 digital_ldo_top_VIA1 $T=64050 37200 0 0 $X=63800 $Y=36960
X2349 2 digital_ldo_top_VIA1 $T=64050 42640 0 0 $X=63800 $Y=42400
X2350 2 digital_ldo_top_VIA1 $T=64050 48080 0 0 $X=63800 $Y=47840
X2351 2 digital_ldo_top_VIA1 $T=64050 53520 0 0 $X=63800 $Y=53280
X2352 2 digital_ldo_top_VIA1 $T=64050 58960 0 0 $X=63800 $Y=58720
X2353 2 digital_ldo_top_VIA1 $T=64050 64400 0 0 $X=63800 $Y=64160
X2354 2 digital_ldo_top_VIA1 $T=64050 69840 0 0 $X=63800 $Y=69600
X2355 2 digital_ldo_top_VIA1 $T=64050 75280 0 0 $X=63800 $Y=75040
X2356 2 digital_ldo_top_VIA1 $T=64050 80720 0 0 $X=63800 $Y=80480
X2357 2 digital_ldo_top_VIA1 $T=64050 86160 0 0 $X=63800 $Y=85920
X2358 2 digital_ldo_top_VIA1 $T=64050 91600 0 0 $X=63800 $Y=91360
X2359 2 digital_ldo_top_VIA1 $T=64050 97040 0 0 $X=63800 $Y=96800
X2360 2 digital_ldo_top_VIA1 $T=64050 102480 0 0 $X=63800 $Y=102240
X2361 2 digital_ldo_top_VIA1 $T=64050 107920 0 0 $X=63800 $Y=107680
X2362 2 digital_ldo_top_VIA1 $T=64050 113360 0 0 $X=63800 $Y=113120
X2363 2 digital_ldo_top_VIA1 $T=64050 118800 0 0 $X=63800 $Y=118560
X2364 2 digital_ldo_top_VIA1 $T=64050 124240 0 0 $X=63800 $Y=124000
X2365 2 digital_ldo_top_VIA1 $T=64050 129680 0 0 $X=63800 $Y=129440
X2366 3 digital_ldo_top_VIA1 $T=66350 12720 0 0 $X=66100 $Y=12480
X2367 3 digital_ldo_top_VIA1 $T=66350 34480 0 0 $X=66100 $Y=34240
X2368 3 digital_ldo_top_VIA1 $T=66350 39920 0 0 $X=66100 $Y=39680
X2369 3 digital_ldo_top_VIA1 $T=66350 45360 0 0 $X=66100 $Y=45120
X2370 3 digital_ldo_top_VIA1 $T=66350 50800 0 0 $X=66100 $Y=50560
X2371 3 digital_ldo_top_VIA1 $T=66350 56240 0 0 $X=66100 $Y=56000
X2372 3 digital_ldo_top_VIA1 $T=66350 61680 0 0 $X=66100 $Y=61440
X2373 3 digital_ldo_top_VIA1 $T=66350 67120 0 0 $X=66100 $Y=66880
X2374 3 digital_ldo_top_VIA1 $T=66350 72560 0 0 $X=66100 $Y=72320
X2375 3 digital_ldo_top_VIA1 $T=66350 78000 0 0 $X=66100 $Y=77760
X2376 3 digital_ldo_top_VIA1 $T=66350 83440 0 0 $X=66100 $Y=83200
X2377 3 digital_ldo_top_VIA1 $T=66350 88880 0 0 $X=66100 $Y=88640
X2378 3 digital_ldo_top_VIA1 $T=66350 94320 0 0 $X=66100 $Y=94080
X2379 3 digital_ldo_top_VIA1 $T=66350 99760 0 0 $X=66100 $Y=99520
X2380 3 digital_ldo_top_VIA1 $T=66350 105200 0 0 $X=66100 $Y=104960
X2381 3 digital_ldo_top_VIA1 $T=66350 110640 0 0 $X=66100 $Y=110400
X2382 3 digital_ldo_top_VIA1 $T=66350 116080 0 0 $X=66100 $Y=115840
X2383 3 digital_ldo_top_VIA1 $T=66350 121520 0 0 $X=66100 $Y=121280
X2384 3 digital_ldo_top_VIA1 $T=66350 126960 0 0 $X=66100 $Y=126720
X2385 2 digital_ldo_top_VIA1 $T=67730 37200 0 0 $X=67480 $Y=36960
X2386 2 digital_ldo_top_VIA1 $T=67730 42640 0 0 $X=67480 $Y=42400
X2387 2 digital_ldo_top_VIA1 $T=67730 48080 0 0 $X=67480 $Y=47840
X2388 2 digital_ldo_top_VIA1 $T=67730 53520 0 0 $X=67480 $Y=53280
X2389 2 digital_ldo_top_VIA1 $T=67730 58960 0 0 $X=67480 $Y=58720
X2390 2 digital_ldo_top_VIA1 $T=67730 64400 0 0 $X=67480 $Y=64160
X2391 2 digital_ldo_top_VIA1 $T=67730 69840 0 0 $X=67480 $Y=69600
X2392 2 digital_ldo_top_VIA1 $T=67730 75280 0 0 $X=67480 $Y=75040
X2393 2 digital_ldo_top_VIA1 $T=67730 80720 0 0 $X=67480 $Y=80480
X2394 2 digital_ldo_top_VIA1 $T=67730 86160 0 0 $X=67480 $Y=85920
X2395 2 digital_ldo_top_VIA1 $T=67730 91600 0 0 $X=67480 $Y=91360
X2396 2 digital_ldo_top_VIA1 $T=67730 97040 0 0 $X=67480 $Y=96800
X2397 2 digital_ldo_top_VIA1 $T=67730 102480 0 0 $X=67480 $Y=102240
X2398 2 digital_ldo_top_VIA1 $T=67730 107920 0 0 $X=67480 $Y=107680
X2399 2 digital_ldo_top_VIA1 $T=67730 113360 0 0 $X=67480 $Y=113120
X2400 2 digital_ldo_top_VIA1 $T=67730 118800 0 0 $X=67480 $Y=118560
X2401 2 digital_ldo_top_VIA1 $T=67730 124240 0 0 $X=67480 $Y=124000
X2402 2 digital_ldo_top_VIA1 $T=67730 129680 0 0 $X=67480 $Y=129440
X2403 3 digital_ldo_top_VIA1 $T=70030 12720 0 0 $X=69780 $Y=12480
X2404 3 digital_ldo_top_VIA1 $T=70030 34480 0 0 $X=69780 $Y=34240
X2405 3 digital_ldo_top_VIA1 $T=70030 39920 0 0 $X=69780 $Y=39680
X2406 3 digital_ldo_top_VIA1 $T=70030 45360 0 0 $X=69780 $Y=45120
X2407 3 digital_ldo_top_VIA1 $T=70030 50800 0 0 $X=69780 $Y=50560
X2408 3 digital_ldo_top_VIA1 $T=70030 56240 0 0 $X=69780 $Y=56000
X2409 3 digital_ldo_top_VIA1 $T=70030 61680 0 0 $X=69780 $Y=61440
X2410 3 digital_ldo_top_VIA1 $T=70030 67120 0 0 $X=69780 $Y=66880
X2411 3 digital_ldo_top_VIA1 $T=70030 72560 0 0 $X=69780 $Y=72320
X2412 3 digital_ldo_top_VIA1 $T=70030 78000 0 0 $X=69780 $Y=77760
X2413 3 digital_ldo_top_VIA1 $T=70030 83440 0 0 $X=69780 $Y=83200
X2414 3 digital_ldo_top_VIA1 $T=70030 88880 0 0 $X=69780 $Y=88640
X2415 3 digital_ldo_top_VIA1 $T=70030 94320 0 0 $X=69780 $Y=94080
X2416 3 digital_ldo_top_VIA1 $T=70030 99760 0 0 $X=69780 $Y=99520
X2417 3 digital_ldo_top_VIA1 $T=70030 105200 0 0 $X=69780 $Y=104960
X2418 3 digital_ldo_top_VIA1 $T=70030 110640 0 0 $X=69780 $Y=110400
X2419 3 digital_ldo_top_VIA1 $T=70030 116080 0 0 $X=69780 $Y=115840
X2420 3 digital_ldo_top_VIA1 $T=70030 121520 0 0 $X=69780 $Y=121280
X2421 3 digital_ldo_top_VIA1 $T=70030 126960 0 0 $X=69780 $Y=126720
X2422 2 digital_ldo_top_VIA1 $T=71410 37200 0 0 $X=71160 $Y=36960
X2423 2 digital_ldo_top_VIA1 $T=71410 42640 0 0 $X=71160 $Y=42400
X2424 2 digital_ldo_top_VIA1 $T=71410 48080 0 0 $X=71160 $Y=47840
X2425 2 digital_ldo_top_VIA1 $T=71410 53520 0 0 $X=71160 $Y=53280
X2426 2 digital_ldo_top_VIA1 $T=71410 58960 0 0 $X=71160 $Y=58720
X2427 2 digital_ldo_top_VIA1 $T=71410 64400 0 0 $X=71160 $Y=64160
X2428 2 digital_ldo_top_VIA1 $T=71410 69840 0 0 $X=71160 $Y=69600
X2429 2 digital_ldo_top_VIA1 $T=71410 75280 0 0 $X=71160 $Y=75040
X2430 2 digital_ldo_top_VIA1 $T=71410 80720 0 0 $X=71160 $Y=80480
X2431 2 digital_ldo_top_VIA1 $T=71410 86160 0 0 $X=71160 $Y=85920
X2432 2 digital_ldo_top_VIA1 $T=71410 91600 0 0 $X=71160 $Y=91360
X2433 2 digital_ldo_top_VIA1 $T=71410 97040 0 0 $X=71160 $Y=96800
X2434 2 digital_ldo_top_VIA1 $T=71410 102480 0 0 $X=71160 $Y=102240
X2435 2 digital_ldo_top_VIA1 $T=71410 107920 0 0 $X=71160 $Y=107680
X2436 2 digital_ldo_top_VIA1 $T=71410 113360 0 0 $X=71160 $Y=113120
X2437 2 digital_ldo_top_VIA1 $T=71410 118800 0 0 $X=71160 $Y=118560
X2438 2 digital_ldo_top_VIA1 $T=71410 124240 0 0 $X=71160 $Y=124000
X2439 2 digital_ldo_top_VIA1 $T=71410 129680 0 0 $X=71160 $Y=129440
X2440 3 digital_ldo_top_VIA1 $T=73710 12720 0 0 $X=73460 $Y=12480
X2441 3 digital_ldo_top_VIA1 $T=73710 34480 0 0 $X=73460 $Y=34240
X2442 3 digital_ldo_top_VIA1 $T=73710 39920 0 0 $X=73460 $Y=39680
X2443 3 digital_ldo_top_VIA1 $T=73710 45360 0 0 $X=73460 $Y=45120
X2444 3 digital_ldo_top_VIA1 $T=73710 50800 0 0 $X=73460 $Y=50560
X2445 3 digital_ldo_top_VIA1 $T=73710 56240 0 0 $X=73460 $Y=56000
X2446 3 digital_ldo_top_VIA1 $T=73710 61680 0 0 $X=73460 $Y=61440
X2447 3 digital_ldo_top_VIA1 $T=73710 67120 0 0 $X=73460 $Y=66880
X2448 3 digital_ldo_top_VIA1 $T=73710 72560 0 0 $X=73460 $Y=72320
X2449 3 digital_ldo_top_VIA1 $T=73710 78000 0 0 $X=73460 $Y=77760
X2450 3 digital_ldo_top_VIA1 $T=73710 83440 0 0 $X=73460 $Y=83200
X2451 3 digital_ldo_top_VIA1 $T=73710 88880 0 0 $X=73460 $Y=88640
X2452 3 digital_ldo_top_VIA1 $T=73710 94320 0 0 $X=73460 $Y=94080
X2453 3 digital_ldo_top_VIA1 $T=73710 99760 0 0 $X=73460 $Y=99520
X2454 3 digital_ldo_top_VIA1 $T=73710 105200 0 0 $X=73460 $Y=104960
X2455 3 digital_ldo_top_VIA1 $T=73710 110640 0 0 $X=73460 $Y=110400
X2456 3 digital_ldo_top_VIA1 $T=73710 116080 0 0 $X=73460 $Y=115840
X2457 3 digital_ldo_top_VIA1 $T=73710 121520 0 0 $X=73460 $Y=121280
X2458 3 digital_ldo_top_VIA1 $T=73710 126960 0 0 $X=73460 $Y=126720
X2459 2 digital_ldo_top_VIA1 $T=75090 37200 0 0 $X=74840 $Y=36960
X2460 2 digital_ldo_top_VIA1 $T=75090 42640 0 0 $X=74840 $Y=42400
X2461 2 digital_ldo_top_VIA1 $T=75090 48080 0 0 $X=74840 $Y=47840
X2462 2 digital_ldo_top_VIA1 $T=75090 53520 0 0 $X=74840 $Y=53280
X2463 2 digital_ldo_top_VIA1 $T=75090 58960 0 0 $X=74840 $Y=58720
X2464 2 digital_ldo_top_VIA1 $T=75090 64400 0 0 $X=74840 $Y=64160
X2465 2 digital_ldo_top_VIA1 $T=75090 69840 0 0 $X=74840 $Y=69600
X2466 2 digital_ldo_top_VIA1 $T=75090 75280 0 0 $X=74840 $Y=75040
X2467 2 digital_ldo_top_VIA1 $T=75090 80720 0 0 $X=74840 $Y=80480
X2468 2 digital_ldo_top_VIA1 $T=75090 86160 0 0 $X=74840 $Y=85920
X2469 2 digital_ldo_top_VIA1 $T=75090 91600 0 0 $X=74840 $Y=91360
X2470 2 digital_ldo_top_VIA1 $T=75090 97040 0 0 $X=74840 $Y=96800
X2471 2 digital_ldo_top_VIA1 $T=75090 102480 0 0 $X=74840 $Y=102240
X2472 2 digital_ldo_top_VIA1 $T=75090 107920 0 0 $X=74840 $Y=107680
X2473 2 digital_ldo_top_VIA1 $T=75090 113360 0 0 $X=74840 $Y=113120
X2474 2 digital_ldo_top_VIA1 $T=75090 118800 0 0 $X=74840 $Y=118560
X2475 2 digital_ldo_top_VIA1 $T=75090 124240 0 0 $X=74840 $Y=124000
X2476 2 digital_ldo_top_VIA1 $T=75090 129680 0 0 $X=74840 $Y=129440
X2477 3 digital_ldo_top_VIA1 $T=77390 12720 0 0 $X=77140 $Y=12480
X2478 3 digital_ldo_top_VIA1 $T=77390 45360 0 0 $X=77140 $Y=45120
X2479 3 digital_ldo_top_VIA1 $T=77390 50800 0 0 $X=77140 $Y=50560
X2480 3 digital_ldo_top_VIA1 $T=77390 56240 0 0 $X=77140 $Y=56000
X2481 3 digital_ldo_top_VIA1 $T=77390 61680 0 0 $X=77140 $Y=61440
X2482 3 digital_ldo_top_VIA1 $T=77390 67120 0 0 $X=77140 $Y=66880
X2483 3 digital_ldo_top_VIA1 $T=77390 72560 0 0 $X=77140 $Y=72320
X2484 3 digital_ldo_top_VIA1 $T=77390 78000 0 0 $X=77140 $Y=77760
X2485 3 digital_ldo_top_VIA1 $T=77390 83440 0 0 $X=77140 $Y=83200
X2486 3 digital_ldo_top_VIA1 $T=77390 88880 0 0 $X=77140 $Y=88640
X2487 3 digital_ldo_top_VIA1 $T=77390 94320 0 0 $X=77140 $Y=94080
X2488 3 digital_ldo_top_VIA1 $T=77390 99760 0 0 $X=77140 $Y=99520
X2489 3 digital_ldo_top_VIA1 $T=77390 105200 0 0 $X=77140 $Y=104960
X2490 3 digital_ldo_top_VIA1 $T=77390 110640 0 0 $X=77140 $Y=110400
X2491 3 digital_ldo_top_VIA1 $T=77390 116080 0 0 $X=77140 $Y=115840
X2492 3 digital_ldo_top_VIA1 $T=77390 121520 0 0 $X=77140 $Y=121280
X2493 3 digital_ldo_top_VIA1 $T=77390 126960 0 0 $X=77140 $Y=126720
X2494 2 digital_ldo_top_VIA1 $T=78770 48080 0 0 $X=78520 $Y=47840
X2495 2 digital_ldo_top_VIA1 $T=78770 53520 0 0 $X=78520 $Y=53280
X2496 2 digital_ldo_top_VIA1 $T=78770 58960 0 0 $X=78520 $Y=58720
X2497 2 digital_ldo_top_VIA1 $T=78770 64400 0 0 $X=78520 $Y=64160
X2498 2 digital_ldo_top_VIA1 $T=78770 69840 0 0 $X=78520 $Y=69600
X2499 2 digital_ldo_top_VIA1 $T=78770 75280 0 0 $X=78520 $Y=75040
X2500 2 digital_ldo_top_VIA1 $T=78770 80720 0 0 $X=78520 $Y=80480
X2501 2 digital_ldo_top_VIA1 $T=78770 86160 0 0 $X=78520 $Y=85920
X2502 2 digital_ldo_top_VIA1 $T=78770 91600 0 0 $X=78520 $Y=91360
X2503 2 digital_ldo_top_VIA1 $T=78770 97040 0 0 $X=78520 $Y=96800
X2504 2 digital_ldo_top_VIA1 $T=78770 102480 0 0 $X=78520 $Y=102240
X2505 2 digital_ldo_top_VIA1 $T=78770 107920 0 0 $X=78520 $Y=107680
X2506 2 digital_ldo_top_VIA1 $T=78770 113360 0 0 $X=78520 $Y=113120
X2507 2 digital_ldo_top_VIA1 $T=78770 118800 0 0 $X=78520 $Y=118560
X2508 2 digital_ldo_top_VIA1 $T=78770 124240 0 0 $X=78520 $Y=124000
X2509 2 digital_ldo_top_VIA1 $T=78770 129680 0 0 $X=78520 $Y=129440
X2510 3 digital_ldo_top_VIA1 $T=81070 12720 0 0 $X=80820 $Y=12480
X2511 3 digital_ldo_top_VIA1 $T=81070 45360 0 0 $X=80820 $Y=45120
X2512 3 digital_ldo_top_VIA1 $T=81070 50800 0 0 $X=80820 $Y=50560
X2513 3 digital_ldo_top_VIA1 $T=81070 56240 0 0 $X=80820 $Y=56000
X2514 3 digital_ldo_top_VIA1 $T=81070 61680 0 0 $X=80820 $Y=61440
X2515 3 digital_ldo_top_VIA1 $T=81070 67120 0 0 $X=80820 $Y=66880
X2516 3 digital_ldo_top_VIA1 $T=81070 72560 0 0 $X=80820 $Y=72320
X2517 3 digital_ldo_top_VIA1 $T=81070 78000 0 0 $X=80820 $Y=77760
X2518 3 digital_ldo_top_VIA1 $T=81070 83440 0 0 $X=80820 $Y=83200
X2519 3 digital_ldo_top_VIA1 $T=81070 88880 0 0 $X=80820 $Y=88640
X2520 3 digital_ldo_top_VIA1 $T=81070 94320 0 0 $X=80820 $Y=94080
X2521 3 digital_ldo_top_VIA1 $T=81070 99760 0 0 $X=80820 $Y=99520
X2522 3 digital_ldo_top_VIA1 $T=81070 105200 0 0 $X=80820 $Y=104960
X2523 3 digital_ldo_top_VIA1 $T=81070 110640 0 0 $X=80820 $Y=110400
X2524 3 digital_ldo_top_VIA1 $T=81070 116080 0 0 $X=80820 $Y=115840
X2525 3 digital_ldo_top_VIA1 $T=81070 121520 0 0 $X=80820 $Y=121280
X2526 3 digital_ldo_top_VIA1 $T=81070 126960 0 0 $X=80820 $Y=126720
X2527 2 digital_ldo_top_VIA1 $T=82450 48080 0 0 $X=82200 $Y=47840
X2528 2 digital_ldo_top_VIA1 $T=82450 53520 0 0 $X=82200 $Y=53280
X2529 2 digital_ldo_top_VIA1 $T=82450 58960 0 0 $X=82200 $Y=58720
X2530 2 digital_ldo_top_VIA1 $T=82450 64400 0 0 $X=82200 $Y=64160
X2531 2 digital_ldo_top_VIA1 $T=82450 69840 0 0 $X=82200 $Y=69600
X2532 2 digital_ldo_top_VIA1 $T=82450 75280 0 0 $X=82200 $Y=75040
X2533 2 digital_ldo_top_VIA1 $T=82450 80720 0 0 $X=82200 $Y=80480
X2534 2 digital_ldo_top_VIA1 $T=82450 86160 0 0 $X=82200 $Y=85920
X2535 2 digital_ldo_top_VIA1 $T=82450 91600 0 0 $X=82200 $Y=91360
X2536 2 digital_ldo_top_VIA1 $T=82450 97040 0 0 $X=82200 $Y=96800
X2537 2 digital_ldo_top_VIA1 $T=82450 102480 0 0 $X=82200 $Y=102240
X2538 2 digital_ldo_top_VIA1 $T=82450 107920 0 0 $X=82200 $Y=107680
X2539 2 digital_ldo_top_VIA1 $T=82450 113360 0 0 $X=82200 $Y=113120
X2540 2 digital_ldo_top_VIA1 $T=82450 118800 0 0 $X=82200 $Y=118560
X2541 2 digital_ldo_top_VIA1 $T=82450 124240 0 0 $X=82200 $Y=124000
X2542 2 digital_ldo_top_VIA1 $T=82450 129680 0 0 $X=82200 $Y=129440
X2543 3 digital_ldo_top_VIA1 $T=84750 12720 0 0 $X=84500 $Y=12480
X2544 3 digital_ldo_top_VIA1 $T=84750 45360 0 0 $X=84500 $Y=45120
X2545 3 digital_ldo_top_VIA1 $T=84750 50800 0 0 $X=84500 $Y=50560
X2546 3 digital_ldo_top_VIA1 $T=84750 56240 0 0 $X=84500 $Y=56000
X2547 3 digital_ldo_top_VIA1 $T=84750 61680 0 0 $X=84500 $Y=61440
X2548 3 digital_ldo_top_VIA1 $T=84750 67120 0 0 $X=84500 $Y=66880
X2549 3 digital_ldo_top_VIA1 $T=84750 72560 0 0 $X=84500 $Y=72320
X2550 3 digital_ldo_top_VIA1 $T=84750 78000 0 0 $X=84500 $Y=77760
X2551 3 digital_ldo_top_VIA1 $T=84750 83440 0 0 $X=84500 $Y=83200
X2552 3 digital_ldo_top_VIA1 $T=84750 88880 0 0 $X=84500 $Y=88640
X2553 3 digital_ldo_top_VIA1 $T=84750 94320 0 0 $X=84500 $Y=94080
X2554 3 digital_ldo_top_VIA1 $T=84750 99760 0 0 $X=84500 $Y=99520
X2555 3 digital_ldo_top_VIA1 $T=84750 105200 0 0 $X=84500 $Y=104960
X2556 3 digital_ldo_top_VIA1 $T=84750 110640 0 0 $X=84500 $Y=110400
X2557 3 digital_ldo_top_VIA1 $T=84750 116080 0 0 $X=84500 $Y=115840
X2558 3 digital_ldo_top_VIA1 $T=84750 121520 0 0 $X=84500 $Y=121280
X2559 3 digital_ldo_top_VIA1 $T=84750 126960 0 0 $X=84500 $Y=126720
X2560 2 digital_ldo_top_VIA1 $T=86130 48080 0 0 $X=85880 $Y=47840
X2561 2 digital_ldo_top_VIA1 $T=86130 53520 0 0 $X=85880 $Y=53280
X2562 2 digital_ldo_top_VIA1 $T=86130 58960 0 0 $X=85880 $Y=58720
X2563 2 digital_ldo_top_VIA1 $T=86130 64400 0 0 $X=85880 $Y=64160
X2564 2 digital_ldo_top_VIA1 $T=86130 69840 0 0 $X=85880 $Y=69600
X2565 2 digital_ldo_top_VIA1 $T=86130 75280 0 0 $X=85880 $Y=75040
X2566 2 digital_ldo_top_VIA1 $T=86130 80720 0 0 $X=85880 $Y=80480
X2567 2 digital_ldo_top_VIA1 $T=86130 86160 0 0 $X=85880 $Y=85920
X2568 2 digital_ldo_top_VIA1 $T=86130 91600 0 0 $X=85880 $Y=91360
X2569 2 digital_ldo_top_VIA1 $T=86130 97040 0 0 $X=85880 $Y=96800
X2570 2 digital_ldo_top_VIA1 $T=86130 102480 0 0 $X=85880 $Y=102240
X2571 2 digital_ldo_top_VIA1 $T=86130 107920 0 0 $X=85880 $Y=107680
X2572 2 digital_ldo_top_VIA1 $T=86130 113360 0 0 $X=85880 $Y=113120
X2573 2 digital_ldo_top_VIA1 $T=86130 118800 0 0 $X=85880 $Y=118560
X2574 2 digital_ldo_top_VIA1 $T=86130 124240 0 0 $X=85880 $Y=124000
X2575 2 digital_ldo_top_VIA1 $T=86130 129680 0 0 $X=85880 $Y=129440
X2576 3 digital_ldo_top_VIA1 $T=88430 12720 0 0 $X=88180 $Y=12480
X2577 3 digital_ldo_top_VIA1 $T=88430 45360 0 0 $X=88180 $Y=45120
X2578 3 digital_ldo_top_VIA1 $T=88430 50800 0 0 $X=88180 $Y=50560
X2579 3 digital_ldo_top_VIA1 $T=88430 56240 0 0 $X=88180 $Y=56000
X2580 3 digital_ldo_top_VIA1 $T=88430 61680 0 0 $X=88180 $Y=61440
X2581 3 digital_ldo_top_VIA1 $T=88430 67120 0 0 $X=88180 $Y=66880
X2582 3 digital_ldo_top_VIA1 $T=88430 72560 0 0 $X=88180 $Y=72320
X2583 3 digital_ldo_top_VIA1 $T=88430 78000 0 0 $X=88180 $Y=77760
X2584 3 digital_ldo_top_VIA1 $T=88430 83440 0 0 $X=88180 $Y=83200
X2585 3 digital_ldo_top_VIA1 $T=88430 88880 0 0 $X=88180 $Y=88640
X2586 3 digital_ldo_top_VIA1 $T=88430 94320 0 0 $X=88180 $Y=94080
X2587 3 digital_ldo_top_VIA1 $T=88430 99760 0 0 $X=88180 $Y=99520
X2588 3 digital_ldo_top_VIA1 $T=88430 105200 0 0 $X=88180 $Y=104960
X2589 3 digital_ldo_top_VIA1 $T=88430 110640 0 0 $X=88180 $Y=110400
X2590 3 digital_ldo_top_VIA1 $T=88430 116080 0 0 $X=88180 $Y=115840
X2591 3 digital_ldo_top_VIA1 $T=88430 121520 0 0 $X=88180 $Y=121280
X2592 3 digital_ldo_top_VIA1 $T=88430 126960 0 0 $X=88180 $Y=126720
X2593 2 digital_ldo_top_VIA1 $T=89810 48080 0 0 $X=89560 $Y=47840
X2594 2 digital_ldo_top_VIA1 $T=89810 53520 0 0 $X=89560 $Y=53280
X2595 2 digital_ldo_top_VIA1 $T=89810 58960 0 0 $X=89560 $Y=58720
X2596 2 digital_ldo_top_VIA1 $T=89810 64400 0 0 $X=89560 $Y=64160
X2597 2 digital_ldo_top_VIA1 $T=89810 69840 0 0 $X=89560 $Y=69600
X2598 2 digital_ldo_top_VIA1 $T=89810 75280 0 0 $X=89560 $Y=75040
X2599 2 digital_ldo_top_VIA1 $T=89810 80720 0 0 $X=89560 $Y=80480
X2600 2 digital_ldo_top_VIA1 $T=89810 86160 0 0 $X=89560 $Y=85920
X2601 2 digital_ldo_top_VIA1 $T=89810 91600 0 0 $X=89560 $Y=91360
X2602 2 digital_ldo_top_VIA1 $T=89810 97040 0 0 $X=89560 $Y=96800
X2603 2 digital_ldo_top_VIA1 $T=89810 102480 0 0 $X=89560 $Y=102240
X2604 2 digital_ldo_top_VIA1 $T=89810 107920 0 0 $X=89560 $Y=107680
X2605 2 digital_ldo_top_VIA1 $T=89810 113360 0 0 $X=89560 $Y=113120
X2606 2 digital_ldo_top_VIA1 $T=89810 118800 0 0 $X=89560 $Y=118560
X2607 2 digital_ldo_top_VIA1 $T=89810 124240 0 0 $X=89560 $Y=124000
X2608 2 digital_ldo_top_VIA1 $T=89810 129680 0 0 $X=89560 $Y=129440
X2609 3 digital_ldo_top_VIA1 $T=92110 12720 0 0 $X=91860 $Y=12480
X2610 3 digital_ldo_top_VIA1 $T=92110 18160 0 0 $X=91860 $Y=17920
X2611 3 digital_ldo_top_VIA1 $T=92110 23600 0 0 $X=91860 $Y=23360
X2612 3 digital_ldo_top_VIA1 $T=92110 29040 0 0 $X=91860 $Y=28800
X2613 3 digital_ldo_top_VIA1 $T=92110 34480 0 0 $X=91860 $Y=34240
X2614 3 digital_ldo_top_VIA1 $T=92110 39920 0 0 $X=91860 $Y=39680
X2615 3 digital_ldo_top_VIA1 $T=92110 45360 0 0 $X=91860 $Y=45120
X2616 3 digital_ldo_top_VIA1 $T=92110 50800 0 0 $X=91860 $Y=50560
X2617 3 digital_ldo_top_VIA1 $T=92110 56240 0 0 $X=91860 $Y=56000
X2618 3 digital_ldo_top_VIA1 $T=92110 61680 0 0 $X=91860 $Y=61440
X2619 3 digital_ldo_top_VIA1 $T=92110 67120 0 0 $X=91860 $Y=66880
X2620 3 digital_ldo_top_VIA1 $T=92110 72560 0 0 $X=91860 $Y=72320
X2621 3 digital_ldo_top_VIA1 $T=92110 78000 0 0 $X=91860 $Y=77760
X2622 3 digital_ldo_top_VIA1 $T=92110 83440 0 0 $X=91860 $Y=83200
X2623 3 digital_ldo_top_VIA1 $T=92110 88880 0 0 $X=91860 $Y=88640
X2624 3 digital_ldo_top_VIA1 $T=92110 94320 0 0 $X=91860 $Y=94080
X2625 3 digital_ldo_top_VIA1 $T=92110 99760 0 0 $X=91860 $Y=99520
X2626 3 digital_ldo_top_VIA1 $T=92110 105200 0 0 $X=91860 $Y=104960
X2627 3 digital_ldo_top_VIA1 $T=92110 110640 0 0 $X=91860 $Y=110400
X2628 3 digital_ldo_top_VIA1 $T=92110 116080 0 0 $X=91860 $Y=115840
X2629 3 digital_ldo_top_VIA1 $T=92110 121520 0 0 $X=91860 $Y=121280
X2630 3 digital_ldo_top_VIA1 $T=92110 126960 0 0 $X=91860 $Y=126720
X2631 2 digital_ldo_top_VIA1 $T=93490 15440 0 0 $X=93240 $Y=15200
X2632 2 digital_ldo_top_VIA1 $T=93490 20880 0 0 $X=93240 $Y=20640
X2633 2 digital_ldo_top_VIA1 $T=93490 26320 0 0 $X=93240 $Y=26080
X2634 2 digital_ldo_top_VIA1 $T=93490 31760 0 0 $X=93240 $Y=31520
X2635 2 digital_ldo_top_VIA1 $T=93490 37200 0 0 $X=93240 $Y=36960
X2636 2 digital_ldo_top_VIA1 $T=93490 42640 0 0 $X=93240 $Y=42400
X2637 2 digital_ldo_top_VIA1 $T=93490 48080 0 0 $X=93240 $Y=47840
X2638 2 digital_ldo_top_VIA1 $T=93490 53520 0 0 $X=93240 $Y=53280
X2639 2 digital_ldo_top_VIA1 $T=93490 58960 0 0 $X=93240 $Y=58720
X2640 2 digital_ldo_top_VIA1 $T=93490 64400 0 0 $X=93240 $Y=64160
X2641 2 digital_ldo_top_VIA1 $T=93490 69840 0 0 $X=93240 $Y=69600
X2642 2 digital_ldo_top_VIA1 $T=93490 75280 0 0 $X=93240 $Y=75040
X2643 2 digital_ldo_top_VIA1 $T=93490 80720 0 0 $X=93240 $Y=80480
X2644 2 digital_ldo_top_VIA1 $T=93490 86160 0 0 $X=93240 $Y=85920
X2645 2 digital_ldo_top_VIA1 $T=93490 91600 0 0 $X=93240 $Y=91360
X2646 2 digital_ldo_top_VIA1 $T=93490 97040 0 0 $X=93240 $Y=96800
X2647 2 digital_ldo_top_VIA1 $T=93490 102480 0 0 $X=93240 $Y=102240
X2648 2 digital_ldo_top_VIA1 $T=93490 107920 0 0 $X=93240 $Y=107680
X2649 2 digital_ldo_top_VIA1 $T=93490 113360 0 0 $X=93240 $Y=113120
X2650 2 digital_ldo_top_VIA1 $T=93490 118800 0 0 $X=93240 $Y=118560
X2651 2 digital_ldo_top_VIA1 $T=93490 124240 0 0 $X=93240 $Y=124000
X2652 2 digital_ldo_top_VIA1 $T=93490 129680 0 0 $X=93240 $Y=129440
X2653 3 digital_ldo_top_VIA1 $T=95790 12720 0 0 $X=95540 $Y=12480
X2654 3 digital_ldo_top_VIA1 $T=95790 18160 0 0 $X=95540 $Y=17920
X2655 3 digital_ldo_top_VIA1 $T=95790 23600 0 0 $X=95540 $Y=23360
X2656 3 digital_ldo_top_VIA1 $T=95790 29040 0 0 $X=95540 $Y=28800
X2657 3 digital_ldo_top_VIA1 $T=95790 34480 0 0 $X=95540 $Y=34240
X2658 3 digital_ldo_top_VIA1 $T=95790 39920 0 0 $X=95540 $Y=39680
X2659 3 digital_ldo_top_VIA1 $T=95790 45360 0 0 $X=95540 $Y=45120
X2660 3 digital_ldo_top_VIA1 $T=95790 50800 0 0 $X=95540 $Y=50560
X2661 3 digital_ldo_top_VIA1 $T=95790 56240 0 0 $X=95540 $Y=56000
X2662 3 digital_ldo_top_VIA1 $T=95790 61680 0 0 $X=95540 $Y=61440
X2663 3 digital_ldo_top_VIA1 $T=95790 67120 0 0 $X=95540 $Y=66880
X2664 3 digital_ldo_top_VIA1 $T=95790 72560 0 0 $X=95540 $Y=72320
X2665 3 digital_ldo_top_VIA1 $T=95790 78000 0 0 $X=95540 $Y=77760
X2666 3 digital_ldo_top_VIA1 $T=95790 83440 0 0 $X=95540 $Y=83200
X2667 3 digital_ldo_top_VIA1 $T=95790 88880 0 0 $X=95540 $Y=88640
X2668 3 digital_ldo_top_VIA1 $T=95790 94320 0 0 $X=95540 $Y=94080
X2669 3 digital_ldo_top_VIA1 $T=95790 99760 0 0 $X=95540 $Y=99520
X2670 3 digital_ldo_top_VIA1 $T=95790 105200 0 0 $X=95540 $Y=104960
X2671 3 digital_ldo_top_VIA1 $T=95790 110640 0 0 $X=95540 $Y=110400
X2672 3 digital_ldo_top_VIA1 $T=95790 116080 0 0 $X=95540 $Y=115840
X2673 3 digital_ldo_top_VIA1 $T=95790 121520 0 0 $X=95540 $Y=121280
X2674 3 digital_ldo_top_VIA1 $T=95790 126960 0 0 $X=95540 $Y=126720
X2675 2 digital_ldo_top_VIA1 $T=97170 15440 0 0 $X=96920 $Y=15200
X2676 2 digital_ldo_top_VIA1 $T=97170 20880 0 0 $X=96920 $Y=20640
X2677 2 digital_ldo_top_VIA1 $T=97170 26320 0 0 $X=96920 $Y=26080
X2678 2 digital_ldo_top_VIA1 $T=97170 31760 0 0 $X=96920 $Y=31520
X2679 2 digital_ldo_top_VIA1 $T=97170 37200 0 0 $X=96920 $Y=36960
X2680 2 digital_ldo_top_VIA1 $T=97170 42640 0 0 $X=96920 $Y=42400
X2681 2 digital_ldo_top_VIA1 $T=97170 48080 0 0 $X=96920 $Y=47840
X2682 2 digital_ldo_top_VIA1 $T=97170 53520 0 0 $X=96920 $Y=53280
X2683 2 digital_ldo_top_VIA1 $T=97170 58960 0 0 $X=96920 $Y=58720
X2684 2 digital_ldo_top_VIA1 $T=97170 64400 0 0 $X=96920 $Y=64160
X2685 2 digital_ldo_top_VIA1 $T=97170 69840 0 0 $X=96920 $Y=69600
X2686 2 digital_ldo_top_VIA1 $T=97170 75280 0 0 $X=96920 $Y=75040
X2687 2 digital_ldo_top_VIA1 $T=97170 80720 0 0 $X=96920 $Y=80480
X2688 2 digital_ldo_top_VIA1 $T=97170 86160 0 0 $X=96920 $Y=85920
X2689 2 digital_ldo_top_VIA1 $T=97170 91600 0 0 $X=96920 $Y=91360
X2690 2 digital_ldo_top_VIA1 $T=97170 97040 0 0 $X=96920 $Y=96800
X2691 2 digital_ldo_top_VIA1 $T=97170 102480 0 0 $X=96920 $Y=102240
X2692 2 digital_ldo_top_VIA1 $T=97170 107920 0 0 $X=96920 $Y=107680
X2693 2 digital_ldo_top_VIA1 $T=97170 113360 0 0 $X=96920 $Y=113120
X2694 2 digital_ldo_top_VIA1 $T=97170 118800 0 0 $X=96920 $Y=118560
X2695 2 digital_ldo_top_VIA1 $T=97170 124240 0 0 $X=96920 $Y=124000
X2696 2 digital_ldo_top_VIA1 $T=97170 129680 0 0 $X=96920 $Y=129440
X2697 3 digital_ldo_top_VIA1 $T=99470 12720 0 0 $X=99220 $Y=12480
X2698 3 digital_ldo_top_VIA1 $T=99470 18160 0 0 $X=99220 $Y=17920
X2699 3 digital_ldo_top_VIA1 $T=99470 23600 0 0 $X=99220 $Y=23360
X2700 3 digital_ldo_top_VIA1 $T=99470 29040 0 0 $X=99220 $Y=28800
X2701 3 digital_ldo_top_VIA1 $T=99470 34480 0 0 $X=99220 $Y=34240
X2702 3 digital_ldo_top_VIA1 $T=99470 39920 0 0 $X=99220 $Y=39680
X2703 3 digital_ldo_top_VIA1 $T=99470 45360 0 0 $X=99220 $Y=45120
X2704 3 digital_ldo_top_VIA1 $T=99470 50800 0 0 $X=99220 $Y=50560
X2705 3 digital_ldo_top_VIA1 $T=99470 56240 0 0 $X=99220 $Y=56000
X2706 3 digital_ldo_top_VIA1 $T=99470 61680 0 0 $X=99220 $Y=61440
X2707 3 digital_ldo_top_VIA1 $T=99470 67120 0 0 $X=99220 $Y=66880
X2708 3 digital_ldo_top_VIA1 $T=99470 72560 0 0 $X=99220 $Y=72320
X2709 3 digital_ldo_top_VIA1 $T=99470 78000 0 0 $X=99220 $Y=77760
X2710 3 digital_ldo_top_VIA1 $T=99470 83440 0 0 $X=99220 $Y=83200
X2711 3 digital_ldo_top_VIA1 $T=99470 88880 0 0 $X=99220 $Y=88640
X2712 3 digital_ldo_top_VIA1 $T=99470 94320 0 0 $X=99220 $Y=94080
X2713 3 digital_ldo_top_VIA1 $T=99470 99760 0 0 $X=99220 $Y=99520
X2714 3 digital_ldo_top_VIA1 $T=99470 105200 0 0 $X=99220 $Y=104960
X2715 3 digital_ldo_top_VIA1 $T=99470 110640 0 0 $X=99220 $Y=110400
X2716 3 digital_ldo_top_VIA1 $T=99470 116080 0 0 $X=99220 $Y=115840
X2717 3 digital_ldo_top_VIA1 $T=99470 121520 0 0 $X=99220 $Y=121280
X2718 3 digital_ldo_top_VIA1 $T=99470 126960 0 0 $X=99220 $Y=126720
X2719 2 digital_ldo_top_VIA1 $T=100850 15440 0 0 $X=100600 $Y=15200
X2720 2 digital_ldo_top_VIA1 $T=100850 20880 0 0 $X=100600 $Y=20640
X2721 2 digital_ldo_top_VIA1 $T=100850 26320 0 0 $X=100600 $Y=26080
X2722 2 digital_ldo_top_VIA1 $T=100850 31760 0 0 $X=100600 $Y=31520
X2723 2 digital_ldo_top_VIA1 $T=100850 37200 0 0 $X=100600 $Y=36960
X2724 2 digital_ldo_top_VIA1 $T=100850 42640 0 0 $X=100600 $Y=42400
X2725 2 digital_ldo_top_VIA1 $T=100850 48080 0 0 $X=100600 $Y=47840
X2726 2 digital_ldo_top_VIA1 $T=100850 53520 0 0 $X=100600 $Y=53280
X2727 2 digital_ldo_top_VIA1 $T=100850 58960 0 0 $X=100600 $Y=58720
X2728 2 digital_ldo_top_VIA1 $T=100850 64400 0 0 $X=100600 $Y=64160
X2729 2 digital_ldo_top_VIA1 $T=100850 69840 0 0 $X=100600 $Y=69600
X2730 2 digital_ldo_top_VIA1 $T=100850 75280 0 0 $X=100600 $Y=75040
X2731 2 digital_ldo_top_VIA1 $T=100850 80720 0 0 $X=100600 $Y=80480
X2732 2 digital_ldo_top_VIA1 $T=100850 86160 0 0 $X=100600 $Y=85920
X2733 2 digital_ldo_top_VIA1 $T=100850 91600 0 0 $X=100600 $Y=91360
X2734 2 digital_ldo_top_VIA1 $T=100850 97040 0 0 $X=100600 $Y=96800
X2735 2 digital_ldo_top_VIA1 $T=100850 102480 0 0 $X=100600 $Y=102240
X2736 2 digital_ldo_top_VIA1 $T=100850 107920 0 0 $X=100600 $Y=107680
X2737 2 digital_ldo_top_VIA1 $T=100850 113360 0 0 $X=100600 $Y=113120
X2738 2 digital_ldo_top_VIA1 $T=100850 118800 0 0 $X=100600 $Y=118560
X2739 2 digital_ldo_top_VIA1 $T=100850 124240 0 0 $X=100600 $Y=124000
X2740 2 digital_ldo_top_VIA1 $T=100850 129680 0 0 $X=100600 $Y=129440
X2741 3 digital_ldo_top_VIA1 $T=103150 12720 0 0 $X=102900 $Y=12480
X2742 3 digital_ldo_top_VIA1 $T=103150 18160 0 0 $X=102900 $Y=17920
X2743 3 digital_ldo_top_VIA1 $T=103150 94320 0 0 $X=102900 $Y=94080
X2744 3 digital_ldo_top_VIA1 $T=103150 99760 0 0 $X=102900 $Y=99520
X2745 3 digital_ldo_top_VIA1 $T=103150 105200 0 0 $X=102900 $Y=104960
X2746 3 digital_ldo_top_VIA1 $T=103150 110640 0 0 $X=102900 $Y=110400
X2747 3 digital_ldo_top_VIA1 $T=103150 116080 0 0 $X=102900 $Y=115840
X2748 3 digital_ldo_top_VIA1 $T=103150 121520 0 0 $X=102900 $Y=121280
X2749 3 digital_ldo_top_VIA1 $T=103150 126960 0 0 $X=102900 $Y=126720
X2750 2 digital_ldo_top_VIA1 $T=104530 15440 0 0 $X=104280 $Y=15200
X2751 2 digital_ldo_top_VIA1 $T=104530 91600 0 0 $X=104280 $Y=91360
X2752 2 digital_ldo_top_VIA1 $T=104530 97040 0 0 $X=104280 $Y=96800
X2753 2 digital_ldo_top_VIA1 $T=104530 102480 0 0 $X=104280 $Y=102240
X2754 2 digital_ldo_top_VIA1 $T=104530 107920 0 0 $X=104280 $Y=107680
X2755 2 digital_ldo_top_VIA1 $T=104530 113360 0 0 $X=104280 $Y=113120
X2756 2 digital_ldo_top_VIA1 $T=104530 118800 0 0 $X=104280 $Y=118560
X2757 2 digital_ldo_top_VIA1 $T=104530 124240 0 0 $X=104280 $Y=124000
X2758 2 digital_ldo_top_VIA1 $T=104530 129680 0 0 $X=104280 $Y=129440
X2759 3 digital_ldo_top_VIA1 $T=106830 12720 0 0 $X=106580 $Y=12480
X2760 3 digital_ldo_top_VIA1 $T=106830 18160 0 0 $X=106580 $Y=17920
X2761 3 digital_ldo_top_VIA1 $T=106830 94320 0 0 $X=106580 $Y=94080
X2762 3 digital_ldo_top_VIA1 $T=106830 99760 0 0 $X=106580 $Y=99520
X2763 3 digital_ldo_top_VIA1 $T=106830 105200 0 0 $X=106580 $Y=104960
X2764 3 digital_ldo_top_VIA1 $T=106830 110640 0 0 $X=106580 $Y=110400
X2765 3 digital_ldo_top_VIA1 $T=106830 116080 0 0 $X=106580 $Y=115840
X2766 3 digital_ldo_top_VIA1 $T=106830 121520 0 0 $X=106580 $Y=121280
X2767 3 digital_ldo_top_VIA1 $T=106830 126960 0 0 $X=106580 $Y=126720
X2768 2 digital_ldo_top_VIA1 $T=108210 15440 0 0 $X=107960 $Y=15200
X2769 2 digital_ldo_top_VIA1 $T=108210 91600 0 0 $X=107960 $Y=91360
X2770 2 digital_ldo_top_VIA1 $T=108210 97040 0 0 $X=107960 $Y=96800
X2771 2 digital_ldo_top_VIA1 $T=108210 102480 0 0 $X=107960 $Y=102240
X2772 2 digital_ldo_top_VIA1 $T=108210 107920 0 0 $X=107960 $Y=107680
X2773 2 digital_ldo_top_VIA1 $T=108210 113360 0 0 $X=107960 $Y=113120
X2774 2 digital_ldo_top_VIA1 $T=108210 118800 0 0 $X=107960 $Y=118560
X2775 2 digital_ldo_top_VIA1 $T=108210 124240 0 0 $X=107960 $Y=124000
X2776 2 digital_ldo_top_VIA1 $T=108210 129680 0 0 $X=107960 $Y=129440
X2777 3 digital_ldo_top_VIA1 $T=110510 12720 0 0 $X=110260 $Y=12480
X2778 3 digital_ldo_top_VIA1 $T=110510 18160 0 0 $X=110260 $Y=17920
X2779 3 digital_ldo_top_VIA1 $T=110510 94320 0 0 $X=110260 $Y=94080
X2780 3 digital_ldo_top_VIA1 $T=110510 99760 0 0 $X=110260 $Y=99520
X2781 3 digital_ldo_top_VIA1 $T=110510 105200 0 0 $X=110260 $Y=104960
X2782 3 digital_ldo_top_VIA1 $T=110510 110640 0 0 $X=110260 $Y=110400
X2783 3 digital_ldo_top_VIA1 $T=110510 116080 0 0 $X=110260 $Y=115840
X2784 3 digital_ldo_top_VIA1 $T=110510 121520 0 0 $X=110260 $Y=121280
X2785 3 digital_ldo_top_VIA1 $T=110510 126960 0 0 $X=110260 $Y=126720
X2786 2 digital_ldo_top_VIA1 $T=111890 15440 0 0 $X=111640 $Y=15200
X2787 2 digital_ldo_top_VIA1 $T=111890 91600 0 0 $X=111640 $Y=91360
X2788 2 digital_ldo_top_VIA1 $T=111890 97040 0 0 $X=111640 $Y=96800
X2789 2 digital_ldo_top_VIA1 $T=111890 102480 0 0 $X=111640 $Y=102240
X2790 2 digital_ldo_top_VIA1 $T=111890 107920 0 0 $X=111640 $Y=107680
X2791 2 digital_ldo_top_VIA1 $T=111890 113360 0 0 $X=111640 $Y=113120
X2792 2 digital_ldo_top_VIA1 $T=111890 118800 0 0 $X=111640 $Y=118560
X2793 2 digital_ldo_top_VIA1 $T=111890 124240 0 0 $X=111640 $Y=124000
X2794 2 digital_ldo_top_VIA1 $T=111890 129680 0 0 $X=111640 $Y=129440
X2795 3 digital_ldo_top_VIA1 $T=114190 12720 0 0 $X=113940 $Y=12480
X2796 3 digital_ldo_top_VIA1 $T=114190 18160 0 0 $X=113940 $Y=17920
X2797 3 digital_ldo_top_VIA1 $T=114190 94320 0 0 $X=113940 $Y=94080
X2798 3 digital_ldo_top_VIA1 $T=114190 99760 0 0 $X=113940 $Y=99520
X2799 3 digital_ldo_top_VIA1 $T=114190 105200 0 0 $X=113940 $Y=104960
X2800 3 digital_ldo_top_VIA1 $T=114190 110640 0 0 $X=113940 $Y=110400
X2801 3 digital_ldo_top_VIA1 $T=114190 116080 0 0 $X=113940 $Y=115840
X2802 3 digital_ldo_top_VIA1 $T=114190 121520 0 0 $X=113940 $Y=121280
X2803 3 digital_ldo_top_VIA1 $T=114190 126960 0 0 $X=113940 $Y=126720
X2804 2 digital_ldo_top_VIA1 $T=115570 15440 0 0 $X=115320 $Y=15200
X2805 2 digital_ldo_top_VIA1 $T=115570 91600 0 0 $X=115320 $Y=91360
X2806 2 digital_ldo_top_VIA1 $T=115570 97040 0 0 $X=115320 $Y=96800
X2807 2 digital_ldo_top_VIA1 $T=115570 102480 0 0 $X=115320 $Y=102240
X2808 2 digital_ldo_top_VIA1 $T=115570 107920 0 0 $X=115320 $Y=107680
X2809 2 digital_ldo_top_VIA1 $T=115570 113360 0 0 $X=115320 $Y=113120
X2810 2 digital_ldo_top_VIA1 $T=115570 118800 0 0 $X=115320 $Y=118560
X2811 2 digital_ldo_top_VIA1 $T=115570 124240 0 0 $X=115320 $Y=124000
X2812 2 digital_ldo_top_VIA1 $T=115570 129680 0 0 $X=115320 $Y=129440
X2813 3 digital_ldo_top_VIA1 $T=117870 12720 0 0 $X=117620 $Y=12480
X2814 3 digital_ldo_top_VIA1 $T=117870 18160 0 0 $X=117620 $Y=17920
X2815 3 digital_ldo_top_VIA1 $T=117870 37720 0 0 $X=117620 $Y=37480
X2816 3 digital_ldo_top_VIA1 $T=117870 43160 0 0 $X=117620 $Y=42920
X2817 3 digital_ldo_top_VIA1 $T=117870 48600 0 0 $X=117620 $Y=48360
X2818 3 digital_ldo_top_VIA1 $T=117870 54040 0 0 $X=117620 $Y=53800
X2819 3 digital_ldo_top_VIA1 $T=117870 59480 0 0 $X=117620 $Y=59240
X2820 3 digital_ldo_top_VIA1 $T=117870 64920 0 0 $X=117620 $Y=64680
X2821 3 digital_ldo_top_VIA1 $T=117870 70360 0 0 $X=117620 $Y=70120
X2822 3 digital_ldo_top_VIA1 $T=117870 75800 0 0 $X=117620 $Y=75560
X2823 3 digital_ldo_top_VIA1 $T=117870 81240 0 0 $X=117620 $Y=81000
X2824 3 digital_ldo_top_VIA1 $T=117870 94320 0 0 $X=117620 $Y=94080
X2825 3 digital_ldo_top_VIA1 $T=117870 99760 0 0 $X=117620 $Y=99520
X2826 3 digital_ldo_top_VIA1 $T=117870 105200 0 0 $X=117620 $Y=104960
X2827 3 digital_ldo_top_VIA1 $T=117870 110640 0 0 $X=117620 $Y=110400
X2828 3 digital_ldo_top_VIA1 $T=117870 116080 0 0 $X=117620 $Y=115840
X2829 3 digital_ldo_top_VIA1 $T=117870 121520 0 0 $X=117620 $Y=121280
X2830 3 digital_ldo_top_VIA1 $T=117870 126960 0 0 $X=117620 $Y=126720
X2831 2 digital_ldo_top_VIA1 $T=119250 15440 0 0 $X=119000 $Y=15200
X2832 2 digital_ldo_top_VIA1 $T=119250 91600 0 0 $X=119000 $Y=91360
X2833 2 digital_ldo_top_VIA1 $T=119250 97040 0 0 $X=119000 $Y=96800
X2834 2 digital_ldo_top_VIA1 $T=119250 102480 0 0 $X=119000 $Y=102240
X2835 2 digital_ldo_top_VIA1 $T=119250 107920 0 0 $X=119000 $Y=107680
X2836 2 digital_ldo_top_VIA1 $T=119250 113360 0 0 $X=119000 $Y=113120
X2837 2 digital_ldo_top_VIA1 $T=119250 118800 0 0 $X=119000 $Y=118560
X2838 2 digital_ldo_top_VIA1 $T=119250 124240 0 0 $X=119000 $Y=124000
X2839 2 digital_ldo_top_VIA1 $T=119250 129680 0 0 $X=119000 $Y=129440
X2840 3 digital_ldo_top_VIA1 $T=121550 12720 0 0 $X=121300 $Y=12480
X2841 3 digital_ldo_top_VIA1 $T=121550 18160 0 0 $X=121300 $Y=17920
X2842 3 digital_ldo_top_VIA1 $T=121550 94320 0 0 $X=121300 $Y=94080
X2843 3 digital_ldo_top_VIA1 $T=121550 99760 0 0 $X=121300 $Y=99520
X2844 3 digital_ldo_top_VIA1 $T=121550 105200 0 0 $X=121300 $Y=104960
X2845 3 digital_ldo_top_VIA1 $T=121550 110640 0 0 $X=121300 $Y=110400
X2846 3 digital_ldo_top_VIA1 $T=121550 116080 0 0 $X=121300 $Y=115840
X2847 3 digital_ldo_top_VIA1 $T=121550 121520 0 0 $X=121300 $Y=121280
X2848 3 digital_ldo_top_VIA1 $T=121550 126960 0 0 $X=121300 $Y=126720
X2849 2 digital_ldo_top_VIA1 $T=122930 15440 0 0 $X=122680 $Y=15200
X2850 2 digital_ldo_top_VIA1 $T=122930 35000 0 0 $X=122680 $Y=34760
X2851 2 digital_ldo_top_VIA1 $T=122930 40440 0 0 $X=122680 $Y=40200
X2852 2 digital_ldo_top_VIA1 $T=122930 45880 0 0 $X=122680 $Y=45640
X2853 2 digital_ldo_top_VIA1 $T=122930 51320 0 0 $X=122680 $Y=51080
X2854 2 digital_ldo_top_VIA1 $T=122930 56760 0 0 $X=122680 $Y=56520
X2855 2 digital_ldo_top_VIA1 $T=122930 62200 0 0 $X=122680 $Y=61960
X2856 2 digital_ldo_top_VIA1 $T=122930 67640 0 0 $X=122680 $Y=67400
X2857 2 digital_ldo_top_VIA1 $T=122930 73080 0 0 $X=122680 $Y=72840
X2858 2 digital_ldo_top_VIA1 $T=122930 78520 0 0 $X=122680 $Y=78280
X2859 2 digital_ldo_top_VIA1 $T=122930 83960 0 0 $X=122680 $Y=83720
X2860 2 digital_ldo_top_VIA1 $T=122930 91600 0 0 $X=122680 $Y=91360
X2861 2 digital_ldo_top_VIA1 $T=122930 97040 0 0 $X=122680 $Y=96800
X2862 2 digital_ldo_top_VIA1 $T=122930 102480 0 0 $X=122680 $Y=102240
X2863 2 digital_ldo_top_VIA1 $T=122930 107920 0 0 $X=122680 $Y=107680
X2864 2 digital_ldo_top_VIA1 $T=122930 113360 0 0 $X=122680 $Y=113120
X2865 2 digital_ldo_top_VIA1 $T=122930 118800 0 0 $X=122680 $Y=118560
X2866 2 digital_ldo_top_VIA1 $T=122930 124240 0 0 $X=122680 $Y=124000
X2867 2 digital_ldo_top_VIA1 $T=122930 129680 0 0 $X=122680 $Y=129440
X2868 3 digital_ldo_top_VIA1 $T=125230 12720 0 0 $X=124980 $Y=12480
X2869 3 digital_ldo_top_VIA1 $T=125230 18160 0 0 $X=124980 $Y=17920
X2870 3 digital_ldo_top_VIA1 $T=125230 94320 0 0 $X=124980 $Y=94080
X2871 3 digital_ldo_top_VIA1 $T=125230 99760 0 0 $X=124980 $Y=99520
X2872 3 digital_ldo_top_VIA1 $T=125230 105200 0 0 $X=124980 $Y=104960
X2873 3 digital_ldo_top_VIA1 $T=125230 110640 0 0 $X=124980 $Y=110400
X2874 3 digital_ldo_top_VIA1 $T=125230 116080 0 0 $X=124980 $Y=115840
X2875 3 digital_ldo_top_VIA1 $T=125230 121520 0 0 $X=124980 $Y=121280
X2876 3 digital_ldo_top_VIA1 $T=125230 126960 0 0 $X=124980 $Y=126720
X2877 2 digital_ldo_top_VIA1 $T=126610 15440 0 0 $X=126360 $Y=15200
X2878 2 digital_ldo_top_VIA1 $T=126610 91600 0 0 $X=126360 $Y=91360
X2879 2 digital_ldo_top_VIA1 $T=126610 97040 0 0 $X=126360 $Y=96800
X2880 2 digital_ldo_top_VIA1 $T=126610 102480 0 0 $X=126360 $Y=102240
X2881 2 digital_ldo_top_VIA1 $T=126610 107920 0 0 $X=126360 $Y=107680
X2882 2 digital_ldo_top_VIA1 $T=126610 113360 0 0 $X=126360 $Y=113120
X2883 2 digital_ldo_top_VIA1 $T=126610 118800 0 0 $X=126360 $Y=118560
X2884 2 digital_ldo_top_VIA1 $T=126610 124240 0 0 $X=126360 $Y=124000
X2885 2 digital_ldo_top_VIA1 $T=126610 129680 0 0 $X=126360 $Y=129440
X2886 3 digital_ldo_top_VIA1 $T=128910 12720 0 0 $X=128660 $Y=12480
X2887 3 digital_ldo_top_VIA1 $T=128910 18160 0 0 $X=128660 $Y=17920
X2888 3 digital_ldo_top_VIA1 $T=128910 37720 0 0 $X=128660 $Y=37480
X2889 3 digital_ldo_top_VIA1 $T=128910 43160 0 0 $X=128660 $Y=42920
X2890 3 digital_ldo_top_VIA1 $T=128910 48600 0 0 $X=128660 $Y=48360
X2891 3 digital_ldo_top_VIA1 $T=128910 54040 0 0 $X=128660 $Y=53800
X2892 3 digital_ldo_top_VIA1 $T=128910 59480 0 0 $X=128660 $Y=59240
X2893 3 digital_ldo_top_VIA1 $T=128910 64920 0 0 $X=128660 $Y=64680
X2894 3 digital_ldo_top_VIA1 $T=128910 70360 0 0 $X=128660 $Y=70120
X2895 3 digital_ldo_top_VIA1 $T=128910 75800 0 0 $X=128660 $Y=75560
X2896 3 digital_ldo_top_VIA1 $T=128910 81240 0 0 $X=128660 $Y=81000
X2897 3 digital_ldo_top_VIA1 $T=128910 94320 0 0 $X=128660 $Y=94080
X2898 3 digital_ldo_top_VIA1 $T=128910 99760 0 0 $X=128660 $Y=99520
X2899 3 digital_ldo_top_VIA1 $T=128910 105200 0 0 $X=128660 $Y=104960
X2900 3 digital_ldo_top_VIA1 $T=128910 110640 0 0 $X=128660 $Y=110400
X2901 3 digital_ldo_top_VIA1 $T=128910 116080 0 0 $X=128660 $Y=115840
X2902 3 digital_ldo_top_VIA1 $T=128910 121520 0 0 $X=128660 $Y=121280
X2903 3 digital_ldo_top_VIA1 $T=128910 126960 0 0 $X=128660 $Y=126720
X2904 2 digital_ldo_top_VIA1 $T=130290 15440 0 0 $X=130040 $Y=15200
X2905 2 digital_ldo_top_VIA1 $T=130290 91600 0 0 $X=130040 $Y=91360
X2906 2 digital_ldo_top_VIA1 $T=130290 97040 0 0 $X=130040 $Y=96800
X2907 2 digital_ldo_top_VIA1 $T=130290 102480 0 0 $X=130040 $Y=102240
X2908 2 digital_ldo_top_VIA1 $T=130290 107920 0 0 $X=130040 $Y=107680
X2909 2 digital_ldo_top_VIA1 $T=130290 113360 0 0 $X=130040 $Y=113120
X2910 2 digital_ldo_top_VIA1 $T=130290 118800 0 0 $X=130040 $Y=118560
X2911 2 digital_ldo_top_VIA1 $T=130290 124240 0 0 $X=130040 $Y=124000
X2912 2 digital_ldo_top_VIA1 $T=130290 129680 0 0 $X=130040 $Y=129440
X2913 3 digital_ldo_top_VIA1 $T=132590 12720 0 0 $X=132340 $Y=12480
X2914 3 digital_ldo_top_VIA1 $T=132590 18160 0 0 $X=132340 $Y=17920
X2915 3 digital_ldo_top_VIA1 $T=132590 94320 0 0 $X=132340 $Y=94080
X2916 3 digital_ldo_top_VIA1 $T=132590 99760 0 0 $X=132340 $Y=99520
X2917 3 digital_ldo_top_VIA1 $T=132590 105200 0 0 $X=132340 $Y=104960
X2918 3 digital_ldo_top_VIA1 $T=132590 110640 0 0 $X=132340 $Y=110400
X2919 3 digital_ldo_top_VIA1 $T=132590 116080 0 0 $X=132340 $Y=115840
X2920 3 digital_ldo_top_VIA1 $T=132590 121520 0 0 $X=132340 $Y=121280
X2921 3 digital_ldo_top_VIA1 $T=132590 126960 0 0 $X=132340 $Y=126720
X2922 2 digital_ldo_top_VIA1 $T=133970 15440 0 0 $X=133720 $Y=15200
X2923 2 digital_ldo_top_VIA1 $T=133970 35000 0 0 $X=133720 $Y=34760
X2924 2 digital_ldo_top_VIA1 $T=133970 40440 0 0 $X=133720 $Y=40200
X2925 2 digital_ldo_top_VIA1 $T=133970 45880 0 0 $X=133720 $Y=45640
X2926 2 digital_ldo_top_VIA1 $T=133970 51320 0 0 $X=133720 $Y=51080
X2927 2 digital_ldo_top_VIA1 $T=133970 56760 0 0 $X=133720 $Y=56520
X2928 2 digital_ldo_top_VIA1 $T=133970 62200 0 0 $X=133720 $Y=61960
X2929 2 digital_ldo_top_VIA1 $T=133970 67640 0 0 $X=133720 $Y=67400
X2930 2 digital_ldo_top_VIA1 $T=133970 73080 0 0 $X=133720 $Y=72840
X2931 2 digital_ldo_top_VIA1 $T=133970 78520 0 0 $X=133720 $Y=78280
X2932 2 digital_ldo_top_VIA1 $T=133970 83960 0 0 $X=133720 $Y=83720
X2933 2 digital_ldo_top_VIA1 $T=133970 91600 0 0 $X=133720 $Y=91360
X2934 2 digital_ldo_top_VIA1 $T=133970 97040 0 0 $X=133720 $Y=96800
X2935 2 digital_ldo_top_VIA1 $T=133970 102480 0 0 $X=133720 $Y=102240
X2936 2 digital_ldo_top_VIA1 $T=133970 107920 0 0 $X=133720 $Y=107680
X2937 2 digital_ldo_top_VIA1 $T=133970 113360 0 0 $X=133720 $Y=113120
X2938 2 digital_ldo_top_VIA1 $T=133970 118800 0 0 $X=133720 $Y=118560
X2939 2 digital_ldo_top_VIA1 $T=133970 124240 0 0 $X=133720 $Y=124000
X2940 2 digital_ldo_top_VIA1 $T=133970 129680 0 0 $X=133720 $Y=129440
X2941 3 digital_ldo_top_VIA1 $T=136270 12720 0 0 $X=136020 $Y=12480
X2942 3 digital_ldo_top_VIA1 $T=136270 18160 0 0 $X=136020 $Y=17920
X2943 3 digital_ldo_top_VIA1 $T=136270 94320 0 0 $X=136020 $Y=94080
X2944 3 digital_ldo_top_VIA1 $T=136270 99760 0 0 $X=136020 $Y=99520
X2945 3 digital_ldo_top_VIA1 $T=136270 105200 0 0 $X=136020 $Y=104960
X2946 3 digital_ldo_top_VIA1 $T=136270 110640 0 0 $X=136020 $Y=110400
X2947 3 digital_ldo_top_VIA1 $T=136270 116080 0 0 $X=136020 $Y=115840
X2948 3 digital_ldo_top_VIA1 $T=136270 121520 0 0 $X=136020 $Y=121280
X2949 3 digital_ldo_top_VIA1 $T=136270 126960 0 0 $X=136020 $Y=126720
X2950 2 digital_ldo_top_VIA1 $T=137650 15440 0 0 $X=137400 $Y=15200
X2951 2 digital_ldo_top_VIA1 $T=137650 91600 0 0 $X=137400 $Y=91360
X2952 2 digital_ldo_top_VIA1 $T=137650 97040 0 0 $X=137400 $Y=96800
X2953 2 digital_ldo_top_VIA1 $T=137650 102480 0 0 $X=137400 $Y=102240
X2954 2 digital_ldo_top_VIA1 $T=137650 107920 0 0 $X=137400 $Y=107680
X2955 2 digital_ldo_top_VIA1 $T=137650 113360 0 0 $X=137400 $Y=113120
X2956 2 digital_ldo_top_VIA1 $T=137650 118800 0 0 $X=137400 $Y=118560
X2957 2 digital_ldo_top_VIA1 $T=137650 124240 0 0 $X=137400 $Y=124000
X2958 2 digital_ldo_top_VIA1 $T=137650 129680 0 0 $X=137400 $Y=129440
X2959 3 digital_ldo_top_VIA1 $T=139950 12720 0 0 $X=139700 $Y=12480
X2960 3 digital_ldo_top_VIA1 $T=139950 18160 0 0 $X=139700 $Y=17920
X2961 3 digital_ldo_top_VIA1 $T=139950 48600 0 0 $X=139700 $Y=48360
X2962 3 digital_ldo_top_VIA1 $T=139950 54040 0 0 $X=139700 $Y=53800
X2963 3 digital_ldo_top_VIA1 $T=139950 59480 0 0 $X=139700 $Y=59240
X2964 3 digital_ldo_top_VIA1 $T=139950 64920 0 0 $X=139700 $Y=64680
X2965 3 digital_ldo_top_VIA1 $T=139950 70360 0 0 $X=139700 $Y=70120
X2966 3 digital_ldo_top_VIA1 $T=139950 75800 0 0 $X=139700 $Y=75560
X2967 3 digital_ldo_top_VIA1 $T=139950 81240 0 0 $X=139700 $Y=81000
X2968 3 digital_ldo_top_VIA1 $T=139950 94320 0 0 $X=139700 $Y=94080
X2969 3 digital_ldo_top_VIA1 $T=139950 99760 0 0 $X=139700 $Y=99520
X2970 3 digital_ldo_top_VIA1 $T=139950 105200 0 0 $X=139700 $Y=104960
X2971 3 digital_ldo_top_VIA1 $T=139950 110640 0 0 $X=139700 $Y=110400
X2972 3 digital_ldo_top_VIA1 $T=139950 116080 0 0 $X=139700 $Y=115840
X2973 3 digital_ldo_top_VIA1 $T=139950 121520 0 0 $X=139700 $Y=121280
X2974 3 digital_ldo_top_VIA1 $T=139950 126960 0 0 $X=139700 $Y=126720
X2975 2 digital_ldo_top_VIA1 $T=141330 15440 0 0 $X=141080 $Y=15200
X2976 2 digital_ldo_top_VIA1 $T=141330 91600 0 0 $X=141080 $Y=91360
X2977 2 digital_ldo_top_VIA1 $T=141330 97040 0 0 $X=141080 $Y=96800
X2978 2 digital_ldo_top_VIA1 $T=141330 102480 0 0 $X=141080 $Y=102240
X2979 2 digital_ldo_top_VIA1 $T=141330 107920 0 0 $X=141080 $Y=107680
X2980 2 digital_ldo_top_VIA1 $T=141330 113360 0 0 $X=141080 $Y=113120
X2981 2 digital_ldo_top_VIA1 $T=141330 118800 0 0 $X=141080 $Y=118560
X2982 2 digital_ldo_top_VIA1 $T=141330 124240 0 0 $X=141080 $Y=124000
X2983 2 digital_ldo_top_VIA1 $T=141330 129680 0 0 $X=141080 $Y=129440
X2984 3 digital_ldo_top_VIA1 $T=143630 12720 0 0 $X=143380 $Y=12480
X2985 3 digital_ldo_top_VIA1 $T=143630 18160 0 0 $X=143380 $Y=17920
X2986 3 digital_ldo_top_VIA1 $T=143630 94320 0 0 $X=143380 $Y=94080
X2987 3 digital_ldo_top_VIA1 $T=143630 99760 0 0 $X=143380 $Y=99520
X2988 3 digital_ldo_top_VIA1 $T=143630 105200 0 0 $X=143380 $Y=104960
X2989 3 digital_ldo_top_VIA1 $T=143630 110640 0 0 $X=143380 $Y=110400
X2990 3 digital_ldo_top_VIA1 $T=143630 116080 0 0 $X=143380 $Y=115840
X2991 3 digital_ldo_top_VIA1 $T=143630 121520 0 0 $X=143380 $Y=121280
X2992 3 digital_ldo_top_VIA1 $T=143630 126960 0 0 $X=143380 $Y=126720
X2993 2 digital_ldo_top_VIA1 $T=145010 15440 0 0 $X=144760 $Y=15200
X2994 2 digital_ldo_top_VIA1 $T=145010 35000 0 0 $X=144760 $Y=34760
X2995 2 digital_ldo_top_VIA1 $T=145010 40440 0 0 $X=144760 $Y=40200
X2996 2 digital_ldo_top_VIA1 $T=145010 45880 0 0 $X=144760 $Y=45640
X2997 2 digital_ldo_top_VIA1 $T=145010 56760 0 0 $X=144760 $Y=56520
X2998 2 digital_ldo_top_VIA1 $T=145010 62200 0 0 $X=144760 $Y=61960
X2999 2 digital_ldo_top_VIA1 $T=145010 67640 0 0 $X=144760 $Y=67400
X3000 2 digital_ldo_top_VIA1 $T=145010 73080 0 0 $X=144760 $Y=72840
X3001 2 digital_ldo_top_VIA1 $T=145010 78520 0 0 $X=144760 $Y=78280
X3002 2 digital_ldo_top_VIA1 $T=145010 83960 0 0 $X=144760 $Y=83720
X3003 2 digital_ldo_top_VIA1 $T=145010 91600 0 0 $X=144760 $Y=91360
X3004 2 digital_ldo_top_VIA1 $T=145010 97040 0 0 $X=144760 $Y=96800
X3005 2 digital_ldo_top_VIA1 $T=145010 102480 0 0 $X=144760 $Y=102240
X3006 2 digital_ldo_top_VIA1 $T=145010 107920 0 0 $X=144760 $Y=107680
X3007 2 digital_ldo_top_VIA1 $T=145010 113360 0 0 $X=144760 $Y=113120
X3008 2 digital_ldo_top_VIA1 $T=145010 118800 0 0 $X=144760 $Y=118560
X3009 2 digital_ldo_top_VIA1 $T=145010 124240 0 0 $X=144760 $Y=124000
X3010 2 digital_ldo_top_VIA1 $T=145010 129680 0 0 $X=144760 $Y=129440
X3011 3 digital_ldo_top_VIA1 $T=147310 12720 0 0 $X=147060 $Y=12480
X3012 3 digital_ldo_top_VIA1 $T=147310 18160 0 0 $X=147060 $Y=17920
X3013 3 digital_ldo_top_VIA1 $T=147310 94320 0 0 $X=147060 $Y=94080
X3014 3 digital_ldo_top_VIA1 $T=147310 99760 0 0 $X=147060 $Y=99520
X3015 3 digital_ldo_top_VIA1 $T=147310 105200 0 0 $X=147060 $Y=104960
X3016 3 digital_ldo_top_VIA1 $T=147310 110640 0 0 $X=147060 $Y=110400
X3017 3 digital_ldo_top_VIA1 $T=147310 116080 0 0 $X=147060 $Y=115840
X3018 3 digital_ldo_top_VIA1 $T=147310 121520 0 0 $X=147060 $Y=121280
X3019 3 digital_ldo_top_VIA1 $T=147310 126960 0 0 $X=147060 $Y=126720
X3020 2 digital_ldo_top_VIA1 $T=148690 15440 0 0 $X=148440 $Y=15200
X3021 2 digital_ldo_top_VIA1 $T=148690 91600 0 0 $X=148440 $Y=91360
X3022 2 digital_ldo_top_VIA1 $T=148690 97040 0 0 $X=148440 $Y=96800
X3023 2 digital_ldo_top_VIA1 $T=148690 102480 0 0 $X=148440 $Y=102240
X3024 2 digital_ldo_top_VIA1 $T=148690 107920 0 0 $X=148440 $Y=107680
X3025 2 digital_ldo_top_VIA1 $T=148690 113360 0 0 $X=148440 $Y=113120
X3026 2 digital_ldo_top_VIA1 $T=148690 118800 0 0 $X=148440 $Y=118560
X3027 2 digital_ldo_top_VIA1 $T=148690 124240 0 0 $X=148440 $Y=124000
X3028 2 digital_ldo_top_VIA1 $T=148690 129680 0 0 $X=148440 $Y=129440
X3029 3 digital_ldo_top_VIA1 $T=150990 12720 0 0 $X=150740 $Y=12480
X3030 3 digital_ldo_top_VIA1 $T=150990 18160 0 0 $X=150740 $Y=17920
X3031 3 digital_ldo_top_VIA1 $T=150990 59480 0 0 $X=150740 $Y=59240
X3032 3 digital_ldo_top_VIA1 $T=150990 64920 0 0 $X=150740 $Y=64680
X3033 3 digital_ldo_top_VIA1 $T=150990 70360 0 0 $X=150740 $Y=70120
X3034 3 digital_ldo_top_VIA1 $T=150990 75800 0 0 $X=150740 $Y=75560
X3035 3 digital_ldo_top_VIA1 $T=150990 81240 0 0 $X=150740 $Y=81000
X3036 3 digital_ldo_top_VIA1 $T=150990 94320 0 0 $X=150740 $Y=94080
X3037 3 digital_ldo_top_VIA1 $T=150990 99760 0 0 $X=150740 $Y=99520
X3038 3 digital_ldo_top_VIA1 $T=150990 105200 0 0 $X=150740 $Y=104960
X3039 3 digital_ldo_top_VIA1 $T=150990 110640 0 0 $X=150740 $Y=110400
X3040 3 digital_ldo_top_VIA1 $T=150990 116080 0 0 $X=150740 $Y=115840
X3041 3 digital_ldo_top_VIA1 $T=150990 121520 0 0 $X=150740 $Y=121280
X3042 3 digital_ldo_top_VIA1 $T=150990 126960 0 0 $X=150740 $Y=126720
X3043 2 digital_ldo_top_VIA1 $T=152370 15440 0 0 $X=152120 $Y=15200
X3044 2 digital_ldo_top_VIA1 $T=152370 91600 0 0 $X=152120 $Y=91360
X3045 2 digital_ldo_top_VIA1 $T=152370 97040 0 0 $X=152120 $Y=96800
X3046 2 digital_ldo_top_VIA1 $T=152370 102480 0 0 $X=152120 $Y=102240
X3047 2 digital_ldo_top_VIA1 $T=152370 107920 0 0 $X=152120 $Y=107680
X3048 2 digital_ldo_top_VIA1 $T=152370 113360 0 0 $X=152120 $Y=113120
X3049 2 digital_ldo_top_VIA1 $T=152370 118800 0 0 $X=152120 $Y=118560
X3050 2 digital_ldo_top_VIA1 $T=152370 124240 0 0 $X=152120 $Y=124000
X3051 2 digital_ldo_top_VIA1 $T=152370 129680 0 0 $X=152120 $Y=129440
X3052 3 digital_ldo_top_VIA1 $T=154670 12720 0 0 $X=154420 $Y=12480
X3053 3 digital_ldo_top_VIA1 $T=154670 18160 0 0 $X=154420 $Y=17920
X3054 3 digital_ldo_top_VIA1 $T=154670 94320 0 0 $X=154420 $Y=94080
X3055 3 digital_ldo_top_VIA1 $T=154670 99760 0 0 $X=154420 $Y=99520
X3056 3 digital_ldo_top_VIA1 $T=154670 105200 0 0 $X=154420 $Y=104960
X3057 3 digital_ldo_top_VIA1 $T=154670 110640 0 0 $X=154420 $Y=110400
X3058 3 digital_ldo_top_VIA1 $T=154670 116080 0 0 $X=154420 $Y=115840
X3059 3 digital_ldo_top_VIA1 $T=154670 121520 0 0 $X=154420 $Y=121280
X3060 3 digital_ldo_top_VIA1 $T=154670 126960 0 0 $X=154420 $Y=126720
X3061 2 digital_ldo_top_VIA1 $T=156050 15440 0 0 $X=155800 $Y=15200
X3062 2 digital_ldo_top_VIA1 $T=156050 35000 0 0 $X=155800 $Y=34760
X3063 2 digital_ldo_top_VIA1 $T=156050 40440 0 0 $X=155800 $Y=40200
X3064 2 digital_ldo_top_VIA1 $T=156050 45880 0 0 $X=155800 $Y=45640
X3065 2 digital_ldo_top_VIA1 $T=156050 51320 0 0 $X=155800 $Y=51080
X3066 2 digital_ldo_top_VIA1 $T=156050 56760 0 0 $X=155800 $Y=56520
X3067 2 digital_ldo_top_VIA1 $T=156050 62200 0 0 $X=155800 $Y=61960
X3068 2 digital_ldo_top_VIA1 $T=156050 67640 0 0 $X=155800 $Y=67400
X3069 2 digital_ldo_top_VIA1 $T=156050 73080 0 0 $X=155800 $Y=72840
X3070 2 digital_ldo_top_VIA1 $T=156050 78520 0 0 $X=155800 $Y=78280
X3071 2 digital_ldo_top_VIA1 $T=156050 83960 0 0 $X=155800 $Y=83720
X3072 2 digital_ldo_top_VIA1 $T=156050 91600 0 0 $X=155800 $Y=91360
X3073 2 digital_ldo_top_VIA1 $T=156050 97040 0 0 $X=155800 $Y=96800
X3074 2 digital_ldo_top_VIA1 $T=156050 102480 0 0 $X=155800 $Y=102240
X3075 2 digital_ldo_top_VIA1 $T=156050 107920 0 0 $X=155800 $Y=107680
X3076 2 digital_ldo_top_VIA1 $T=156050 113360 0 0 $X=155800 $Y=113120
X3077 2 digital_ldo_top_VIA1 $T=156050 118800 0 0 $X=155800 $Y=118560
X3078 2 digital_ldo_top_VIA1 $T=156050 124240 0 0 $X=155800 $Y=124000
X3079 2 digital_ldo_top_VIA1 $T=156050 129680 0 0 $X=155800 $Y=129440
X3080 3 digital_ldo_top_VIA1 $T=158350 12720 0 0 $X=158100 $Y=12480
X3081 3 digital_ldo_top_VIA1 $T=158350 18160 0 0 $X=158100 $Y=17920
X3082 3 digital_ldo_top_VIA1 $T=158350 94320 0 0 $X=158100 $Y=94080
X3083 3 digital_ldo_top_VIA1 $T=158350 99760 0 0 $X=158100 $Y=99520
X3084 3 digital_ldo_top_VIA1 $T=158350 105200 0 0 $X=158100 $Y=104960
X3085 3 digital_ldo_top_VIA1 $T=158350 110640 0 0 $X=158100 $Y=110400
X3086 3 digital_ldo_top_VIA1 $T=158350 116080 0 0 $X=158100 $Y=115840
X3087 3 digital_ldo_top_VIA1 $T=158350 121520 0 0 $X=158100 $Y=121280
X3088 3 digital_ldo_top_VIA1 $T=158350 126960 0 0 $X=158100 $Y=126720
X3089 2 digital_ldo_top_VIA1 $T=159730 15440 0 0 $X=159480 $Y=15200
X3090 2 digital_ldo_top_VIA1 $T=159730 91600 0 0 $X=159480 $Y=91360
X3091 2 digital_ldo_top_VIA1 $T=159730 97040 0 0 $X=159480 $Y=96800
X3092 2 digital_ldo_top_VIA1 $T=159730 102480 0 0 $X=159480 $Y=102240
X3093 2 digital_ldo_top_VIA1 $T=159730 107920 0 0 $X=159480 $Y=107680
X3094 2 digital_ldo_top_VIA1 $T=159730 113360 0 0 $X=159480 $Y=113120
X3095 2 digital_ldo_top_VIA1 $T=159730 118800 0 0 $X=159480 $Y=118560
X3096 2 digital_ldo_top_VIA1 $T=159730 124240 0 0 $X=159480 $Y=124000
X3097 2 digital_ldo_top_VIA1 $T=159730 129680 0 0 $X=159480 $Y=129440
X3098 3 digital_ldo_top_VIA1 $T=162030 12720 0 0 $X=161780 $Y=12480
X3099 3 digital_ldo_top_VIA1 $T=162030 18160 0 0 $X=161780 $Y=17920
X3100 3 digital_ldo_top_VIA1 $T=162030 59480 0 0 $X=161780 $Y=59240
X3101 3 digital_ldo_top_VIA1 $T=162030 64920 0 0 $X=161780 $Y=64680
X3102 3 digital_ldo_top_VIA1 $T=162030 70360 0 0 $X=161780 $Y=70120
X3103 3 digital_ldo_top_VIA1 $T=162030 75800 0 0 $X=161780 $Y=75560
X3104 3 digital_ldo_top_VIA1 $T=162030 81240 0 0 $X=161780 $Y=81000
X3105 3 digital_ldo_top_VIA1 $T=162030 94320 0 0 $X=161780 $Y=94080
X3106 3 digital_ldo_top_VIA1 $T=162030 99760 0 0 $X=161780 $Y=99520
X3107 3 digital_ldo_top_VIA1 $T=162030 105200 0 0 $X=161780 $Y=104960
X3108 3 digital_ldo_top_VIA1 $T=162030 110640 0 0 $X=161780 $Y=110400
X3109 3 digital_ldo_top_VIA1 $T=162030 116080 0 0 $X=161780 $Y=115840
X3110 3 digital_ldo_top_VIA1 $T=162030 121520 0 0 $X=161780 $Y=121280
X3111 3 digital_ldo_top_VIA1 $T=162030 126960 0 0 $X=161780 $Y=126720
X3112 2 digital_ldo_top_VIA1 $T=163410 15440 0 0 $X=163160 $Y=15200
X3113 2 digital_ldo_top_VIA1 $T=163410 91600 0 0 $X=163160 $Y=91360
X3114 2 digital_ldo_top_VIA1 $T=163410 97040 0 0 $X=163160 $Y=96800
X3115 2 digital_ldo_top_VIA1 $T=163410 102480 0 0 $X=163160 $Y=102240
X3116 2 digital_ldo_top_VIA1 $T=163410 107920 0 0 $X=163160 $Y=107680
X3117 2 digital_ldo_top_VIA1 $T=163410 113360 0 0 $X=163160 $Y=113120
X3118 2 digital_ldo_top_VIA1 $T=163410 118800 0 0 $X=163160 $Y=118560
X3119 2 digital_ldo_top_VIA1 $T=163410 124240 0 0 $X=163160 $Y=124000
X3120 2 digital_ldo_top_VIA1 $T=163410 129680 0 0 $X=163160 $Y=129440
X3121 3 digital_ldo_top_VIA1 $T=165710 12720 0 0 $X=165460 $Y=12480
X3122 3 digital_ldo_top_VIA1 $T=165710 18160 0 0 $X=165460 $Y=17920
X3123 3 digital_ldo_top_VIA1 $T=165710 94320 0 0 $X=165460 $Y=94080
X3124 3 digital_ldo_top_VIA1 $T=165710 99760 0 0 $X=165460 $Y=99520
X3125 3 digital_ldo_top_VIA1 $T=165710 105200 0 0 $X=165460 $Y=104960
X3126 3 digital_ldo_top_VIA1 $T=165710 110640 0 0 $X=165460 $Y=110400
X3127 3 digital_ldo_top_VIA1 $T=165710 116080 0 0 $X=165460 $Y=115840
X3128 3 digital_ldo_top_VIA1 $T=165710 121520 0 0 $X=165460 $Y=121280
X3129 3 digital_ldo_top_VIA1 $T=165710 126960 0 0 $X=165460 $Y=126720
X3130 2 digital_ldo_top_VIA1 $T=167090 15440 0 0 $X=166840 $Y=15200
X3131 2 digital_ldo_top_VIA1 $T=167090 35000 0 0 $X=166840 $Y=34760
X3132 2 digital_ldo_top_VIA1 $T=167090 45880 0 0 $X=166840 $Y=45640
X3133 2 digital_ldo_top_VIA1 $T=167090 51320 0 0 $X=166840 $Y=51080
X3134 2 digital_ldo_top_VIA1 $T=167090 56760 0 0 $X=166840 $Y=56520
X3135 2 digital_ldo_top_VIA1 $T=167090 62200 0 0 $X=166840 $Y=61960
X3136 2 digital_ldo_top_VIA1 $T=167090 67640 0 0 $X=166840 $Y=67400
X3137 2 digital_ldo_top_VIA1 $T=167090 73080 0 0 $X=166840 $Y=72840
X3138 2 digital_ldo_top_VIA1 $T=167090 78520 0 0 $X=166840 $Y=78280
X3139 2 digital_ldo_top_VIA1 $T=167090 83960 0 0 $X=166840 $Y=83720
X3140 2 digital_ldo_top_VIA1 $T=167090 91600 0 0 $X=166840 $Y=91360
X3141 2 digital_ldo_top_VIA1 $T=167090 97040 0 0 $X=166840 $Y=96800
X3142 2 digital_ldo_top_VIA1 $T=167090 102480 0 0 $X=166840 $Y=102240
X3143 2 digital_ldo_top_VIA1 $T=167090 107920 0 0 $X=166840 $Y=107680
X3144 2 digital_ldo_top_VIA1 $T=167090 113360 0 0 $X=166840 $Y=113120
X3145 2 digital_ldo_top_VIA1 $T=167090 118800 0 0 $X=166840 $Y=118560
X3146 2 digital_ldo_top_VIA1 $T=167090 124240 0 0 $X=166840 $Y=124000
X3147 2 digital_ldo_top_VIA1 $T=167090 129680 0 0 $X=166840 $Y=129440
X3148 3 digital_ldo_top_VIA1 $T=169390 12720 0 0 $X=169140 $Y=12480
X3149 3 digital_ldo_top_VIA1 $T=169390 18160 0 0 $X=169140 $Y=17920
X3150 3 digital_ldo_top_VIA1 $T=169390 94320 0 0 $X=169140 $Y=94080
X3151 3 digital_ldo_top_VIA1 $T=169390 99760 0 0 $X=169140 $Y=99520
X3152 3 digital_ldo_top_VIA1 $T=169390 105200 0 0 $X=169140 $Y=104960
X3153 3 digital_ldo_top_VIA1 $T=169390 110640 0 0 $X=169140 $Y=110400
X3154 3 digital_ldo_top_VIA1 $T=169390 116080 0 0 $X=169140 $Y=115840
X3155 3 digital_ldo_top_VIA1 $T=169390 121520 0 0 $X=169140 $Y=121280
X3156 3 digital_ldo_top_VIA1 $T=169390 126960 0 0 $X=169140 $Y=126720
X3157 2 digital_ldo_top_VIA1 $T=170770 15440 0 0 $X=170520 $Y=15200
X3158 2 digital_ldo_top_VIA1 $T=170770 91600 0 0 $X=170520 $Y=91360
X3159 2 digital_ldo_top_VIA1 $T=170770 97040 0 0 $X=170520 $Y=96800
X3160 2 digital_ldo_top_VIA1 $T=170770 102480 0 0 $X=170520 $Y=102240
X3161 2 digital_ldo_top_VIA1 $T=170770 107920 0 0 $X=170520 $Y=107680
X3162 2 digital_ldo_top_VIA1 $T=170770 113360 0 0 $X=170520 $Y=113120
X3163 2 digital_ldo_top_VIA1 $T=170770 118800 0 0 $X=170520 $Y=118560
X3164 2 digital_ldo_top_VIA1 $T=170770 124240 0 0 $X=170520 $Y=124000
X3165 2 digital_ldo_top_VIA1 $T=170770 129680 0 0 $X=170520 $Y=129440
X3166 3 digital_ldo_top_VIA1 $T=173070 12720 0 0 $X=172820 $Y=12480
X3167 3 digital_ldo_top_VIA1 $T=173070 18160 0 0 $X=172820 $Y=17920
X3168 3 digital_ldo_top_VIA1 $T=173070 54040 0 0 $X=172820 $Y=53800
X3169 3 digital_ldo_top_VIA1 $T=173070 59480 0 0 $X=172820 $Y=59240
X3170 3 digital_ldo_top_VIA1 $T=173070 64920 0 0 $X=172820 $Y=64680
X3171 3 digital_ldo_top_VIA1 $T=173070 70360 0 0 $X=172820 $Y=70120
X3172 3 digital_ldo_top_VIA1 $T=173070 75800 0 0 $X=172820 $Y=75560
X3173 3 digital_ldo_top_VIA1 $T=173070 81240 0 0 $X=172820 $Y=81000
X3174 3 digital_ldo_top_VIA1 $T=173070 94320 0 0 $X=172820 $Y=94080
X3175 3 digital_ldo_top_VIA1 $T=173070 99760 0 0 $X=172820 $Y=99520
X3176 3 digital_ldo_top_VIA1 $T=173070 105200 0 0 $X=172820 $Y=104960
X3177 3 digital_ldo_top_VIA1 $T=173070 110640 0 0 $X=172820 $Y=110400
X3178 3 digital_ldo_top_VIA1 $T=173070 116080 0 0 $X=172820 $Y=115840
X3179 3 digital_ldo_top_VIA1 $T=173070 121520 0 0 $X=172820 $Y=121280
X3180 3 digital_ldo_top_VIA1 $T=173070 126960 0 0 $X=172820 $Y=126720
X3181 2 digital_ldo_top_VIA1 $T=174450 15440 0 0 $X=174200 $Y=15200
X3182 2 digital_ldo_top_VIA1 $T=174450 91600 0 0 $X=174200 $Y=91360
X3183 2 digital_ldo_top_VIA1 $T=174450 97040 0 0 $X=174200 $Y=96800
X3184 2 digital_ldo_top_VIA1 $T=174450 102480 0 0 $X=174200 $Y=102240
X3185 2 digital_ldo_top_VIA1 $T=174450 107920 0 0 $X=174200 $Y=107680
X3186 2 digital_ldo_top_VIA1 $T=174450 113360 0 0 $X=174200 $Y=113120
X3187 2 digital_ldo_top_VIA1 $T=174450 118800 0 0 $X=174200 $Y=118560
X3188 2 digital_ldo_top_VIA1 $T=174450 124240 0 0 $X=174200 $Y=124000
X3189 2 digital_ldo_top_VIA1 $T=174450 129680 0 0 $X=174200 $Y=129440
X3190 3 digital_ldo_top_VIA1 $T=176750 12720 0 0 $X=176500 $Y=12480
X3191 3 digital_ldo_top_VIA1 $T=176750 18160 0 0 $X=176500 $Y=17920
X3192 3 digital_ldo_top_VIA1 $T=176750 94320 0 0 $X=176500 $Y=94080
X3193 3 digital_ldo_top_VIA1 $T=176750 99760 0 0 $X=176500 $Y=99520
X3194 3 digital_ldo_top_VIA1 $T=176750 105200 0 0 $X=176500 $Y=104960
X3195 3 digital_ldo_top_VIA1 $T=176750 110640 0 0 $X=176500 $Y=110400
X3196 3 digital_ldo_top_VIA1 $T=176750 116080 0 0 $X=176500 $Y=115840
X3197 3 digital_ldo_top_VIA1 $T=176750 121520 0 0 $X=176500 $Y=121280
X3198 3 digital_ldo_top_VIA1 $T=176750 126960 0 0 $X=176500 $Y=126720
X3199 2 digital_ldo_top_VIA1 $T=178130 15440 0 0 $X=177880 $Y=15200
X3200 2 digital_ldo_top_VIA1 $T=178130 35000 0 0 $X=177880 $Y=34760
X3201 2 digital_ldo_top_VIA1 $T=178130 40440 0 0 $X=177880 $Y=40200
X3202 2 digital_ldo_top_VIA1 $T=178130 45880 0 0 $X=177880 $Y=45640
X3203 2 digital_ldo_top_VIA1 $T=178130 51320 0 0 $X=177880 $Y=51080
X3204 2 digital_ldo_top_VIA1 $T=178130 56760 0 0 $X=177880 $Y=56520
X3205 2 digital_ldo_top_VIA1 $T=178130 62200 0 0 $X=177880 $Y=61960
X3206 2 digital_ldo_top_VIA1 $T=178130 67640 0 0 $X=177880 $Y=67400
X3207 2 digital_ldo_top_VIA1 $T=178130 73080 0 0 $X=177880 $Y=72840
X3208 2 digital_ldo_top_VIA1 $T=178130 78520 0 0 $X=177880 $Y=78280
X3209 2 digital_ldo_top_VIA1 $T=178130 83960 0 0 $X=177880 $Y=83720
X3210 2 digital_ldo_top_VIA1 $T=178130 91600 0 0 $X=177880 $Y=91360
X3211 2 digital_ldo_top_VIA1 $T=178130 97040 0 0 $X=177880 $Y=96800
X3212 2 digital_ldo_top_VIA1 $T=178130 102480 0 0 $X=177880 $Y=102240
X3213 2 digital_ldo_top_VIA1 $T=178130 107920 0 0 $X=177880 $Y=107680
X3214 2 digital_ldo_top_VIA1 $T=178130 113360 0 0 $X=177880 $Y=113120
X3215 2 digital_ldo_top_VIA1 $T=178130 118800 0 0 $X=177880 $Y=118560
X3216 2 digital_ldo_top_VIA1 $T=178130 124240 0 0 $X=177880 $Y=124000
X3217 2 digital_ldo_top_VIA1 $T=178130 129680 0 0 $X=177880 $Y=129440
X3218 3 digital_ldo_top_VIA1 $T=180430 12720 0 0 $X=180180 $Y=12480
X3219 3 digital_ldo_top_VIA1 $T=180430 18160 0 0 $X=180180 $Y=17920
X3220 3 digital_ldo_top_VIA1 $T=180430 94320 0 0 $X=180180 $Y=94080
X3221 3 digital_ldo_top_VIA1 $T=180430 99760 0 0 $X=180180 $Y=99520
X3222 3 digital_ldo_top_VIA1 $T=180430 105200 0 0 $X=180180 $Y=104960
X3223 3 digital_ldo_top_VIA1 $T=180430 110640 0 0 $X=180180 $Y=110400
X3224 3 digital_ldo_top_VIA1 $T=180430 116080 0 0 $X=180180 $Y=115840
X3225 3 digital_ldo_top_VIA1 $T=180430 121520 0 0 $X=180180 $Y=121280
X3226 3 digital_ldo_top_VIA1 $T=180430 126960 0 0 $X=180180 $Y=126720
X3227 2 digital_ldo_top_VIA1 $T=181810 15440 0 0 $X=181560 $Y=15200
X3228 2 digital_ldo_top_VIA1 $T=181810 91600 0 0 $X=181560 $Y=91360
X3229 2 digital_ldo_top_VIA1 $T=181810 97040 0 0 $X=181560 $Y=96800
X3230 2 digital_ldo_top_VIA1 $T=181810 102480 0 0 $X=181560 $Y=102240
X3231 2 digital_ldo_top_VIA1 $T=181810 107920 0 0 $X=181560 $Y=107680
X3232 2 digital_ldo_top_VIA1 $T=181810 113360 0 0 $X=181560 $Y=113120
X3233 2 digital_ldo_top_VIA1 $T=181810 118800 0 0 $X=181560 $Y=118560
X3234 2 digital_ldo_top_VIA1 $T=181810 124240 0 0 $X=181560 $Y=124000
X3235 2 digital_ldo_top_VIA1 $T=181810 129680 0 0 $X=181560 $Y=129440
X3236 3 digital_ldo_top_VIA1 $T=184110 12720 0 0 $X=183860 $Y=12480
X3237 3 digital_ldo_top_VIA1 $T=184110 18160 0 0 $X=183860 $Y=17920
X3238 3 digital_ldo_top_VIA1 $T=184110 59480 0 0 $X=183860 $Y=59240
X3239 3 digital_ldo_top_VIA1 $T=184110 64920 0 0 $X=183860 $Y=64680
X3240 3 digital_ldo_top_VIA1 $T=184110 70360 0 0 $X=183860 $Y=70120
X3241 3 digital_ldo_top_VIA1 $T=184110 75800 0 0 $X=183860 $Y=75560
X3242 3 digital_ldo_top_VIA1 $T=184110 81240 0 0 $X=183860 $Y=81000
X3243 3 digital_ldo_top_VIA1 $T=184110 94320 0 0 $X=183860 $Y=94080
X3244 3 digital_ldo_top_VIA1 $T=184110 99760 0 0 $X=183860 $Y=99520
X3245 3 digital_ldo_top_VIA1 $T=184110 105200 0 0 $X=183860 $Y=104960
X3246 3 digital_ldo_top_VIA1 $T=184110 110640 0 0 $X=183860 $Y=110400
X3247 3 digital_ldo_top_VIA1 $T=184110 116080 0 0 $X=183860 $Y=115840
X3248 3 digital_ldo_top_VIA1 $T=184110 121520 0 0 $X=183860 $Y=121280
X3249 3 digital_ldo_top_VIA1 $T=184110 126960 0 0 $X=183860 $Y=126720
X3250 2 digital_ldo_top_VIA1 $T=185490 15440 0 0 $X=185240 $Y=15200
X3251 2 digital_ldo_top_VIA1 $T=185490 91600 0 0 $X=185240 $Y=91360
X3252 2 digital_ldo_top_VIA1 $T=185490 97040 0 0 $X=185240 $Y=96800
X3253 2 digital_ldo_top_VIA1 $T=185490 102480 0 0 $X=185240 $Y=102240
X3254 2 digital_ldo_top_VIA1 $T=185490 107920 0 0 $X=185240 $Y=107680
X3255 2 digital_ldo_top_VIA1 $T=185490 113360 0 0 $X=185240 $Y=113120
X3256 2 digital_ldo_top_VIA1 $T=185490 118800 0 0 $X=185240 $Y=118560
X3257 2 digital_ldo_top_VIA1 $T=185490 124240 0 0 $X=185240 $Y=124000
X3258 2 digital_ldo_top_VIA1 $T=185490 129680 0 0 $X=185240 $Y=129440
X3259 3 digital_ldo_top_VIA1 $T=187790 12720 0 0 $X=187540 $Y=12480
X3260 3 digital_ldo_top_VIA1 $T=187790 18160 0 0 $X=187540 $Y=17920
X3261 3 digital_ldo_top_VIA1 $T=187790 94320 0 0 $X=187540 $Y=94080
X3262 3 digital_ldo_top_VIA1 $T=187790 99760 0 0 $X=187540 $Y=99520
X3263 3 digital_ldo_top_VIA1 $T=187790 105200 0 0 $X=187540 $Y=104960
X3264 3 digital_ldo_top_VIA1 $T=187790 110640 0 0 $X=187540 $Y=110400
X3265 3 digital_ldo_top_VIA1 $T=187790 116080 0 0 $X=187540 $Y=115840
X3266 3 digital_ldo_top_VIA1 $T=187790 121520 0 0 $X=187540 $Y=121280
X3267 3 digital_ldo_top_VIA1 $T=187790 126960 0 0 $X=187540 $Y=126720
X3268 2 digital_ldo_top_VIA1 $T=189170 15440 0 0 $X=188920 $Y=15200
X3269 2 digital_ldo_top_VIA1 $T=189170 35000 0 0 $X=188920 $Y=34760
X3270 2 digital_ldo_top_VIA1 $T=189170 40440 0 0 $X=188920 $Y=40200
X3271 2 digital_ldo_top_VIA1 $T=189170 51320 0 0 $X=188920 $Y=51080
X3272 2 digital_ldo_top_VIA1 $T=189170 56760 0 0 $X=188920 $Y=56520
X3273 2 digital_ldo_top_VIA1 $T=189170 62200 0 0 $X=188920 $Y=61960
X3274 2 digital_ldo_top_VIA1 $T=189170 67640 0 0 $X=188920 $Y=67400
X3275 2 digital_ldo_top_VIA1 $T=189170 73080 0 0 $X=188920 $Y=72840
X3276 2 digital_ldo_top_VIA1 $T=189170 78520 0 0 $X=188920 $Y=78280
X3277 2 digital_ldo_top_VIA1 $T=189170 83960 0 0 $X=188920 $Y=83720
X3278 2 digital_ldo_top_VIA1 $T=189170 91600 0 0 $X=188920 $Y=91360
X3279 2 digital_ldo_top_VIA1 $T=189170 97040 0 0 $X=188920 $Y=96800
X3280 2 digital_ldo_top_VIA1 $T=189170 102480 0 0 $X=188920 $Y=102240
X3281 2 digital_ldo_top_VIA1 $T=189170 107920 0 0 $X=188920 $Y=107680
X3282 2 digital_ldo_top_VIA1 $T=189170 113360 0 0 $X=188920 $Y=113120
X3283 2 digital_ldo_top_VIA1 $T=189170 118800 0 0 $X=188920 $Y=118560
X3284 2 digital_ldo_top_VIA1 $T=189170 124240 0 0 $X=188920 $Y=124000
X3285 2 digital_ldo_top_VIA1 $T=189170 129680 0 0 $X=188920 $Y=129440
X3286 3 digital_ldo_top_VIA1 $T=191470 12720 0 0 $X=191220 $Y=12480
X3287 3 digital_ldo_top_VIA1 $T=191470 18160 0 0 $X=191220 $Y=17920
X3288 3 digital_ldo_top_VIA1 $T=191470 94320 0 0 $X=191220 $Y=94080
X3289 3 digital_ldo_top_VIA1 $T=191470 99760 0 0 $X=191220 $Y=99520
X3290 3 digital_ldo_top_VIA1 $T=191470 105200 0 0 $X=191220 $Y=104960
X3291 3 digital_ldo_top_VIA1 $T=191470 110640 0 0 $X=191220 $Y=110400
X3292 3 digital_ldo_top_VIA1 $T=191470 116080 0 0 $X=191220 $Y=115840
X3293 3 digital_ldo_top_VIA1 $T=191470 121520 0 0 $X=191220 $Y=121280
X3294 3 digital_ldo_top_VIA1 $T=191470 126960 0 0 $X=191220 $Y=126720
X3295 2 digital_ldo_top_VIA1 $T=192850 15440 0 0 $X=192600 $Y=15200
X3296 2 digital_ldo_top_VIA1 $T=192850 91600 0 0 $X=192600 $Y=91360
X3297 2 digital_ldo_top_VIA1 $T=192850 97040 0 0 $X=192600 $Y=96800
X3298 2 digital_ldo_top_VIA1 $T=192850 102480 0 0 $X=192600 $Y=102240
X3299 2 digital_ldo_top_VIA1 $T=192850 107920 0 0 $X=192600 $Y=107680
X3300 2 digital_ldo_top_VIA1 $T=192850 113360 0 0 $X=192600 $Y=113120
X3301 2 digital_ldo_top_VIA1 $T=192850 118800 0 0 $X=192600 $Y=118560
X3302 2 digital_ldo_top_VIA1 $T=192850 124240 0 0 $X=192600 $Y=124000
X3303 2 digital_ldo_top_VIA1 $T=192850 129680 0 0 $X=192600 $Y=129440
X3304 3 digital_ldo_top_VIA1 $T=195150 12720 0 0 $X=194900 $Y=12480
X3305 3 digital_ldo_top_VIA1 $T=195150 18160 0 0 $X=194900 $Y=17920
X3306 3 digital_ldo_top_VIA1 $T=195150 59480 0 0 $X=194900 $Y=59240
X3307 3 digital_ldo_top_VIA1 $T=195150 64920 0 0 $X=194900 $Y=64680
X3308 3 digital_ldo_top_VIA1 $T=195150 70360 0 0 $X=194900 $Y=70120
X3309 3 digital_ldo_top_VIA1 $T=195150 75800 0 0 $X=194900 $Y=75560
X3310 3 digital_ldo_top_VIA1 $T=195150 81240 0 0 $X=194900 $Y=81000
X3311 3 digital_ldo_top_VIA1 $T=195150 94320 0 0 $X=194900 $Y=94080
X3312 3 digital_ldo_top_VIA1 $T=195150 99760 0 0 $X=194900 $Y=99520
X3313 3 digital_ldo_top_VIA1 $T=195150 105200 0 0 $X=194900 $Y=104960
X3314 3 digital_ldo_top_VIA1 $T=195150 110640 0 0 $X=194900 $Y=110400
X3315 3 digital_ldo_top_VIA1 $T=195150 116080 0 0 $X=194900 $Y=115840
X3316 3 digital_ldo_top_VIA1 $T=195150 121520 0 0 $X=194900 $Y=121280
X3317 3 digital_ldo_top_VIA1 $T=195150 126960 0 0 $X=194900 $Y=126720
X3318 2 digital_ldo_top_VIA1 $T=196530 15440 0 0 $X=196280 $Y=15200
X3319 2 digital_ldo_top_VIA1 $T=196530 91600 0 0 $X=196280 $Y=91360
X3320 2 digital_ldo_top_VIA1 $T=196530 97040 0 0 $X=196280 $Y=96800
X3321 2 digital_ldo_top_VIA1 $T=196530 102480 0 0 $X=196280 $Y=102240
X3322 2 digital_ldo_top_VIA1 $T=196530 107920 0 0 $X=196280 $Y=107680
X3323 2 digital_ldo_top_VIA1 $T=196530 113360 0 0 $X=196280 $Y=113120
X3324 2 digital_ldo_top_VIA1 $T=196530 118800 0 0 $X=196280 $Y=118560
X3325 2 digital_ldo_top_VIA1 $T=196530 124240 0 0 $X=196280 $Y=124000
X3326 2 digital_ldo_top_VIA1 $T=196530 129680 0 0 $X=196280 $Y=129440
X3327 3 digital_ldo_top_VIA1 $T=198830 12720 0 0 $X=198580 $Y=12480
X3328 3 digital_ldo_top_VIA1 $T=198830 18160 0 0 $X=198580 $Y=17920
X3329 3 digital_ldo_top_VIA1 $T=198830 94320 0 0 $X=198580 $Y=94080
X3330 3 digital_ldo_top_VIA1 $T=198830 99760 0 0 $X=198580 $Y=99520
X3331 3 digital_ldo_top_VIA1 $T=198830 105200 0 0 $X=198580 $Y=104960
X3332 3 digital_ldo_top_VIA1 $T=198830 110640 0 0 $X=198580 $Y=110400
X3333 3 digital_ldo_top_VIA1 $T=198830 116080 0 0 $X=198580 $Y=115840
X3334 3 digital_ldo_top_VIA1 $T=198830 121520 0 0 $X=198580 $Y=121280
X3335 3 digital_ldo_top_VIA1 $T=198830 126960 0 0 $X=198580 $Y=126720
X3336 2 digital_ldo_top_VIA1 $T=200210 15440 0 0 $X=199960 $Y=15200
X3337 2 digital_ldo_top_VIA1 $T=200210 51320 0 0 $X=199960 $Y=51080
X3338 2 digital_ldo_top_VIA1 $T=200210 56760 0 0 $X=199960 $Y=56520
X3339 2 digital_ldo_top_VIA1 $T=200210 62200 0 0 $X=199960 $Y=61960
X3340 2 digital_ldo_top_VIA1 $T=200210 67640 0 0 $X=199960 $Y=67400
X3341 2 digital_ldo_top_VIA1 $T=200210 73080 0 0 $X=199960 $Y=72840
X3342 2 digital_ldo_top_VIA1 $T=200210 78520 0 0 $X=199960 $Y=78280
X3343 2 digital_ldo_top_VIA1 $T=200210 83960 0 0 $X=199960 $Y=83720
X3344 2 digital_ldo_top_VIA1 $T=200210 91600 0 0 $X=199960 $Y=91360
X3345 2 digital_ldo_top_VIA1 $T=200210 97040 0 0 $X=199960 $Y=96800
X3346 2 digital_ldo_top_VIA1 $T=200210 102480 0 0 $X=199960 $Y=102240
X3347 2 digital_ldo_top_VIA1 $T=200210 107920 0 0 $X=199960 $Y=107680
X3348 2 digital_ldo_top_VIA1 $T=200210 113360 0 0 $X=199960 $Y=113120
X3349 2 digital_ldo_top_VIA1 $T=200210 118800 0 0 $X=199960 $Y=118560
X3350 2 digital_ldo_top_VIA1 $T=200210 124240 0 0 $X=199960 $Y=124000
X3351 2 digital_ldo_top_VIA1 $T=200210 129680 0 0 $X=199960 $Y=129440
X3352 3 digital_ldo_top_VIA1 $T=202510 12720 0 0 $X=202260 $Y=12480
X3353 3 digital_ldo_top_VIA1 $T=202510 18160 0 0 $X=202260 $Y=17920
X3354 3 digital_ldo_top_VIA1 $T=202510 94320 0 0 $X=202260 $Y=94080
X3355 3 digital_ldo_top_VIA1 $T=202510 99760 0 0 $X=202260 $Y=99520
X3356 3 digital_ldo_top_VIA1 $T=202510 105200 0 0 $X=202260 $Y=104960
X3357 3 digital_ldo_top_VIA1 $T=202510 110640 0 0 $X=202260 $Y=110400
X3358 3 digital_ldo_top_VIA1 $T=202510 116080 0 0 $X=202260 $Y=115840
X3359 3 digital_ldo_top_VIA1 $T=202510 121520 0 0 $X=202260 $Y=121280
X3360 3 digital_ldo_top_VIA1 $T=202510 126960 0 0 $X=202260 $Y=126720
X3361 2 digital_ldo_top_VIA1 $T=203890 15440 0 0 $X=203640 $Y=15200
X3362 2 digital_ldo_top_VIA1 $T=203890 91600 0 0 $X=203640 $Y=91360
X3363 2 digital_ldo_top_VIA1 $T=203890 97040 0 0 $X=203640 $Y=96800
X3364 2 digital_ldo_top_VIA1 $T=203890 102480 0 0 $X=203640 $Y=102240
X3365 2 digital_ldo_top_VIA1 $T=203890 107920 0 0 $X=203640 $Y=107680
X3366 2 digital_ldo_top_VIA1 $T=203890 113360 0 0 $X=203640 $Y=113120
X3367 2 digital_ldo_top_VIA1 $T=203890 118800 0 0 $X=203640 $Y=118560
X3368 2 digital_ldo_top_VIA1 $T=203890 124240 0 0 $X=203640 $Y=124000
X3369 2 digital_ldo_top_VIA1 $T=203890 129680 0 0 $X=203640 $Y=129440
X3370 3 digital_ldo_top_VIA1 $T=206190 12720 0 0 $X=205940 $Y=12480
X3371 3 digital_ldo_top_VIA1 $T=206190 18160 0 0 $X=205940 $Y=17920
X3372 3 digital_ldo_top_VIA1 $T=206190 59480 0 0 $X=205940 $Y=59240
X3373 3 digital_ldo_top_VIA1 $T=206190 64920 0 0 $X=205940 $Y=64680
X3374 3 digital_ldo_top_VIA1 $T=206190 70360 0 0 $X=205940 $Y=70120
X3375 3 digital_ldo_top_VIA1 $T=206190 75800 0 0 $X=205940 $Y=75560
X3376 3 digital_ldo_top_VIA1 $T=206190 81240 0 0 $X=205940 $Y=81000
X3377 3 digital_ldo_top_VIA1 $T=206190 94320 0 0 $X=205940 $Y=94080
X3378 3 digital_ldo_top_VIA1 $T=206190 99760 0 0 $X=205940 $Y=99520
X3379 3 digital_ldo_top_VIA1 $T=206190 105200 0 0 $X=205940 $Y=104960
X3380 3 digital_ldo_top_VIA1 $T=206190 110640 0 0 $X=205940 $Y=110400
X3381 3 digital_ldo_top_VIA1 $T=206190 116080 0 0 $X=205940 $Y=115840
X3382 3 digital_ldo_top_VIA1 $T=206190 121520 0 0 $X=205940 $Y=121280
X3383 3 digital_ldo_top_VIA1 $T=206190 126960 0 0 $X=205940 $Y=126720
X3384 2 digital_ldo_top_VIA1 $T=207570 15440 0 0 $X=207320 $Y=15200
X3385 2 digital_ldo_top_VIA1 $T=207570 91600 0 0 $X=207320 $Y=91360
X3386 2 digital_ldo_top_VIA1 $T=207570 97040 0 0 $X=207320 $Y=96800
X3387 2 digital_ldo_top_VIA1 $T=207570 102480 0 0 $X=207320 $Y=102240
X3388 2 digital_ldo_top_VIA1 $T=207570 107920 0 0 $X=207320 $Y=107680
X3389 2 digital_ldo_top_VIA1 $T=207570 113360 0 0 $X=207320 $Y=113120
X3390 2 digital_ldo_top_VIA1 $T=207570 118800 0 0 $X=207320 $Y=118560
X3391 2 digital_ldo_top_VIA1 $T=207570 124240 0 0 $X=207320 $Y=124000
X3392 2 digital_ldo_top_VIA1 $T=207570 129680 0 0 $X=207320 $Y=129440
X3393 3 digital_ldo_top_VIA1 $T=209870 12720 0 0 $X=209620 $Y=12480
X3394 3 digital_ldo_top_VIA1 $T=209870 18160 0 0 $X=209620 $Y=17920
X3395 3 digital_ldo_top_VIA1 $T=209870 94320 0 0 $X=209620 $Y=94080
X3396 3 digital_ldo_top_VIA1 $T=209870 99760 0 0 $X=209620 $Y=99520
X3397 3 digital_ldo_top_VIA1 $T=209870 105200 0 0 $X=209620 $Y=104960
X3398 3 digital_ldo_top_VIA1 $T=209870 110640 0 0 $X=209620 $Y=110400
X3399 3 digital_ldo_top_VIA1 $T=209870 116080 0 0 $X=209620 $Y=115840
X3400 3 digital_ldo_top_VIA1 $T=209870 121520 0 0 $X=209620 $Y=121280
X3401 3 digital_ldo_top_VIA1 $T=209870 126960 0 0 $X=209620 $Y=126720
X3402 2 digital_ldo_top_VIA1 $T=211250 15440 0 0 $X=211000 $Y=15200
X3403 2 digital_ldo_top_VIA1 $T=211250 35000 0 0 $X=211000 $Y=34760
X3404 2 digital_ldo_top_VIA1 $T=211250 40440 0 0 $X=211000 $Y=40200
X3405 2 digital_ldo_top_VIA1 $T=211250 45880 0 0 $X=211000 $Y=45640
X3406 2 digital_ldo_top_VIA1 $T=211250 51320 0 0 $X=211000 $Y=51080
X3407 2 digital_ldo_top_VIA1 $T=211250 56760 0 0 $X=211000 $Y=56520
X3408 2 digital_ldo_top_VIA1 $T=211250 62200 0 0 $X=211000 $Y=61960
X3409 2 digital_ldo_top_VIA1 $T=211250 67640 0 0 $X=211000 $Y=67400
X3410 2 digital_ldo_top_VIA1 $T=211250 73080 0 0 $X=211000 $Y=72840
X3411 2 digital_ldo_top_VIA1 $T=211250 78520 0 0 $X=211000 $Y=78280
X3412 2 digital_ldo_top_VIA1 $T=211250 83960 0 0 $X=211000 $Y=83720
X3413 2 digital_ldo_top_VIA1 $T=211250 91600 0 0 $X=211000 $Y=91360
X3414 2 digital_ldo_top_VIA1 $T=211250 97040 0 0 $X=211000 $Y=96800
X3415 2 digital_ldo_top_VIA1 $T=211250 102480 0 0 $X=211000 $Y=102240
X3416 2 digital_ldo_top_VIA1 $T=211250 107920 0 0 $X=211000 $Y=107680
X3417 2 digital_ldo_top_VIA1 $T=211250 113360 0 0 $X=211000 $Y=113120
X3418 2 digital_ldo_top_VIA1 $T=211250 118800 0 0 $X=211000 $Y=118560
X3419 2 digital_ldo_top_VIA1 $T=211250 124240 0 0 $X=211000 $Y=124000
X3420 2 digital_ldo_top_VIA1 $T=211250 129680 0 0 $X=211000 $Y=129440
X3421 3 digital_ldo_top_VIA1 $T=213550 12720 0 0 $X=213300 $Y=12480
X3422 3 digital_ldo_top_VIA1 $T=213550 18160 0 0 $X=213300 $Y=17920
X3423 3 digital_ldo_top_VIA1 $T=213550 94320 0 0 $X=213300 $Y=94080
X3424 3 digital_ldo_top_VIA1 $T=213550 99760 0 0 $X=213300 $Y=99520
X3425 3 digital_ldo_top_VIA1 $T=213550 105200 0 0 $X=213300 $Y=104960
X3426 3 digital_ldo_top_VIA1 $T=213550 110640 0 0 $X=213300 $Y=110400
X3427 3 digital_ldo_top_VIA1 $T=213550 116080 0 0 $X=213300 $Y=115840
X3428 3 digital_ldo_top_VIA1 $T=213550 121520 0 0 $X=213300 $Y=121280
X3429 3 digital_ldo_top_VIA1 $T=213550 126960 0 0 $X=213300 $Y=126720
X3430 2 digital_ldo_top_VIA1 $T=214930 15440 0 0 $X=214680 $Y=15200
X3431 2 digital_ldo_top_VIA1 $T=214930 91600 0 0 $X=214680 $Y=91360
X3432 2 digital_ldo_top_VIA1 $T=214930 97040 0 0 $X=214680 $Y=96800
X3433 2 digital_ldo_top_VIA1 $T=214930 102480 0 0 $X=214680 $Y=102240
X3434 2 digital_ldo_top_VIA1 $T=214930 107920 0 0 $X=214680 $Y=107680
X3435 2 digital_ldo_top_VIA1 $T=214930 113360 0 0 $X=214680 $Y=113120
X3436 2 digital_ldo_top_VIA1 $T=214930 118800 0 0 $X=214680 $Y=118560
X3437 2 digital_ldo_top_VIA1 $T=214930 124240 0 0 $X=214680 $Y=124000
X3438 2 digital_ldo_top_VIA1 $T=214930 129680 0 0 $X=214680 $Y=129440
X3439 3 digital_ldo_top_VIA1 $T=217230 12720 0 0 $X=216980 $Y=12480
X3440 3 digital_ldo_top_VIA1 $T=217230 18160 0 0 $X=216980 $Y=17920
X3441 3 digital_ldo_top_VIA1 $T=217230 37720 0 0 $X=216980 $Y=37480
X3442 3 digital_ldo_top_VIA1 $T=217230 59480 0 0 $X=216980 $Y=59240
X3443 3 digital_ldo_top_VIA1 $T=217230 64920 0 0 $X=216980 $Y=64680
X3444 3 digital_ldo_top_VIA1 $T=217230 70360 0 0 $X=216980 $Y=70120
X3445 3 digital_ldo_top_VIA1 $T=217230 75800 0 0 $X=216980 $Y=75560
X3446 3 digital_ldo_top_VIA1 $T=217230 81240 0 0 $X=216980 $Y=81000
X3447 3 digital_ldo_top_VIA1 $T=217230 94320 0 0 $X=216980 $Y=94080
X3448 3 digital_ldo_top_VIA1 $T=217230 99760 0 0 $X=216980 $Y=99520
X3449 3 digital_ldo_top_VIA1 $T=217230 105200 0 0 $X=216980 $Y=104960
X3450 3 digital_ldo_top_VIA1 $T=217230 110640 0 0 $X=216980 $Y=110400
X3451 3 digital_ldo_top_VIA1 $T=217230 116080 0 0 $X=216980 $Y=115840
X3452 3 digital_ldo_top_VIA1 $T=217230 121520 0 0 $X=216980 $Y=121280
X3453 3 digital_ldo_top_VIA1 $T=217230 126960 0 0 $X=216980 $Y=126720
X3454 2 digital_ldo_top_VIA1 $T=218610 15440 0 0 $X=218360 $Y=15200
X3455 2 digital_ldo_top_VIA1 $T=218610 91600 0 0 $X=218360 $Y=91360
X3456 2 digital_ldo_top_VIA1 $T=218610 97040 0 0 $X=218360 $Y=96800
X3457 2 digital_ldo_top_VIA1 $T=218610 102480 0 0 $X=218360 $Y=102240
X3458 2 digital_ldo_top_VIA1 $T=218610 107920 0 0 $X=218360 $Y=107680
X3459 2 digital_ldo_top_VIA1 $T=218610 113360 0 0 $X=218360 $Y=113120
X3460 2 digital_ldo_top_VIA1 $T=218610 118800 0 0 $X=218360 $Y=118560
X3461 2 digital_ldo_top_VIA1 $T=218610 124240 0 0 $X=218360 $Y=124000
X3462 2 digital_ldo_top_VIA1 $T=218610 129680 0 0 $X=218360 $Y=129440
X3463 3 digital_ldo_top_VIA1 $T=220910 12720 0 0 $X=220660 $Y=12480
X3464 3 digital_ldo_top_VIA1 $T=220910 18160 0 0 $X=220660 $Y=17920
X3465 3 digital_ldo_top_VIA1 $T=220910 94320 0 0 $X=220660 $Y=94080
X3466 3 digital_ldo_top_VIA1 $T=220910 99760 0 0 $X=220660 $Y=99520
X3467 3 digital_ldo_top_VIA1 $T=220910 105200 0 0 $X=220660 $Y=104960
X3468 3 digital_ldo_top_VIA1 $T=220910 110640 0 0 $X=220660 $Y=110400
X3469 3 digital_ldo_top_VIA1 $T=220910 116080 0 0 $X=220660 $Y=115840
X3470 3 digital_ldo_top_VIA1 $T=220910 121520 0 0 $X=220660 $Y=121280
X3471 3 digital_ldo_top_VIA1 $T=220910 126960 0 0 $X=220660 $Y=126720
X3472 2 digital_ldo_top_VIA1 $T=222290 15440 0 0 $X=222040 $Y=15200
X3473 2 digital_ldo_top_VIA1 $T=222290 35000 0 0 $X=222040 $Y=34760
X3474 2 digital_ldo_top_VIA1 $T=222290 40440 0 0 $X=222040 $Y=40200
X3475 2 digital_ldo_top_VIA1 $T=222290 45880 0 0 $X=222040 $Y=45640
X3476 2 digital_ldo_top_VIA1 $T=222290 51320 0 0 $X=222040 $Y=51080
X3477 2 digital_ldo_top_VIA1 $T=222290 56760 0 0 $X=222040 $Y=56520
X3478 2 digital_ldo_top_VIA1 $T=222290 62200 0 0 $X=222040 $Y=61960
X3479 2 digital_ldo_top_VIA1 $T=222290 67640 0 0 $X=222040 $Y=67400
X3480 2 digital_ldo_top_VIA1 $T=222290 73080 0 0 $X=222040 $Y=72840
X3481 2 digital_ldo_top_VIA1 $T=222290 78520 0 0 $X=222040 $Y=78280
X3482 2 digital_ldo_top_VIA1 $T=222290 83960 0 0 $X=222040 $Y=83720
X3483 2 digital_ldo_top_VIA1 $T=222290 91600 0 0 $X=222040 $Y=91360
X3484 2 digital_ldo_top_VIA1 $T=222290 97040 0 0 $X=222040 $Y=96800
X3485 2 digital_ldo_top_VIA1 $T=222290 102480 0 0 $X=222040 $Y=102240
X3486 2 digital_ldo_top_VIA1 $T=222290 107920 0 0 $X=222040 $Y=107680
X3487 2 digital_ldo_top_VIA1 $T=222290 113360 0 0 $X=222040 $Y=113120
X3488 2 digital_ldo_top_VIA1 $T=222290 118800 0 0 $X=222040 $Y=118560
X3489 2 digital_ldo_top_VIA1 $T=222290 124240 0 0 $X=222040 $Y=124000
X3490 2 digital_ldo_top_VIA1 $T=222290 129680 0 0 $X=222040 $Y=129440
X3491 3 digital_ldo_top_VIA1 $T=224590 12720 0 0 $X=224340 $Y=12480
X3492 3 digital_ldo_top_VIA1 $T=224590 18160 0 0 $X=224340 $Y=17920
X3493 3 digital_ldo_top_VIA1 $T=224590 94320 0 0 $X=224340 $Y=94080
X3494 3 digital_ldo_top_VIA1 $T=224590 99760 0 0 $X=224340 $Y=99520
X3495 3 digital_ldo_top_VIA1 $T=224590 105200 0 0 $X=224340 $Y=104960
X3496 3 digital_ldo_top_VIA1 $T=224590 110640 0 0 $X=224340 $Y=110400
X3497 3 digital_ldo_top_VIA1 $T=224590 116080 0 0 $X=224340 $Y=115840
X3498 3 digital_ldo_top_VIA1 $T=224590 121520 0 0 $X=224340 $Y=121280
X3499 3 digital_ldo_top_VIA1 $T=224590 126960 0 0 $X=224340 $Y=126720
X3500 2 digital_ldo_top_VIA1 $T=225970 15440 0 0 $X=225720 $Y=15200
X3501 2 digital_ldo_top_VIA1 $T=225970 91600 0 0 $X=225720 $Y=91360
X3502 2 digital_ldo_top_VIA1 $T=225970 97040 0 0 $X=225720 $Y=96800
X3503 2 digital_ldo_top_VIA1 $T=225970 102480 0 0 $X=225720 $Y=102240
X3504 2 digital_ldo_top_VIA1 $T=225970 107920 0 0 $X=225720 $Y=107680
X3505 2 digital_ldo_top_VIA1 $T=225970 113360 0 0 $X=225720 $Y=113120
X3506 2 digital_ldo_top_VIA1 $T=225970 118800 0 0 $X=225720 $Y=118560
X3507 2 digital_ldo_top_VIA1 $T=225970 124240 0 0 $X=225720 $Y=124000
X3508 2 digital_ldo_top_VIA1 $T=225970 129680 0 0 $X=225720 $Y=129440
X3509 3 digital_ldo_top_VIA1 $T=228270 12720 0 0 $X=228020 $Y=12480
X3510 3 digital_ldo_top_VIA1 $T=228270 18160 0 0 $X=228020 $Y=17920
X3511 3 digital_ldo_top_VIA1 $T=228270 59480 0 0 $X=228020 $Y=59240
X3512 3 digital_ldo_top_VIA1 $T=228270 64920 0 0 $X=228020 $Y=64680
X3513 3 digital_ldo_top_VIA1 $T=228270 70360 0 0 $X=228020 $Y=70120
X3514 3 digital_ldo_top_VIA1 $T=228270 75800 0 0 $X=228020 $Y=75560
X3515 3 digital_ldo_top_VIA1 $T=228270 81240 0 0 $X=228020 $Y=81000
X3516 3 digital_ldo_top_VIA1 $T=228270 94320 0 0 $X=228020 $Y=94080
X3517 3 digital_ldo_top_VIA1 $T=228270 99760 0 0 $X=228020 $Y=99520
X3518 3 digital_ldo_top_VIA1 $T=228270 105200 0 0 $X=228020 $Y=104960
X3519 3 digital_ldo_top_VIA1 $T=228270 110640 0 0 $X=228020 $Y=110400
X3520 3 digital_ldo_top_VIA1 $T=228270 116080 0 0 $X=228020 $Y=115840
X3521 3 digital_ldo_top_VIA1 $T=228270 121520 0 0 $X=228020 $Y=121280
X3522 3 digital_ldo_top_VIA1 $T=228270 126960 0 0 $X=228020 $Y=126720
X3523 2 digital_ldo_top_VIA1 $T=229650 15440 0 0 $X=229400 $Y=15200
X3524 2 digital_ldo_top_VIA1 $T=229650 91600 0 0 $X=229400 $Y=91360
X3525 2 digital_ldo_top_VIA1 $T=229650 97040 0 0 $X=229400 $Y=96800
X3526 2 digital_ldo_top_VIA1 $T=229650 102480 0 0 $X=229400 $Y=102240
X3527 2 digital_ldo_top_VIA1 $T=229650 107920 0 0 $X=229400 $Y=107680
X3528 2 digital_ldo_top_VIA1 $T=229650 113360 0 0 $X=229400 $Y=113120
X3529 2 digital_ldo_top_VIA1 $T=229650 118800 0 0 $X=229400 $Y=118560
X3530 2 digital_ldo_top_VIA1 $T=229650 124240 0 0 $X=229400 $Y=124000
X3531 2 digital_ldo_top_VIA1 $T=229650 129680 0 0 $X=229400 $Y=129440
X3532 3 digital_ldo_top_VIA1 $T=231950 12720 0 0 $X=231700 $Y=12480
X3533 3 digital_ldo_top_VIA1 $T=231950 18160 0 0 $X=231700 $Y=17920
X3534 3 digital_ldo_top_VIA1 $T=231950 94320 0 0 $X=231700 $Y=94080
X3535 3 digital_ldo_top_VIA1 $T=231950 99760 0 0 $X=231700 $Y=99520
X3536 3 digital_ldo_top_VIA1 $T=231950 105200 0 0 $X=231700 $Y=104960
X3537 3 digital_ldo_top_VIA1 $T=231950 110640 0 0 $X=231700 $Y=110400
X3538 3 digital_ldo_top_VIA1 $T=231950 116080 0 0 $X=231700 $Y=115840
X3539 3 digital_ldo_top_VIA1 $T=231950 121520 0 0 $X=231700 $Y=121280
X3540 3 digital_ldo_top_VIA1 $T=231950 126960 0 0 $X=231700 $Y=126720
X3541 2 digital_ldo_top_VIA1 $T=233330 15440 0 0 $X=233080 $Y=15200
X3542 2 digital_ldo_top_VIA1 $T=233330 35000 0 0 $X=233080 $Y=34760
X3543 2 digital_ldo_top_VIA1 $T=233330 51320 0 0 $X=233080 $Y=51080
X3544 2 digital_ldo_top_VIA1 $T=233330 56760 0 0 $X=233080 $Y=56520
X3545 2 digital_ldo_top_VIA1 $T=233330 62200 0 0 $X=233080 $Y=61960
X3546 2 digital_ldo_top_VIA1 $T=233330 67640 0 0 $X=233080 $Y=67400
X3547 2 digital_ldo_top_VIA1 $T=233330 73080 0 0 $X=233080 $Y=72840
X3548 2 digital_ldo_top_VIA1 $T=233330 78520 0 0 $X=233080 $Y=78280
X3549 2 digital_ldo_top_VIA1 $T=233330 83960 0 0 $X=233080 $Y=83720
X3550 2 digital_ldo_top_VIA1 $T=233330 91600 0 0 $X=233080 $Y=91360
X3551 2 digital_ldo_top_VIA1 $T=233330 97040 0 0 $X=233080 $Y=96800
X3552 2 digital_ldo_top_VIA1 $T=233330 102480 0 0 $X=233080 $Y=102240
X3553 2 digital_ldo_top_VIA1 $T=233330 107920 0 0 $X=233080 $Y=107680
X3554 2 digital_ldo_top_VIA1 $T=233330 113360 0 0 $X=233080 $Y=113120
X3555 2 digital_ldo_top_VIA1 $T=233330 118800 0 0 $X=233080 $Y=118560
X3556 2 digital_ldo_top_VIA1 $T=233330 124240 0 0 $X=233080 $Y=124000
X3557 2 digital_ldo_top_VIA1 $T=233330 129680 0 0 $X=233080 $Y=129440
X3558 3 digital_ldo_top_VIA1 $T=235630 12720 0 0 $X=235380 $Y=12480
X3559 3 digital_ldo_top_VIA1 $T=235630 18160 0 0 $X=235380 $Y=17920
X3560 3 digital_ldo_top_VIA1 $T=235630 94320 0 0 $X=235380 $Y=94080
X3561 3 digital_ldo_top_VIA1 $T=235630 99760 0 0 $X=235380 $Y=99520
X3562 3 digital_ldo_top_VIA1 $T=235630 105200 0 0 $X=235380 $Y=104960
X3563 3 digital_ldo_top_VIA1 $T=235630 110640 0 0 $X=235380 $Y=110400
X3564 3 digital_ldo_top_VIA1 $T=235630 116080 0 0 $X=235380 $Y=115840
X3565 3 digital_ldo_top_VIA1 $T=235630 121520 0 0 $X=235380 $Y=121280
X3566 3 digital_ldo_top_VIA1 $T=235630 126960 0 0 $X=235380 $Y=126720
X3567 2 digital_ldo_top_VIA1 $T=237010 15440 0 0 $X=236760 $Y=15200
X3568 2 digital_ldo_top_VIA1 $T=237010 91600 0 0 $X=236760 $Y=91360
X3569 2 digital_ldo_top_VIA1 $T=237010 97040 0 0 $X=236760 $Y=96800
X3570 2 digital_ldo_top_VIA1 $T=237010 102480 0 0 $X=236760 $Y=102240
X3571 2 digital_ldo_top_VIA1 $T=237010 107920 0 0 $X=236760 $Y=107680
X3572 2 digital_ldo_top_VIA1 $T=237010 113360 0 0 $X=236760 $Y=113120
X3573 2 digital_ldo_top_VIA1 $T=237010 118800 0 0 $X=236760 $Y=118560
X3574 2 digital_ldo_top_VIA1 $T=237010 124240 0 0 $X=236760 $Y=124000
X3575 2 digital_ldo_top_VIA1 $T=237010 129680 0 0 $X=236760 $Y=129440
X3576 3 digital_ldo_top_VIA1 $T=239310 12720 0 0 $X=239060 $Y=12480
X3577 3 digital_ldo_top_VIA1 $T=239310 18160 0 0 $X=239060 $Y=17920
X3578 3 digital_ldo_top_VIA1 $T=239310 54040 0 0 $X=239060 $Y=53800
X3579 3 digital_ldo_top_VIA1 $T=239310 59480 0 0 $X=239060 $Y=59240
X3580 3 digital_ldo_top_VIA1 $T=239310 64920 0 0 $X=239060 $Y=64680
X3581 3 digital_ldo_top_VIA1 $T=239310 70360 0 0 $X=239060 $Y=70120
X3582 3 digital_ldo_top_VIA1 $T=239310 75800 0 0 $X=239060 $Y=75560
X3583 3 digital_ldo_top_VIA1 $T=239310 81240 0 0 $X=239060 $Y=81000
X3584 3 digital_ldo_top_VIA1 $T=239310 94320 0 0 $X=239060 $Y=94080
X3585 3 digital_ldo_top_VIA1 $T=239310 99760 0 0 $X=239060 $Y=99520
X3586 3 digital_ldo_top_VIA1 $T=239310 105200 0 0 $X=239060 $Y=104960
X3587 3 digital_ldo_top_VIA1 $T=239310 110640 0 0 $X=239060 $Y=110400
X3588 3 digital_ldo_top_VIA1 $T=239310 116080 0 0 $X=239060 $Y=115840
X3589 3 digital_ldo_top_VIA1 $T=239310 121520 0 0 $X=239060 $Y=121280
X3590 3 digital_ldo_top_VIA1 $T=239310 126960 0 0 $X=239060 $Y=126720
X3591 2 digital_ldo_top_VIA1 $T=240690 15440 0 0 $X=240440 $Y=15200
X3592 2 digital_ldo_top_VIA1 $T=240690 91600 0 0 $X=240440 $Y=91360
X3593 2 digital_ldo_top_VIA1 $T=240690 97040 0 0 $X=240440 $Y=96800
X3594 2 digital_ldo_top_VIA1 $T=240690 102480 0 0 $X=240440 $Y=102240
X3595 2 digital_ldo_top_VIA1 $T=240690 107920 0 0 $X=240440 $Y=107680
X3596 2 digital_ldo_top_VIA1 $T=240690 113360 0 0 $X=240440 $Y=113120
X3597 2 digital_ldo_top_VIA1 $T=240690 118800 0 0 $X=240440 $Y=118560
X3598 2 digital_ldo_top_VIA1 $T=240690 124240 0 0 $X=240440 $Y=124000
X3599 2 digital_ldo_top_VIA1 $T=240690 129680 0 0 $X=240440 $Y=129440
X3600 3 digital_ldo_top_VIA1 $T=242990 12720 0 0 $X=242740 $Y=12480
X3601 3 digital_ldo_top_VIA1 $T=242990 18160 0 0 $X=242740 $Y=17920
X3602 3 digital_ldo_top_VIA1 $T=242990 94320 0 0 $X=242740 $Y=94080
X3603 3 digital_ldo_top_VIA1 $T=242990 99760 0 0 $X=242740 $Y=99520
X3604 3 digital_ldo_top_VIA1 $T=242990 105200 0 0 $X=242740 $Y=104960
X3605 3 digital_ldo_top_VIA1 $T=242990 110640 0 0 $X=242740 $Y=110400
X3606 3 digital_ldo_top_VIA1 $T=242990 116080 0 0 $X=242740 $Y=115840
X3607 3 digital_ldo_top_VIA1 $T=242990 121520 0 0 $X=242740 $Y=121280
X3608 3 digital_ldo_top_VIA1 $T=242990 126960 0 0 $X=242740 $Y=126720
X3609 2 digital_ldo_top_VIA1 $T=244370 15440 0 0 $X=244120 $Y=15200
X3610 2 digital_ldo_top_VIA1 $T=244370 35000 0 0 $X=244120 $Y=34760
X3611 2 digital_ldo_top_VIA1 $T=244370 45880 0 0 $X=244120 $Y=45640
X3612 2 digital_ldo_top_VIA1 $T=244370 51320 0 0 $X=244120 $Y=51080
X3613 2 digital_ldo_top_VIA1 $T=244370 56760 0 0 $X=244120 $Y=56520
X3614 2 digital_ldo_top_VIA1 $T=244370 62200 0 0 $X=244120 $Y=61960
X3615 2 digital_ldo_top_VIA1 $T=244370 67640 0 0 $X=244120 $Y=67400
X3616 2 digital_ldo_top_VIA1 $T=244370 73080 0 0 $X=244120 $Y=72840
X3617 2 digital_ldo_top_VIA1 $T=244370 78520 0 0 $X=244120 $Y=78280
X3618 2 digital_ldo_top_VIA1 $T=244370 83960 0 0 $X=244120 $Y=83720
X3619 2 digital_ldo_top_VIA1 $T=244370 91600 0 0 $X=244120 $Y=91360
X3620 2 digital_ldo_top_VIA1 $T=244370 97040 0 0 $X=244120 $Y=96800
X3621 2 digital_ldo_top_VIA1 $T=244370 102480 0 0 $X=244120 $Y=102240
X3622 2 digital_ldo_top_VIA1 $T=244370 107920 0 0 $X=244120 $Y=107680
X3623 2 digital_ldo_top_VIA1 $T=244370 113360 0 0 $X=244120 $Y=113120
X3624 2 digital_ldo_top_VIA1 $T=244370 118800 0 0 $X=244120 $Y=118560
X3625 2 digital_ldo_top_VIA1 $T=244370 124240 0 0 $X=244120 $Y=124000
X3626 2 digital_ldo_top_VIA1 $T=244370 129680 0 0 $X=244120 $Y=129440
X3627 3 digital_ldo_top_VIA1 $T=246670 12720 0 0 $X=246420 $Y=12480
X3628 3 digital_ldo_top_VIA1 $T=246670 18160 0 0 $X=246420 $Y=17920
X3629 3 digital_ldo_top_VIA1 $T=246670 94320 0 0 $X=246420 $Y=94080
X3630 3 digital_ldo_top_VIA1 $T=246670 99760 0 0 $X=246420 $Y=99520
X3631 3 digital_ldo_top_VIA1 $T=246670 105200 0 0 $X=246420 $Y=104960
X3632 3 digital_ldo_top_VIA1 $T=246670 110640 0 0 $X=246420 $Y=110400
X3633 3 digital_ldo_top_VIA1 $T=246670 116080 0 0 $X=246420 $Y=115840
X3634 3 digital_ldo_top_VIA1 $T=246670 121520 0 0 $X=246420 $Y=121280
X3635 3 digital_ldo_top_VIA1 $T=246670 126960 0 0 $X=246420 $Y=126720
X3636 2 digital_ldo_top_VIA1 $T=248050 15440 0 0 $X=247800 $Y=15200
X3637 2 digital_ldo_top_VIA1 $T=248050 91600 0 0 $X=247800 $Y=91360
X3638 2 digital_ldo_top_VIA1 $T=248050 97040 0 0 $X=247800 $Y=96800
X3639 2 digital_ldo_top_VIA1 $T=248050 102480 0 0 $X=247800 $Y=102240
X3640 2 digital_ldo_top_VIA1 $T=248050 107920 0 0 $X=247800 $Y=107680
X3641 2 digital_ldo_top_VIA1 $T=248050 113360 0 0 $X=247800 $Y=113120
X3642 2 digital_ldo_top_VIA1 $T=248050 118800 0 0 $X=247800 $Y=118560
X3643 2 digital_ldo_top_VIA1 $T=248050 124240 0 0 $X=247800 $Y=124000
X3644 2 digital_ldo_top_VIA1 $T=248050 129680 0 0 $X=247800 $Y=129440
X3645 3 digital_ldo_top_VIA1 $T=250350 12720 0 0 $X=250100 $Y=12480
X3646 3 digital_ldo_top_VIA1 $T=250350 18160 0 0 $X=250100 $Y=17920
X3647 3 digital_ldo_top_VIA1 $T=250350 37720 0 0 $X=250100 $Y=37480
X3648 3 digital_ldo_top_VIA1 $T=250350 54040 0 0 $X=250100 $Y=53800
X3649 3 digital_ldo_top_VIA1 $T=250350 59480 0 0 $X=250100 $Y=59240
X3650 3 digital_ldo_top_VIA1 $T=250350 64920 0 0 $X=250100 $Y=64680
X3651 3 digital_ldo_top_VIA1 $T=250350 70360 0 0 $X=250100 $Y=70120
X3652 3 digital_ldo_top_VIA1 $T=250350 75800 0 0 $X=250100 $Y=75560
X3653 3 digital_ldo_top_VIA1 $T=250350 81240 0 0 $X=250100 $Y=81000
X3654 3 digital_ldo_top_VIA1 $T=250350 94320 0 0 $X=250100 $Y=94080
X3655 3 digital_ldo_top_VIA1 $T=250350 99760 0 0 $X=250100 $Y=99520
X3656 3 digital_ldo_top_VIA1 $T=250350 105200 0 0 $X=250100 $Y=104960
X3657 3 digital_ldo_top_VIA1 $T=250350 110640 0 0 $X=250100 $Y=110400
X3658 3 digital_ldo_top_VIA1 $T=250350 116080 0 0 $X=250100 $Y=115840
X3659 3 digital_ldo_top_VIA1 $T=250350 121520 0 0 $X=250100 $Y=121280
X3660 3 digital_ldo_top_VIA1 $T=250350 126960 0 0 $X=250100 $Y=126720
X3661 2 digital_ldo_top_VIA1 $T=251730 15440 0 0 $X=251480 $Y=15200
X3662 2 digital_ldo_top_VIA1 $T=251730 91600 0 0 $X=251480 $Y=91360
X3663 2 digital_ldo_top_VIA1 $T=251730 97040 0 0 $X=251480 $Y=96800
X3664 2 digital_ldo_top_VIA1 $T=251730 102480 0 0 $X=251480 $Y=102240
X3665 2 digital_ldo_top_VIA1 $T=251730 107920 0 0 $X=251480 $Y=107680
X3666 2 digital_ldo_top_VIA1 $T=251730 113360 0 0 $X=251480 $Y=113120
X3667 2 digital_ldo_top_VIA1 $T=251730 118800 0 0 $X=251480 $Y=118560
X3668 2 digital_ldo_top_VIA1 $T=251730 124240 0 0 $X=251480 $Y=124000
X3669 2 digital_ldo_top_VIA1 $T=251730 129680 0 0 $X=251480 $Y=129440
X3670 3 digital_ldo_top_VIA1 $T=254030 12720 0 0 $X=253780 $Y=12480
X3671 3 digital_ldo_top_VIA1 $T=254030 18160 0 0 $X=253780 $Y=17920
X3672 3 digital_ldo_top_VIA1 $T=254030 94320 0 0 $X=253780 $Y=94080
X3673 3 digital_ldo_top_VIA1 $T=254030 99760 0 0 $X=253780 $Y=99520
X3674 3 digital_ldo_top_VIA1 $T=254030 105200 0 0 $X=253780 $Y=104960
X3675 3 digital_ldo_top_VIA1 $T=254030 110640 0 0 $X=253780 $Y=110400
X3676 3 digital_ldo_top_VIA1 $T=254030 116080 0 0 $X=253780 $Y=115840
X3677 3 digital_ldo_top_VIA1 $T=254030 121520 0 0 $X=253780 $Y=121280
X3678 3 digital_ldo_top_VIA1 $T=254030 126960 0 0 $X=253780 $Y=126720
X3679 2 digital_ldo_top_VIA1 $T=255410 15440 0 0 $X=255160 $Y=15200
X3680 2 digital_ldo_top_VIA1 $T=255410 45880 0 0 $X=255160 $Y=45640
X3681 2 digital_ldo_top_VIA1 $T=255410 51320 0 0 $X=255160 $Y=51080
X3682 2 digital_ldo_top_VIA1 $T=255410 56760 0 0 $X=255160 $Y=56520
X3683 2 digital_ldo_top_VIA1 $T=255410 62200 0 0 $X=255160 $Y=61960
X3684 2 digital_ldo_top_VIA1 $T=255410 67640 0 0 $X=255160 $Y=67400
X3685 2 digital_ldo_top_VIA1 $T=255410 73080 0 0 $X=255160 $Y=72840
X3686 2 digital_ldo_top_VIA1 $T=255410 78520 0 0 $X=255160 $Y=78280
X3687 2 digital_ldo_top_VIA1 $T=255410 83960 0 0 $X=255160 $Y=83720
X3688 2 digital_ldo_top_VIA1 $T=255410 91600 0 0 $X=255160 $Y=91360
X3689 2 digital_ldo_top_VIA1 $T=255410 97040 0 0 $X=255160 $Y=96800
X3690 2 digital_ldo_top_VIA1 $T=255410 102480 0 0 $X=255160 $Y=102240
X3691 2 digital_ldo_top_VIA1 $T=255410 107920 0 0 $X=255160 $Y=107680
X3692 2 digital_ldo_top_VIA1 $T=255410 113360 0 0 $X=255160 $Y=113120
X3693 2 digital_ldo_top_VIA1 $T=255410 118800 0 0 $X=255160 $Y=118560
X3694 2 digital_ldo_top_VIA1 $T=255410 124240 0 0 $X=255160 $Y=124000
X3695 2 digital_ldo_top_VIA1 $T=255410 129680 0 0 $X=255160 $Y=129440
X3696 3 digital_ldo_top_VIA1 $T=257710 12720 0 0 $X=257460 $Y=12480
X3697 3 digital_ldo_top_VIA1 $T=257710 18160 0 0 $X=257460 $Y=17920
X3698 3 digital_ldo_top_VIA1 $T=257710 94320 0 0 $X=257460 $Y=94080
X3699 3 digital_ldo_top_VIA1 $T=257710 99760 0 0 $X=257460 $Y=99520
X3700 3 digital_ldo_top_VIA1 $T=257710 105200 0 0 $X=257460 $Y=104960
X3701 3 digital_ldo_top_VIA1 $T=257710 110640 0 0 $X=257460 $Y=110400
X3702 3 digital_ldo_top_VIA1 $T=257710 116080 0 0 $X=257460 $Y=115840
X3703 3 digital_ldo_top_VIA1 $T=257710 121520 0 0 $X=257460 $Y=121280
X3704 3 digital_ldo_top_VIA1 $T=257710 126960 0 0 $X=257460 $Y=126720
X3705 2 digital_ldo_top_VIA1 $T=259090 15440 0 0 $X=258840 $Y=15200
X3706 2 digital_ldo_top_VIA1 $T=259090 91600 0 0 $X=258840 $Y=91360
X3707 2 digital_ldo_top_VIA1 $T=259090 97040 0 0 $X=258840 $Y=96800
X3708 2 digital_ldo_top_VIA1 $T=259090 102480 0 0 $X=258840 $Y=102240
X3709 2 digital_ldo_top_VIA1 $T=259090 107920 0 0 $X=258840 $Y=107680
X3710 2 digital_ldo_top_VIA1 $T=259090 113360 0 0 $X=258840 $Y=113120
X3711 2 digital_ldo_top_VIA1 $T=259090 118800 0 0 $X=258840 $Y=118560
X3712 2 digital_ldo_top_VIA1 $T=259090 124240 0 0 $X=258840 $Y=124000
X3713 2 digital_ldo_top_VIA1 $T=259090 129680 0 0 $X=258840 $Y=129440
X3714 3 digital_ldo_top_VIA1 $T=261390 12720 0 0 $X=261140 $Y=12480
X3715 3 digital_ldo_top_VIA1 $T=261390 18160 0 0 $X=261140 $Y=17920
X3716 3 digital_ldo_top_VIA1 $T=261390 37720 0 0 $X=261140 $Y=37480
X3717 3 digital_ldo_top_VIA1 $T=261390 59480 0 0 $X=261140 $Y=59240
X3718 3 digital_ldo_top_VIA1 $T=261390 64920 0 0 $X=261140 $Y=64680
X3719 3 digital_ldo_top_VIA1 $T=261390 70360 0 0 $X=261140 $Y=70120
X3720 3 digital_ldo_top_VIA1 $T=261390 75800 0 0 $X=261140 $Y=75560
X3721 3 digital_ldo_top_VIA1 $T=261390 81240 0 0 $X=261140 $Y=81000
X3722 3 digital_ldo_top_VIA1 $T=261390 94320 0 0 $X=261140 $Y=94080
X3723 3 digital_ldo_top_VIA1 $T=261390 99760 0 0 $X=261140 $Y=99520
X3724 3 digital_ldo_top_VIA1 $T=261390 105200 0 0 $X=261140 $Y=104960
X3725 3 digital_ldo_top_VIA1 $T=261390 110640 0 0 $X=261140 $Y=110400
X3726 3 digital_ldo_top_VIA1 $T=261390 116080 0 0 $X=261140 $Y=115840
X3727 3 digital_ldo_top_VIA1 $T=261390 121520 0 0 $X=261140 $Y=121280
X3728 3 digital_ldo_top_VIA1 $T=261390 126960 0 0 $X=261140 $Y=126720
X3729 2 digital_ldo_top_VIA1 $T=262770 15440 0 0 $X=262520 $Y=15200
X3730 2 digital_ldo_top_VIA1 $T=262770 91600 0 0 $X=262520 $Y=91360
X3731 2 digital_ldo_top_VIA1 $T=262770 97040 0 0 $X=262520 $Y=96800
X3732 2 digital_ldo_top_VIA1 $T=262770 102480 0 0 $X=262520 $Y=102240
X3733 2 digital_ldo_top_VIA1 $T=262770 107920 0 0 $X=262520 $Y=107680
X3734 2 digital_ldo_top_VIA1 $T=262770 113360 0 0 $X=262520 $Y=113120
X3735 2 digital_ldo_top_VIA1 $T=262770 118800 0 0 $X=262520 $Y=118560
X3736 2 digital_ldo_top_VIA1 $T=262770 124240 0 0 $X=262520 $Y=124000
X3737 2 digital_ldo_top_VIA1 $T=262770 129680 0 0 $X=262520 $Y=129440
X3738 3 digital_ldo_top_VIA1 $T=265070 12720 0 0 $X=264820 $Y=12480
X3739 3 digital_ldo_top_VIA1 $T=265070 18160 0 0 $X=264820 $Y=17920
X3740 3 digital_ldo_top_VIA1 $T=265070 94320 0 0 $X=264820 $Y=94080
X3741 3 digital_ldo_top_VIA1 $T=265070 99760 0 0 $X=264820 $Y=99520
X3742 3 digital_ldo_top_VIA1 $T=265070 105200 0 0 $X=264820 $Y=104960
X3743 3 digital_ldo_top_VIA1 $T=265070 110640 0 0 $X=264820 $Y=110400
X3744 3 digital_ldo_top_VIA1 $T=265070 116080 0 0 $X=264820 $Y=115840
X3745 3 digital_ldo_top_VIA1 $T=265070 121520 0 0 $X=264820 $Y=121280
X3746 3 digital_ldo_top_VIA1 $T=265070 126960 0 0 $X=264820 $Y=126720
X3747 2 digital_ldo_top_VIA1 $T=266450 15440 0 0 $X=266200 $Y=15200
X3748 2 digital_ldo_top_VIA1 $T=266450 40440 0 0 $X=266200 $Y=40200
X3749 2 digital_ldo_top_VIA1 $T=266450 45880 0 0 $X=266200 $Y=45640
X3750 2 digital_ldo_top_VIA1 $T=266450 51320 0 0 $X=266200 $Y=51080
X3751 2 digital_ldo_top_VIA1 $T=266450 56760 0 0 $X=266200 $Y=56520
X3752 2 digital_ldo_top_VIA1 $T=266450 62200 0 0 $X=266200 $Y=61960
X3753 2 digital_ldo_top_VIA1 $T=266450 67640 0 0 $X=266200 $Y=67400
X3754 2 digital_ldo_top_VIA1 $T=266450 73080 0 0 $X=266200 $Y=72840
X3755 2 digital_ldo_top_VIA1 $T=266450 78520 0 0 $X=266200 $Y=78280
X3756 2 digital_ldo_top_VIA1 $T=266450 83960 0 0 $X=266200 $Y=83720
X3757 2 digital_ldo_top_VIA1 $T=266450 91600 0 0 $X=266200 $Y=91360
X3758 2 digital_ldo_top_VIA1 $T=266450 97040 0 0 $X=266200 $Y=96800
X3759 2 digital_ldo_top_VIA1 $T=266450 102480 0 0 $X=266200 $Y=102240
X3760 2 digital_ldo_top_VIA1 $T=266450 107920 0 0 $X=266200 $Y=107680
X3761 2 digital_ldo_top_VIA1 $T=266450 113360 0 0 $X=266200 $Y=113120
X3762 2 digital_ldo_top_VIA1 $T=266450 118800 0 0 $X=266200 $Y=118560
X3763 2 digital_ldo_top_VIA1 $T=266450 124240 0 0 $X=266200 $Y=124000
X3764 2 digital_ldo_top_VIA1 $T=266450 129680 0 0 $X=266200 $Y=129440
X3765 3 digital_ldo_top_VIA1 $T=268750 12720 0 0 $X=268500 $Y=12480
X3766 3 digital_ldo_top_VIA1 $T=268750 18160 0 0 $X=268500 $Y=17920
X3767 3 digital_ldo_top_VIA1 $T=268750 94320 0 0 $X=268500 $Y=94080
X3768 3 digital_ldo_top_VIA1 $T=268750 99760 0 0 $X=268500 $Y=99520
X3769 3 digital_ldo_top_VIA1 $T=268750 105200 0 0 $X=268500 $Y=104960
X3770 3 digital_ldo_top_VIA1 $T=268750 110640 0 0 $X=268500 $Y=110400
X3771 3 digital_ldo_top_VIA1 $T=268750 116080 0 0 $X=268500 $Y=115840
X3772 3 digital_ldo_top_VIA1 $T=268750 121520 0 0 $X=268500 $Y=121280
X3773 3 digital_ldo_top_VIA1 $T=268750 126960 0 0 $X=268500 $Y=126720
X3774 2 digital_ldo_top_VIA1 $T=270130 15440 0 0 $X=269880 $Y=15200
X3775 2 digital_ldo_top_VIA1 $T=270130 91600 0 0 $X=269880 $Y=91360
X3776 2 digital_ldo_top_VIA1 $T=270130 97040 0 0 $X=269880 $Y=96800
X3777 2 digital_ldo_top_VIA1 $T=270130 102480 0 0 $X=269880 $Y=102240
X3778 2 digital_ldo_top_VIA1 $T=270130 107920 0 0 $X=269880 $Y=107680
X3779 2 digital_ldo_top_VIA1 $T=270130 113360 0 0 $X=269880 $Y=113120
X3780 2 digital_ldo_top_VIA1 $T=270130 118800 0 0 $X=269880 $Y=118560
X3781 2 digital_ldo_top_VIA1 $T=270130 124240 0 0 $X=269880 $Y=124000
X3782 2 digital_ldo_top_VIA1 $T=270130 129680 0 0 $X=269880 $Y=129440
X3783 3 digital_ldo_top_VIA1 $T=272430 12720 0 0 $X=272180 $Y=12480
X3784 3 digital_ldo_top_VIA1 $T=272430 18160 0 0 $X=272180 $Y=17920
X3785 3 digital_ldo_top_VIA1 $T=272430 54040 0 0 $X=272180 $Y=53800
X3786 3 digital_ldo_top_VIA1 $T=272430 59480 0 0 $X=272180 $Y=59240
X3787 3 digital_ldo_top_VIA1 $T=272430 64920 0 0 $X=272180 $Y=64680
X3788 3 digital_ldo_top_VIA1 $T=272430 70360 0 0 $X=272180 $Y=70120
X3789 3 digital_ldo_top_VIA1 $T=272430 75800 0 0 $X=272180 $Y=75560
X3790 3 digital_ldo_top_VIA1 $T=272430 81240 0 0 $X=272180 $Y=81000
X3791 3 digital_ldo_top_VIA1 $T=272430 94320 0 0 $X=272180 $Y=94080
X3792 3 digital_ldo_top_VIA1 $T=272430 99760 0 0 $X=272180 $Y=99520
X3793 3 digital_ldo_top_VIA1 $T=272430 105200 0 0 $X=272180 $Y=104960
X3794 3 digital_ldo_top_VIA1 $T=272430 110640 0 0 $X=272180 $Y=110400
X3795 3 digital_ldo_top_VIA1 $T=272430 116080 0 0 $X=272180 $Y=115840
X3796 3 digital_ldo_top_VIA1 $T=272430 121520 0 0 $X=272180 $Y=121280
X3797 3 digital_ldo_top_VIA1 $T=272430 126960 0 0 $X=272180 $Y=126720
X3798 2 digital_ldo_top_VIA1 $T=273810 15440 0 0 $X=273560 $Y=15200
X3799 2 digital_ldo_top_VIA1 $T=273810 91600 0 0 $X=273560 $Y=91360
X3800 2 digital_ldo_top_VIA1 $T=273810 97040 0 0 $X=273560 $Y=96800
X3801 2 digital_ldo_top_VIA1 $T=273810 102480 0 0 $X=273560 $Y=102240
X3802 2 digital_ldo_top_VIA1 $T=273810 107920 0 0 $X=273560 $Y=107680
X3803 2 digital_ldo_top_VIA1 $T=273810 113360 0 0 $X=273560 $Y=113120
X3804 2 digital_ldo_top_VIA1 $T=273810 118800 0 0 $X=273560 $Y=118560
X3805 2 digital_ldo_top_VIA1 $T=273810 124240 0 0 $X=273560 $Y=124000
X3806 2 digital_ldo_top_VIA1 $T=273810 129680 0 0 $X=273560 $Y=129440
X3807 3 digital_ldo_top_VIA1 $T=276110 12720 0 0 $X=275860 $Y=12480
X3808 3 digital_ldo_top_VIA1 $T=276110 18160 0 0 $X=275860 $Y=17920
X3809 3 digital_ldo_top_VIA1 $T=276110 94320 0 0 $X=275860 $Y=94080
X3810 3 digital_ldo_top_VIA1 $T=276110 99760 0 0 $X=275860 $Y=99520
X3811 3 digital_ldo_top_VIA1 $T=276110 105200 0 0 $X=275860 $Y=104960
X3812 3 digital_ldo_top_VIA1 $T=276110 110640 0 0 $X=275860 $Y=110400
X3813 3 digital_ldo_top_VIA1 $T=276110 116080 0 0 $X=275860 $Y=115840
X3814 3 digital_ldo_top_VIA1 $T=276110 121520 0 0 $X=275860 $Y=121280
X3815 3 digital_ldo_top_VIA1 $T=276110 126960 0 0 $X=275860 $Y=126720
X3816 2 digital_ldo_top_VIA1 $T=277490 15440 0 0 $X=277240 $Y=15200
X3817 2 digital_ldo_top_VIA1 $T=277490 35000 0 0 $X=277240 $Y=34760
X3818 2 digital_ldo_top_VIA1 $T=277490 51320 0 0 $X=277240 $Y=51080
X3819 2 digital_ldo_top_VIA1 $T=277490 56760 0 0 $X=277240 $Y=56520
X3820 2 digital_ldo_top_VIA1 $T=277490 62200 0 0 $X=277240 $Y=61960
X3821 2 digital_ldo_top_VIA1 $T=277490 67640 0 0 $X=277240 $Y=67400
X3822 2 digital_ldo_top_VIA1 $T=277490 73080 0 0 $X=277240 $Y=72840
X3823 2 digital_ldo_top_VIA1 $T=277490 78520 0 0 $X=277240 $Y=78280
X3824 2 digital_ldo_top_VIA1 $T=277490 83960 0 0 $X=277240 $Y=83720
X3825 2 digital_ldo_top_VIA1 $T=277490 91600 0 0 $X=277240 $Y=91360
X3826 2 digital_ldo_top_VIA1 $T=277490 97040 0 0 $X=277240 $Y=96800
X3827 2 digital_ldo_top_VIA1 $T=277490 102480 0 0 $X=277240 $Y=102240
X3828 2 digital_ldo_top_VIA1 $T=277490 107920 0 0 $X=277240 $Y=107680
X3829 2 digital_ldo_top_VIA1 $T=277490 113360 0 0 $X=277240 $Y=113120
X3830 2 digital_ldo_top_VIA1 $T=277490 118800 0 0 $X=277240 $Y=118560
X3831 2 digital_ldo_top_VIA1 $T=277490 124240 0 0 $X=277240 $Y=124000
X3832 2 digital_ldo_top_VIA1 $T=277490 129680 0 0 $X=277240 $Y=129440
X3833 3 digital_ldo_top_VIA1 $T=279790 12720 0 0 $X=279540 $Y=12480
X3834 3 digital_ldo_top_VIA1 $T=279790 18160 0 0 $X=279540 $Y=17920
X3835 3 digital_ldo_top_VIA1 $T=279790 94320 0 0 $X=279540 $Y=94080
X3836 3 digital_ldo_top_VIA1 $T=279790 99760 0 0 $X=279540 $Y=99520
X3837 3 digital_ldo_top_VIA1 $T=279790 105200 0 0 $X=279540 $Y=104960
X3838 3 digital_ldo_top_VIA1 $T=279790 110640 0 0 $X=279540 $Y=110400
X3839 3 digital_ldo_top_VIA1 $T=279790 116080 0 0 $X=279540 $Y=115840
X3840 3 digital_ldo_top_VIA1 $T=279790 121520 0 0 $X=279540 $Y=121280
X3841 3 digital_ldo_top_VIA1 $T=279790 126960 0 0 $X=279540 $Y=126720
X3842 2 digital_ldo_top_VIA1 $T=281170 15440 0 0 $X=280920 $Y=15200
X3843 2 digital_ldo_top_VIA1 $T=281170 91600 0 0 $X=280920 $Y=91360
X3844 2 digital_ldo_top_VIA1 $T=281170 97040 0 0 $X=280920 $Y=96800
X3845 2 digital_ldo_top_VIA1 $T=281170 102480 0 0 $X=280920 $Y=102240
X3846 2 digital_ldo_top_VIA1 $T=281170 107920 0 0 $X=280920 $Y=107680
X3847 2 digital_ldo_top_VIA1 $T=281170 113360 0 0 $X=280920 $Y=113120
X3848 2 digital_ldo_top_VIA1 $T=281170 118800 0 0 $X=280920 $Y=118560
X3849 2 digital_ldo_top_VIA1 $T=281170 124240 0 0 $X=280920 $Y=124000
X3850 2 digital_ldo_top_VIA1 $T=281170 129680 0 0 $X=280920 $Y=129440
X3851 3 digital_ldo_top_VIA1 $T=283470 12720 0 0 $X=283220 $Y=12480
X3852 3 digital_ldo_top_VIA1 $T=283470 18160 0 0 $X=283220 $Y=17920
X3853 3 digital_ldo_top_VIA1 $T=283470 43160 0 0 $X=283220 $Y=42920
X3854 3 digital_ldo_top_VIA1 $T=283470 48600 0 0 $X=283220 $Y=48360
X3855 3 digital_ldo_top_VIA1 $T=283470 54040 0 0 $X=283220 $Y=53800
X3856 3 digital_ldo_top_VIA1 $T=283470 59480 0 0 $X=283220 $Y=59240
X3857 3 digital_ldo_top_VIA1 $T=283470 64920 0 0 $X=283220 $Y=64680
X3858 3 digital_ldo_top_VIA1 $T=283470 70360 0 0 $X=283220 $Y=70120
X3859 3 digital_ldo_top_VIA1 $T=283470 75800 0 0 $X=283220 $Y=75560
X3860 3 digital_ldo_top_VIA1 $T=283470 81240 0 0 $X=283220 $Y=81000
X3861 3 digital_ldo_top_VIA1 $T=283470 94320 0 0 $X=283220 $Y=94080
X3862 3 digital_ldo_top_VIA1 $T=283470 99760 0 0 $X=283220 $Y=99520
X3863 3 digital_ldo_top_VIA1 $T=283470 105200 0 0 $X=283220 $Y=104960
X3864 3 digital_ldo_top_VIA1 $T=283470 110640 0 0 $X=283220 $Y=110400
X3865 3 digital_ldo_top_VIA1 $T=283470 116080 0 0 $X=283220 $Y=115840
X3866 3 digital_ldo_top_VIA1 $T=283470 121520 0 0 $X=283220 $Y=121280
X3867 3 digital_ldo_top_VIA1 $T=283470 126960 0 0 $X=283220 $Y=126720
X3868 2 digital_ldo_top_VIA1 $T=284850 15440 0 0 $X=284600 $Y=15200
X3869 2 digital_ldo_top_VIA1 $T=284850 91600 0 0 $X=284600 $Y=91360
X3870 2 digital_ldo_top_VIA1 $T=284850 97040 0 0 $X=284600 $Y=96800
X3871 2 digital_ldo_top_VIA1 $T=284850 102480 0 0 $X=284600 $Y=102240
X3872 2 digital_ldo_top_VIA1 $T=284850 107920 0 0 $X=284600 $Y=107680
X3873 2 digital_ldo_top_VIA1 $T=284850 113360 0 0 $X=284600 $Y=113120
X3874 2 digital_ldo_top_VIA1 $T=284850 118800 0 0 $X=284600 $Y=118560
X3875 2 digital_ldo_top_VIA1 $T=284850 124240 0 0 $X=284600 $Y=124000
X3876 2 digital_ldo_top_VIA1 $T=284850 129680 0 0 $X=284600 $Y=129440
X3877 3 digital_ldo_top_VIA1 $T=287150 12720 0 0 $X=286900 $Y=12480
X3878 3 digital_ldo_top_VIA1 $T=287150 18160 0 0 $X=286900 $Y=17920
X3879 3 digital_ldo_top_VIA1 $T=287150 94320 0 0 $X=286900 $Y=94080
X3880 3 digital_ldo_top_VIA1 $T=287150 99760 0 0 $X=286900 $Y=99520
X3881 3 digital_ldo_top_VIA1 $T=287150 105200 0 0 $X=286900 $Y=104960
X3882 3 digital_ldo_top_VIA1 $T=287150 110640 0 0 $X=286900 $Y=110400
X3883 3 digital_ldo_top_VIA1 $T=287150 116080 0 0 $X=286900 $Y=115840
X3884 3 digital_ldo_top_VIA1 $T=287150 121520 0 0 $X=286900 $Y=121280
X3885 3 digital_ldo_top_VIA1 $T=287150 126960 0 0 $X=286900 $Y=126720
X3886 2 digital_ldo_top_VIA1 $T=288530 15440 0 0 $X=288280 $Y=15200
X3887 2 digital_ldo_top_VIA1 $T=288530 35000 0 0 $X=288280 $Y=34760
X3888 2 digital_ldo_top_VIA1 $T=288530 40440 0 0 $X=288280 $Y=40200
X3889 2 digital_ldo_top_VIA1 $T=288530 45880 0 0 $X=288280 $Y=45640
X3890 2 digital_ldo_top_VIA1 $T=288530 51320 0 0 $X=288280 $Y=51080
X3891 2 digital_ldo_top_VIA1 $T=288530 56760 0 0 $X=288280 $Y=56520
X3892 2 digital_ldo_top_VIA1 $T=288530 62200 0 0 $X=288280 $Y=61960
X3893 2 digital_ldo_top_VIA1 $T=288530 67640 0 0 $X=288280 $Y=67400
X3894 2 digital_ldo_top_VIA1 $T=288530 73080 0 0 $X=288280 $Y=72840
X3895 2 digital_ldo_top_VIA1 $T=288530 78520 0 0 $X=288280 $Y=78280
X3896 2 digital_ldo_top_VIA1 $T=288530 83960 0 0 $X=288280 $Y=83720
X3897 2 digital_ldo_top_VIA1 $T=288530 91600 0 0 $X=288280 $Y=91360
X3898 2 digital_ldo_top_VIA1 $T=288530 97040 0 0 $X=288280 $Y=96800
X3899 2 digital_ldo_top_VIA1 $T=288530 102480 0 0 $X=288280 $Y=102240
X3900 2 digital_ldo_top_VIA1 $T=288530 107920 0 0 $X=288280 $Y=107680
X3901 2 digital_ldo_top_VIA1 $T=288530 113360 0 0 $X=288280 $Y=113120
X3902 2 digital_ldo_top_VIA1 $T=288530 118800 0 0 $X=288280 $Y=118560
X3903 2 digital_ldo_top_VIA1 $T=288530 124240 0 0 $X=288280 $Y=124000
X3904 2 digital_ldo_top_VIA1 $T=288530 129680 0 0 $X=288280 $Y=129440
X3905 3 digital_ldo_top_VIA1 $T=290830 12720 0 0 $X=290580 $Y=12480
X3906 3 digital_ldo_top_VIA1 $T=290830 18160 0 0 $X=290580 $Y=17920
X3907 3 digital_ldo_top_VIA1 $T=290830 94320 0 0 $X=290580 $Y=94080
X3908 3 digital_ldo_top_VIA1 $T=290830 99760 0 0 $X=290580 $Y=99520
X3909 3 digital_ldo_top_VIA1 $T=290830 105200 0 0 $X=290580 $Y=104960
X3910 3 digital_ldo_top_VIA1 $T=290830 110640 0 0 $X=290580 $Y=110400
X3911 3 digital_ldo_top_VIA1 $T=290830 116080 0 0 $X=290580 $Y=115840
X3912 3 digital_ldo_top_VIA1 $T=290830 121520 0 0 $X=290580 $Y=121280
X3913 3 digital_ldo_top_VIA1 $T=290830 126960 0 0 $X=290580 $Y=126720
X3914 2 digital_ldo_top_VIA1 $T=292210 15440 0 0 $X=291960 $Y=15200
X3915 2 digital_ldo_top_VIA1 $T=292210 91600 0 0 $X=291960 $Y=91360
X3916 2 digital_ldo_top_VIA1 $T=292210 97040 0 0 $X=291960 $Y=96800
X3917 2 digital_ldo_top_VIA1 $T=292210 102480 0 0 $X=291960 $Y=102240
X3918 2 digital_ldo_top_VIA1 $T=292210 107920 0 0 $X=291960 $Y=107680
X3919 2 digital_ldo_top_VIA1 $T=292210 113360 0 0 $X=291960 $Y=113120
X3920 2 digital_ldo_top_VIA1 $T=292210 118800 0 0 $X=291960 $Y=118560
X3921 2 digital_ldo_top_VIA1 $T=292210 124240 0 0 $X=291960 $Y=124000
X3922 2 digital_ldo_top_VIA1 $T=292210 129680 0 0 $X=291960 $Y=129440
X3923 3 digital_ldo_top_VIA1 $T=294510 12720 0 0 $X=294260 $Y=12480
X3924 3 digital_ldo_top_VIA1 $T=294510 18160 0 0 $X=294260 $Y=17920
X3925 3 digital_ldo_top_VIA1 $T=294510 37720 0 0 $X=294260 $Y=37480
X3926 3 digital_ldo_top_VIA1 $T=294510 43160 0 0 $X=294260 $Y=42920
X3927 3 digital_ldo_top_VIA1 $T=294510 48600 0 0 $X=294260 $Y=48360
X3928 3 digital_ldo_top_VIA1 $T=294510 54040 0 0 $X=294260 $Y=53800
X3929 3 digital_ldo_top_VIA1 $T=294510 59480 0 0 $X=294260 $Y=59240
X3930 3 digital_ldo_top_VIA1 $T=294510 64920 0 0 $X=294260 $Y=64680
X3931 3 digital_ldo_top_VIA1 $T=294510 70360 0 0 $X=294260 $Y=70120
X3932 3 digital_ldo_top_VIA1 $T=294510 75800 0 0 $X=294260 $Y=75560
X3933 3 digital_ldo_top_VIA1 $T=294510 81240 0 0 $X=294260 $Y=81000
X3934 3 digital_ldo_top_VIA1 $T=294510 94320 0 0 $X=294260 $Y=94080
X3935 3 digital_ldo_top_VIA1 $T=294510 99760 0 0 $X=294260 $Y=99520
X3936 3 digital_ldo_top_VIA1 $T=294510 105200 0 0 $X=294260 $Y=104960
X3937 3 digital_ldo_top_VIA1 $T=294510 110640 0 0 $X=294260 $Y=110400
X3938 3 digital_ldo_top_VIA1 $T=294510 116080 0 0 $X=294260 $Y=115840
X3939 3 digital_ldo_top_VIA1 $T=294510 121520 0 0 $X=294260 $Y=121280
X3940 3 digital_ldo_top_VIA1 $T=294510 126960 0 0 $X=294260 $Y=126720
X3941 2 digital_ldo_top_VIA1 $T=295890 15440 0 0 $X=295640 $Y=15200
X3942 2 digital_ldo_top_VIA1 $T=295890 91600 0 0 $X=295640 $Y=91360
X3943 2 digital_ldo_top_VIA1 $T=295890 97040 0 0 $X=295640 $Y=96800
X3944 2 digital_ldo_top_VIA1 $T=295890 102480 0 0 $X=295640 $Y=102240
X3945 2 digital_ldo_top_VIA1 $T=295890 107920 0 0 $X=295640 $Y=107680
X3946 2 digital_ldo_top_VIA1 $T=295890 113360 0 0 $X=295640 $Y=113120
X3947 2 digital_ldo_top_VIA1 $T=295890 118800 0 0 $X=295640 $Y=118560
X3948 2 digital_ldo_top_VIA1 $T=295890 124240 0 0 $X=295640 $Y=124000
X3949 2 digital_ldo_top_VIA1 $T=295890 129680 0 0 $X=295640 $Y=129440
X3950 3 digital_ldo_top_VIA1 $T=298190 12720 0 0 $X=297940 $Y=12480
X3951 3 digital_ldo_top_VIA1 $T=298190 18160 0 0 $X=297940 $Y=17920
X3952 3 digital_ldo_top_VIA1 $T=298190 94320 0 0 $X=297940 $Y=94080
X3953 3 digital_ldo_top_VIA1 $T=298190 99760 0 0 $X=297940 $Y=99520
X3954 3 digital_ldo_top_VIA1 $T=298190 105200 0 0 $X=297940 $Y=104960
X3955 3 digital_ldo_top_VIA1 $T=298190 110640 0 0 $X=297940 $Y=110400
X3956 3 digital_ldo_top_VIA1 $T=298190 116080 0 0 $X=297940 $Y=115840
X3957 3 digital_ldo_top_VIA1 $T=298190 121520 0 0 $X=297940 $Y=121280
X3958 3 digital_ldo_top_VIA1 $T=298190 126960 0 0 $X=297940 $Y=126720
X3959 2 digital_ldo_top_VIA1 $T=299570 15440 0 0 $X=299320 $Y=15200
X3960 2 digital_ldo_top_VIA1 $T=299570 91600 0 0 $X=299320 $Y=91360
X3961 2 digital_ldo_top_VIA1 $T=299570 97040 0 0 $X=299320 $Y=96800
X3962 2 digital_ldo_top_VIA1 $T=299570 102480 0 0 $X=299320 $Y=102240
X3963 2 digital_ldo_top_VIA1 $T=299570 107920 0 0 $X=299320 $Y=107680
X3964 2 digital_ldo_top_VIA1 $T=299570 113360 0 0 $X=299320 $Y=113120
X3965 2 digital_ldo_top_VIA1 $T=299570 118800 0 0 $X=299320 $Y=118560
X3966 2 digital_ldo_top_VIA1 $T=299570 124240 0 0 $X=299320 $Y=124000
X3967 2 digital_ldo_top_VIA1 $T=299570 129680 0 0 $X=299320 $Y=129440
X3968 3 digital_ldo_top_VIA1 $T=301870 12720 0 0 $X=301620 $Y=12480
X3969 3 digital_ldo_top_VIA1 $T=301870 18160 0 0 $X=301620 $Y=17920
X3970 3 digital_ldo_top_VIA1 $T=301870 94320 0 0 $X=301620 $Y=94080
X3971 3 digital_ldo_top_VIA1 $T=301870 99760 0 0 $X=301620 $Y=99520
X3972 3 digital_ldo_top_VIA1 $T=301870 105200 0 0 $X=301620 $Y=104960
X3973 3 digital_ldo_top_VIA1 $T=301870 110640 0 0 $X=301620 $Y=110400
X3974 3 digital_ldo_top_VIA1 $T=301870 116080 0 0 $X=301620 $Y=115840
X3975 3 digital_ldo_top_VIA1 $T=301870 121520 0 0 $X=301620 $Y=121280
X3976 3 digital_ldo_top_VIA1 $T=301870 126960 0 0 $X=301620 $Y=126720
X3977 2 digital_ldo_top_VIA1 $T=303250 15440 0 0 $X=303000 $Y=15200
X3978 2 digital_ldo_top_VIA1 $T=303250 91600 0 0 $X=303000 $Y=91360
X3979 2 digital_ldo_top_VIA1 $T=303250 97040 0 0 $X=303000 $Y=96800
X3980 2 digital_ldo_top_VIA1 $T=303250 102480 0 0 $X=303000 $Y=102240
X3981 2 digital_ldo_top_VIA1 $T=303250 107920 0 0 $X=303000 $Y=107680
X3982 2 digital_ldo_top_VIA1 $T=303250 113360 0 0 $X=303000 $Y=113120
X3983 2 digital_ldo_top_VIA1 $T=303250 118800 0 0 $X=303000 $Y=118560
X3984 2 digital_ldo_top_VIA1 $T=303250 124240 0 0 $X=303000 $Y=124000
X3985 2 digital_ldo_top_VIA1 $T=303250 129680 0 0 $X=303000 $Y=129440
X3986 3 digital_ldo_top_VIA1 $T=305550 12720 0 0 $X=305300 $Y=12480
X3987 3 digital_ldo_top_VIA1 $T=305550 18160 0 0 $X=305300 $Y=17920
X3988 3 digital_ldo_top_VIA1 $T=305550 94320 0 0 $X=305300 $Y=94080
X3989 3 digital_ldo_top_VIA1 $T=305550 99760 0 0 $X=305300 $Y=99520
X3990 3 digital_ldo_top_VIA1 $T=305550 105200 0 0 $X=305300 $Y=104960
X3991 3 digital_ldo_top_VIA1 $T=305550 110640 0 0 $X=305300 $Y=110400
X3992 3 digital_ldo_top_VIA1 $T=305550 116080 0 0 $X=305300 $Y=115840
X3993 3 digital_ldo_top_VIA1 $T=305550 121520 0 0 $X=305300 $Y=121280
X3994 3 digital_ldo_top_VIA1 $T=305550 126960 0 0 $X=305300 $Y=126720
X3995 2 digital_ldo_top_VIA1 $T=306930 15440 0 0 $X=306680 $Y=15200
X3996 2 digital_ldo_top_VIA1 $T=306930 91600 0 0 $X=306680 $Y=91360
X3997 2 digital_ldo_top_VIA1 $T=306930 97040 0 0 $X=306680 $Y=96800
X3998 2 digital_ldo_top_VIA1 $T=306930 102480 0 0 $X=306680 $Y=102240
X3999 2 digital_ldo_top_VIA1 $T=306930 107920 0 0 $X=306680 $Y=107680
X4000 2 digital_ldo_top_VIA1 $T=306930 113360 0 0 $X=306680 $Y=113120
X4001 2 digital_ldo_top_VIA1 $T=306930 118800 0 0 $X=306680 $Y=118560
X4002 2 digital_ldo_top_VIA1 $T=306930 124240 0 0 $X=306680 $Y=124000
X4003 2 digital_ldo_top_VIA1 $T=306930 129680 0 0 $X=306680 $Y=129440
X4004 3 digital_ldo_top_VIA1 $T=309230 12720 0 0 $X=308980 $Y=12480
X4005 3 digital_ldo_top_VIA1 $T=309230 18160 0 0 $X=308980 $Y=17920
X4006 3 digital_ldo_top_VIA1 $T=309230 23600 0 0 $X=308980 $Y=23360
X4007 3 digital_ldo_top_VIA1 $T=309230 29040 0 0 $X=308980 $Y=28800
X4008 3 digital_ldo_top_VIA1 $T=309230 34480 0 0 $X=308980 $Y=34240
X4009 3 digital_ldo_top_VIA1 $T=309230 39920 0 0 $X=308980 $Y=39680
X4010 3 digital_ldo_top_VIA1 $T=309230 45360 0 0 $X=308980 $Y=45120
X4011 3 digital_ldo_top_VIA1 $T=309230 50800 0 0 $X=308980 $Y=50560
X4012 3 digital_ldo_top_VIA1 $T=309230 56240 0 0 $X=308980 $Y=56000
X4013 3 digital_ldo_top_VIA1 $T=309230 61680 0 0 $X=308980 $Y=61440
X4014 3 digital_ldo_top_VIA1 $T=309230 67120 0 0 $X=308980 $Y=66880
X4015 3 digital_ldo_top_VIA1 $T=309230 72560 0 0 $X=308980 $Y=72320
X4016 3 digital_ldo_top_VIA1 $T=309230 78000 0 0 $X=308980 $Y=77760
X4017 3 digital_ldo_top_VIA1 $T=309230 83440 0 0 $X=308980 $Y=83200
X4018 3 digital_ldo_top_VIA1 $T=309230 88880 0 0 $X=308980 $Y=88640
X4019 3 digital_ldo_top_VIA1 $T=309230 94320 0 0 $X=308980 $Y=94080
X4020 3 digital_ldo_top_VIA1 $T=309230 99760 0 0 $X=308980 $Y=99520
X4021 3 digital_ldo_top_VIA1 $T=309230 105200 0 0 $X=308980 $Y=104960
X4022 3 digital_ldo_top_VIA1 $T=309230 110640 0 0 $X=308980 $Y=110400
X4023 3 digital_ldo_top_VIA1 $T=309230 116080 0 0 $X=308980 $Y=115840
X4024 3 digital_ldo_top_VIA1 $T=309230 121520 0 0 $X=308980 $Y=121280
X4025 3 digital_ldo_top_VIA1 $T=309230 126960 0 0 $X=308980 $Y=126720
X4026 2 digital_ldo_top_VIA1 $T=310610 15440 0 0 $X=310360 $Y=15200
X4027 2 digital_ldo_top_VIA1 $T=310610 20880 0 0 $X=310360 $Y=20640
X4028 2 digital_ldo_top_VIA1 $T=310610 26320 0 0 $X=310360 $Y=26080
X4029 2 digital_ldo_top_VIA1 $T=310610 31760 0 0 $X=310360 $Y=31520
X4030 2 digital_ldo_top_VIA1 $T=310610 37200 0 0 $X=310360 $Y=36960
X4031 2 digital_ldo_top_VIA1 $T=310610 42640 0 0 $X=310360 $Y=42400
X4032 2 digital_ldo_top_VIA1 $T=310610 48080 0 0 $X=310360 $Y=47840
X4033 2 digital_ldo_top_VIA1 $T=310610 53520 0 0 $X=310360 $Y=53280
X4034 2 digital_ldo_top_VIA1 $T=310610 58960 0 0 $X=310360 $Y=58720
X4035 2 digital_ldo_top_VIA1 $T=310610 64400 0 0 $X=310360 $Y=64160
X4036 2 digital_ldo_top_VIA1 $T=310610 69840 0 0 $X=310360 $Y=69600
X4037 2 digital_ldo_top_VIA1 $T=310610 75280 0 0 $X=310360 $Y=75040
X4038 2 digital_ldo_top_VIA1 $T=310610 80720 0 0 $X=310360 $Y=80480
X4039 2 digital_ldo_top_VIA1 $T=310610 86160 0 0 $X=310360 $Y=85920
X4040 2 digital_ldo_top_VIA1 $T=310610 91600 0 0 $X=310360 $Y=91360
X4041 2 digital_ldo_top_VIA1 $T=310610 97040 0 0 $X=310360 $Y=96800
X4042 2 digital_ldo_top_VIA1 $T=310610 102480 0 0 $X=310360 $Y=102240
X4043 2 digital_ldo_top_VIA1 $T=310610 107920 0 0 $X=310360 $Y=107680
X4044 2 digital_ldo_top_VIA1 $T=310610 113360 0 0 $X=310360 $Y=113120
X4045 2 digital_ldo_top_VIA1 $T=310610 118800 0 0 $X=310360 $Y=118560
X4046 2 digital_ldo_top_VIA1 $T=310610 124240 0 0 $X=310360 $Y=124000
X4047 2 digital_ldo_top_VIA1 $T=310610 129680 0 0 $X=310360 $Y=129440
X4048 3 digital_ldo_top_VIA1 $T=312910 12720 0 0 $X=312660 $Y=12480
X4049 3 digital_ldo_top_VIA1 $T=312910 18160 0 0 $X=312660 $Y=17920
X4050 3 digital_ldo_top_VIA1 $T=312910 23600 0 0 $X=312660 $Y=23360
X4051 3 digital_ldo_top_VIA1 $T=312910 29040 0 0 $X=312660 $Y=28800
X4052 3 digital_ldo_top_VIA1 $T=312910 34480 0 0 $X=312660 $Y=34240
X4053 3 digital_ldo_top_VIA1 $T=312910 39920 0 0 $X=312660 $Y=39680
X4054 3 digital_ldo_top_VIA1 $T=312910 45360 0 0 $X=312660 $Y=45120
X4055 3 digital_ldo_top_VIA1 $T=312910 50800 0 0 $X=312660 $Y=50560
X4056 3 digital_ldo_top_VIA1 $T=312910 56240 0 0 $X=312660 $Y=56000
X4057 3 digital_ldo_top_VIA1 $T=312910 61680 0 0 $X=312660 $Y=61440
X4058 3 digital_ldo_top_VIA1 $T=312910 67120 0 0 $X=312660 $Y=66880
X4059 3 digital_ldo_top_VIA1 $T=312910 72560 0 0 $X=312660 $Y=72320
X4060 3 digital_ldo_top_VIA1 $T=312910 78000 0 0 $X=312660 $Y=77760
X4061 3 digital_ldo_top_VIA1 $T=312910 83440 0 0 $X=312660 $Y=83200
X4062 3 digital_ldo_top_VIA1 $T=312910 88880 0 0 $X=312660 $Y=88640
X4063 3 digital_ldo_top_VIA1 $T=312910 94320 0 0 $X=312660 $Y=94080
X4064 3 digital_ldo_top_VIA1 $T=312910 99760 0 0 $X=312660 $Y=99520
X4065 3 digital_ldo_top_VIA1 $T=312910 105200 0 0 $X=312660 $Y=104960
X4066 3 digital_ldo_top_VIA1 $T=312910 110640 0 0 $X=312660 $Y=110400
X4067 3 digital_ldo_top_VIA1 $T=312910 116080 0 0 $X=312660 $Y=115840
X4068 3 digital_ldo_top_VIA1 $T=312910 121520 0 0 $X=312660 $Y=121280
X4069 3 digital_ldo_top_VIA1 $T=312910 126960 0 0 $X=312660 $Y=126720
X4070 2 digital_ldo_top_VIA1 $T=314290 15440 0 0 $X=314040 $Y=15200
X4071 2 digital_ldo_top_VIA1 $T=314290 20880 0 0 $X=314040 $Y=20640
X4072 2 digital_ldo_top_VIA1 $T=314290 26320 0 0 $X=314040 $Y=26080
X4073 2 digital_ldo_top_VIA1 $T=314290 31760 0 0 $X=314040 $Y=31520
X4074 2 digital_ldo_top_VIA1 $T=314290 37200 0 0 $X=314040 $Y=36960
X4075 2 digital_ldo_top_VIA1 $T=314290 42640 0 0 $X=314040 $Y=42400
X4076 2 digital_ldo_top_VIA1 $T=314290 48080 0 0 $X=314040 $Y=47840
X4077 2 digital_ldo_top_VIA1 $T=314290 53520 0 0 $X=314040 $Y=53280
X4078 2 digital_ldo_top_VIA1 $T=314290 58960 0 0 $X=314040 $Y=58720
X4079 2 digital_ldo_top_VIA1 $T=314290 64400 0 0 $X=314040 $Y=64160
X4080 2 digital_ldo_top_VIA1 $T=314290 69840 0 0 $X=314040 $Y=69600
X4081 2 digital_ldo_top_VIA1 $T=314290 75280 0 0 $X=314040 $Y=75040
X4082 2 digital_ldo_top_VIA1 $T=314290 80720 0 0 $X=314040 $Y=80480
X4083 2 digital_ldo_top_VIA1 $T=314290 86160 0 0 $X=314040 $Y=85920
X4084 2 digital_ldo_top_VIA1 $T=314290 91600 0 0 $X=314040 $Y=91360
X4085 2 digital_ldo_top_VIA1 $T=314290 97040 0 0 $X=314040 $Y=96800
X4086 2 digital_ldo_top_VIA1 $T=314290 102480 0 0 $X=314040 $Y=102240
X4087 2 digital_ldo_top_VIA1 $T=314290 107920 0 0 $X=314040 $Y=107680
X4088 2 digital_ldo_top_VIA1 $T=314290 113360 0 0 $X=314040 $Y=113120
X4089 2 digital_ldo_top_VIA1 $T=314290 118800 0 0 $X=314040 $Y=118560
X4090 2 digital_ldo_top_VIA1 $T=314290 124240 0 0 $X=314040 $Y=124000
X4091 2 digital_ldo_top_VIA1 $T=314290 129680 0 0 $X=314040 $Y=129440
X4092 3 digital_ldo_top_VIA1 $T=316590 12720 0 0 $X=316340 $Y=12480
X4093 3 digital_ldo_top_VIA1 $T=316590 18160 0 0 $X=316340 $Y=17920
X4094 3 digital_ldo_top_VIA1 $T=316590 23600 0 0 $X=316340 $Y=23360
X4095 3 digital_ldo_top_VIA1 $T=316590 29040 0 0 $X=316340 $Y=28800
X4096 3 digital_ldo_top_VIA1 $T=316590 34480 0 0 $X=316340 $Y=34240
X4097 3 digital_ldo_top_VIA1 $T=316590 39920 0 0 $X=316340 $Y=39680
X4098 3 digital_ldo_top_VIA1 $T=316590 45360 0 0 $X=316340 $Y=45120
X4099 3 digital_ldo_top_VIA1 $T=316590 50800 0 0 $X=316340 $Y=50560
X4100 3 digital_ldo_top_VIA1 $T=316590 56240 0 0 $X=316340 $Y=56000
X4101 3 digital_ldo_top_VIA1 $T=316590 61680 0 0 $X=316340 $Y=61440
X4102 3 digital_ldo_top_VIA1 $T=316590 67120 0 0 $X=316340 $Y=66880
X4103 3 digital_ldo_top_VIA1 $T=316590 72560 0 0 $X=316340 $Y=72320
X4104 3 digital_ldo_top_VIA1 $T=316590 78000 0 0 $X=316340 $Y=77760
X4105 3 digital_ldo_top_VIA1 $T=316590 83440 0 0 $X=316340 $Y=83200
X4106 3 digital_ldo_top_VIA1 $T=316590 88880 0 0 $X=316340 $Y=88640
X4107 3 digital_ldo_top_VIA1 $T=316590 94320 0 0 $X=316340 $Y=94080
X4108 3 digital_ldo_top_VIA1 $T=316590 99760 0 0 $X=316340 $Y=99520
X4109 3 digital_ldo_top_VIA1 $T=316590 105200 0 0 $X=316340 $Y=104960
X4110 3 digital_ldo_top_VIA1 $T=316590 110640 0 0 $X=316340 $Y=110400
X4111 3 digital_ldo_top_VIA1 $T=316590 116080 0 0 $X=316340 $Y=115840
X4112 3 digital_ldo_top_VIA1 $T=316590 121520 0 0 $X=316340 $Y=121280
X4113 3 digital_ldo_top_VIA1 $T=316590 126960 0 0 $X=316340 $Y=126720
X4114 2 digital_ldo_top_VIA1 $T=317970 15440 0 0 $X=317720 $Y=15200
X4115 2 digital_ldo_top_VIA1 $T=317970 20880 0 0 $X=317720 $Y=20640
X4116 2 digital_ldo_top_VIA1 $T=317970 26320 0 0 $X=317720 $Y=26080
X4117 2 digital_ldo_top_VIA1 $T=317970 31760 0 0 $X=317720 $Y=31520
X4118 2 digital_ldo_top_VIA1 $T=317970 37200 0 0 $X=317720 $Y=36960
X4119 2 digital_ldo_top_VIA1 $T=317970 42640 0 0 $X=317720 $Y=42400
X4120 2 digital_ldo_top_VIA1 $T=317970 48080 0 0 $X=317720 $Y=47840
X4121 2 digital_ldo_top_VIA1 $T=317970 53520 0 0 $X=317720 $Y=53280
X4122 2 digital_ldo_top_VIA1 $T=317970 58960 0 0 $X=317720 $Y=58720
X4123 2 digital_ldo_top_VIA1 $T=317970 64400 0 0 $X=317720 $Y=64160
X4124 2 digital_ldo_top_VIA1 $T=317970 69840 0 0 $X=317720 $Y=69600
X4125 2 digital_ldo_top_VIA1 $T=317970 75280 0 0 $X=317720 $Y=75040
X4126 2 digital_ldo_top_VIA1 $T=317970 80720 0 0 $X=317720 $Y=80480
X4127 2 digital_ldo_top_VIA1 $T=317970 86160 0 0 $X=317720 $Y=85920
X4128 2 digital_ldo_top_VIA1 $T=317970 91600 0 0 $X=317720 $Y=91360
X4129 2 digital_ldo_top_VIA1 $T=317970 97040 0 0 $X=317720 $Y=96800
X4130 2 digital_ldo_top_VIA1 $T=317970 102480 0 0 $X=317720 $Y=102240
X4131 2 digital_ldo_top_VIA1 $T=317970 107920 0 0 $X=317720 $Y=107680
X4132 2 digital_ldo_top_VIA1 $T=317970 113360 0 0 $X=317720 $Y=113120
X4133 2 digital_ldo_top_VIA1 $T=317970 118800 0 0 $X=317720 $Y=118560
X4134 2 digital_ldo_top_VIA1 $T=317970 124240 0 0 $X=317720 $Y=124000
X4135 2 digital_ldo_top_VIA1 $T=317970 129680 0 0 $X=317720 $Y=129440
X4136 3 digital_ldo_top_VIA1 $T=320270 12720 0 0 $X=320020 $Y=12480
X4137 3 digital_ldo_top_VIA1 $T=320270 18160 0 0 $X=320020 $Y=17920
X4138 3 digital_ldo_top_VIA1 $T=320270 23600 0 0 $X=320020 $Y=23360
X4139 3 digital_ldo_top_VIA1 $T=320270 29040 0 0 $X=320020 $Y=28800
X4140 3 digital_ldo_top_VIA1 $T=320270 34480 0 0 $X=320020 $Y=34240
X4141 3 digital_ldo_top_VIA1 $T=320270 39920 0 0 $X=320020 $Y=39680
X4142 3 digital_ldo_top_VIA1 $T=320270 45360 0 0 $X=320020 $Y=45120
X4143 3 digital_ldo_top_VIA1 $T=320270 50800 0 0 $X=320020 $Y=50560
X4144 3 digital_ldo_top_VIA1 $T=320270 56240 0 0 $X=320020 $Y=56000
X4145 3 digital_ldo_top_VIA1 $T=320270 61680 0 0 $X=320020 $Y=61440
X4146 3 digital_ldo_top_VIA1 $T=320270 67120 0 0 $X=320020 $Y=66880
X4147 3 digital_ldo_top_VIA1 $T=320270 72560 0 0 $X=320020 $Y=72320
X4148 3 digital_ldo_top_VIA1 $T=320270 78000 0 0 $X=320020 $Y=77760
X4149 3 digital_ldo_top_VIA1 $T=320270 83440 0 0 $X=320020 $Y=83200
X4150 3 digital_ldo_top_VIA1 $T=320270 88880 0 0 $X=320020 $Y=88640
X4151 3 digital_ldo_top_VIA1 $T=320270 94320 0 0 $X=320020 $Y=94080
X4152 3 digital_ldo_top_VIA1 $T=320270 99760 0 0 $X=320020 $Y=99520
X4153 3 digital_ldo_top_VIA1 $T=320270 105200 0 0 $X=320020 $Y=104960
X4154 3 digital_ldo_top_VIA1 $T=320270 110640 0 0 $X=320020 $Y=110400
X4155 3 digital_ldo_top_VIA1 $T=320270 116080 0 0 $X=320020 $Y=115840
X4156 3 digital_ldo_top_VIA1 $T=320270 121520 0 0 $X=320020 $Y=121280
X4157 3 digital_ldo_top_VIA1 $T=320270 126960 0 0 $X=320020 $Y=126720
X4158 2 digital_ldo_top_VIA1 $T=321650 15440 0 0 $X=321400 $Y=15200
X4159 2 digital_ldo_top_VIA1 $T=321650 20880 0 0 $X=321400 $Y=20640
X4160 2 digital_ldo_top_VIA1 $T=321650 26320 0 0 $X=321400 $Y=26080
X4161 2 digital_ldo_top_VIA1 $T=321650 31760 0 0 $X=321400 $Y=31520
X4162 2 digital_ldo_top_VIA1 $T=321650 37200 0 0 $X=321400 $Y=36960
X4163 2 digital_ldo_top_VIA1 $T=321650 42640 0 0 $X=321400 $Y=42400
X4164 2 digital_ldo_top_VIA1 $T=321650 48080 0 0 $X=321400 $Y=47840
X4165 2 digital_ldo_top_VIA1 $T=321650 53520 0 0 $X=321400 $Y=53280
X4166 2 digital_ldo_top_VIA1 $T=321650 58960 0 0 $X=321400 $Y=58720
X4167 2 digital_ldo_top_VIA1 $T=321650 64400 0 0 $X=321400 $Y=64160
X4168 2 digital_ldo_top_VIA1 $T=321650 69840 0 0 $X=321400 $Y=69600
X4169 2 digital_ldo_top_VIA1 $T=321650 75280 0 0 $X=321400 $Y=75040
X4170 2 digital_ldo_top_VIA1 $T=321650 80720 0 0 $X=321400 $Y=80480
X4171 2 digital_ldo_top_VIA1 $T=321650 86160 0 0 $X=321400 $Y=85920
X4172 2 digital_ldo_top_VIA1 $T=321650 91600 0 0 $X=321400 $Y=91360
X4173 2 digital_ldo_top_VIA1 $T=321650 97040 0 0 $X=321400 $Y=96800
X4174 2 digital_ldo_top_VIA1 $T=321650 102480 0 0 $X=321400 $Y=102240
X4175 2 digital_ldo_top_VIA1 $T=321650 107920 0 0 $X=321400 $Y=107680
X4176 2 digital_ldo_top_VIA1 $T=321650 113360 0 0 $X=321400 $Y=113120
X4177 2 digital_ldo_top_VIA1 $T=321650 118800 0 0 $X=321400 $Y=118560
X4178 2 digital_ldo_top_VIA1 $T=321650 124240 0 0 $X=321400 $Y=124000
X4179 2 digital_ldo_top_VIA1 $T=321650 129680 0 0 $X=321400 $Y=129440
X4180 3 digital_ldo_top_VIA1 $T=323950 12720 0 0 $X=323700 $Y=12480
X4181 3 digital_ldo_top_VIA1 $T=323950 50800 0 0 $X=323700 $Y=50560
X4182 3 digital_ldo_top_VIA1 $T=323950 56240 0 0 $X=323700 $Y=56000
X4183 3 digital_ldo_top_VIA1 $T=323950 61680 0 0 $X=323700 $Y=61440
X4184 3 digital_ldo_top_VIA1 $T=323950 67120 0 0 $X=323700 $Y=66880
X4185 3 digital_ldo_top_VIA1 $T=323950 72560 0 0 $X=323700 $Y=72320
X4186 3 digital_ldo_top_VIA1 $T=323950 78000 0 0 $X=323700 $Y=77760
X4187 3 digital_ldo_top_VIA1 $T=323950 83440 0 0 $X=323700 $Y=83200
X4188 3 digital_ldo_top_VIA1 $T=323950 88880 0 0 $X=323700 $Y=88640
X4189 3 digital_ldo_top_VIA1 $T=323950 94320 0 0 $X=323700 $Y=94080
X4190 3 digital_ldo_top_VIA1 $T=323950 99760 0 0 $X=323700 $Y=99520
X4191 3 digital_ldo_top_VIA1 $T=323950 105200 0 0 $X=323700 $Y=104960
X4192 3 digital_ldo_top_VIA1 $T=323950 110640 0 0 $X=323700 $Y=110400
X4193 3 digital_ldo_top_VIA1 $T=323950 116080 0 0 $X=323700 $Y=115840
X4194 3 digital_ldo_top_VIA1 $T=323950 121520 0 0 $X=323700 $Y=121280
X4195 3 digital_ldo_top_VIA1 $T=323950 126960 0 0 $X=323700 $Y=126720
X4196 2 digital_ldo_top_VIA1 $T=325330 53520 0 0 $X=325080 $Y=53280
X4197 2 digital_ldo_top_VIA1 $T=325330 58960 0 0 $X=325080 $Y=58720
X4198 2 digital_ldo_top_VIA1 $T=325330 64400 0 0 $X=325080 $Y=64160
X4199 2 digital_ldo_top_VIA1 $T=325330 69840 0 0 $X=325080 $Y=69600
X4200 2 digital_ldo_top_VIA1 $T=325330 75280 0 0 $X=325080 $Y=75040
X4201 2 digital_ldo_top_VIA1 $T=325330 80720 0 0 $X=325080 $Y=80480
X4202 2 digital_ldo_top_VIA1 $T=325330 86160 0 0 $X=325080 $Y=85920
X4203 2 digital_ldo_top_VIA1 $T=325330 91600 0 0 $X=325080 $Y=91360
X4204 2 digital_ldo_top_VIA1 $T=325330 97040 0 0 $X=325080 $Y=96800
X4205 2 digital_ldo_top_VIA1 $T=325330 102480 0 0 $X=325080 $Y=102240
X4206 2 digital_ldo_top_VIA1 $T=325330 107920 0 0 $X=325080 $Y=107680
X4207 2 digital_ldo_top_VIA1 $T=325330 113360 0 0 $X=325080 $Y=113120
X4208 2 digital_ldo_top_VIA1 $T=325330 118800 0 0 $X=325080 $Y=118560
X4209 2 digital_ldo_top_VIA1 $T=325330 124240 0 0 $X=325080 $Y=124000
X4210 2 digital_ldo_top_VIA1 $T=325330 129680 0 0 $X=325080 $Y=129440
X4211 3 digital_ldo_top_VIA1 $T=327630 12720 0 0 $X=327380 $Y=12480
X4212 3 digital_ldo_top_VIA1 $T=327630 50800 0 0 $X=327380 $Y=50560
X4213 3 digital_ldo_top_VIA1 $T=327630 56240 0 0 $X=327380 $Y=56000
X4214 3 digital_ldo_top_VIA1 $T=327630 61680 0 0 $X=327380 $Y=61440
X4215 3 digital_ldo_top_VIA1 $T=327630 67120 0 0 $X=327380 $Y=66880
X4216 3 digital_ldo_top_VIA1 $T=327630 72560 0 0 $X=327380 $Y=72320
X4217 3 digital_ldo_top_VIA1 $T=327630 78000 0 0 $X=327380 $Y=77760
X4218 3 digital_ldo_top_VIA1 $T=327630 83440 0 0 $X=327380 $Y=83200
X4219 3 digital_ldo_top_VIA1 $T=327630 88880 0 0 $X=327380 $Y=88640
X4220 3 digital_ldo_top_VIA1 $T=327630 94320 0 0 $X=327380 $Y=94080
X4221 3 digital_ldo_top_VIA1 $T=327630 99760 0 0 $X=327380 $Y=99520
X4222 3 digital_ldo_top_VIA1 $T=327630 105200 0 0 $X=327380 $Y=104960
X4223 3 digital_ldo_top_VIA1 $T=327630 110640 0 0 $X=327380 $Y=110400
X4224 3 digital_ldo_top_VIA1 $T=327630 116080 0 0 $X=327380 $Y=115840
X4225 3 digital_ldo_top_VIA1 $T=327630 121520 0 0 $X=327380 $Y=121280
X4226 3 digital_ldo_top_VIA1 $T=327630 126960 0 0 $X=327380 $Y=126720
X4227 2 digital_ldo_top_VIA1 $T=329010 53520 0 0 $X=328760 $Y=53280
X4228 2 digital_ldo_top_VIA1 $T=329010 58960 0 0 $X=328760 $Y=58720
X4229 2 digital_ldo_top_VIA1 $T=329010 64400 0 0 $X=328760 $Y=64160
X4230 2 digital_ldo_top_VIA1 $T=329010 69840 0 0 $X=328760 $Y=69600
X4231 2 digital_ldo_top_VIA1 $T=329010 75280 0 0 $X=328760 $Y=75040
X4232 2 digital_ldo_top_VIA1 $T=329010 80720 0 0 $X=328760 $Y=80480
X4233 2 digital_ldo_top_VIA1 $T=329010 86160 0 0 $X=328760 $Y=85920
X4234 2 digital_ldo_top_VIA1 $T=329010 91600 0 0 $X=328760 $Y=91360
X4235 2 digital_ldo_top_VIA1 $T=329010 97040 0 0 $X=328760 $Y=96800
X4236 2 digital_ldo_top_VIA1 $T=329010 102480 0 0 $X=328760 $Y=102240
X4237 2 digital_ldo_top_VIA1 $T=329010 107920 0 0 $X=328760 $Y=107680
X4238 2 digital_ldo_top_VIA1 $T=329010 113360 0 0 $X=328760 $Y=113120
X4239 2 digital_ldo_top_VIA1 $T=329010 118800 0 0 $X=328760 $Y=118560
X4240 2 digital_ldo_top_VIA1 $T=329010 124240 0 0 $X=328760 $Y=124000
X4241 2 digital_ldo_top_VIA1 $T=329010 129680 0 0 $X=328760 $Y=129440
X4242 3 digital_ldo_top_VIA1 $T=331310 12720 0 0 $X=331060 $Y=12480
X4243 3 digital_ldo_top_VIA1 $T=331310 50800 0 0 $X=331060 $Y=50560
X4244 3 digital_ldo_top_VIA1 $T=331310 56240 0 0 $X=331060 $Y=56000
X4245 3 digital_ldo_top_VIA1 $T=331310 61680 0 0 $X=331060 $Y=61440
X4246 3 digital_ldo_top_VIA1 $T=331310 67120 0 0 $X=331060 $Y=66880
X4247 3 digital_ldo_top_VIA1 $T=331310 72560 0 0 $X=331060 $Y=72320
X4248 3 digital_ldo_top_VIA1 $T=331310 78000 0 0 $X=331060 $Y=77760
X4249 3 digital_ldo_top_VIA1 $T=331310 83440 0 0 $X=331060 $Y=83200
X4250 3 digital_ldo_top_VIA1 $T=331310 88880 0 0 $X=331060 $Y=88640
X4251 3 digital_ldo_top_VIA1 $T=331310 94320 0 0 $X=331060 $Y=94080
X4252 3 digital_ldo_top_VIA1 $T=331310 99760 0 0 $X=331060 $Y=99520
X4253 3 digital_ldo_top_VIA1 $T=331310 105200 0 0 $X=331060 $Y=104960
X4254 3 digital_ldo_top_VIA1 $T=331310 110640 0 0 $X=331060 $Y=110400
X4255 3 digital_ldo_top_VIA1 $T=331310 116080 0 0 $X=331060 $Y=115840
X4256 3 digital_ldo_top_VIA1 $T=331310 121520 0 0 $X=331060 $Y=121280
X4257 3 digital_ldo_top_VIA1 $T=331310 126960 0 0 $X=331060 $Y=126720
X4258 2 digital_ldo_top_VIA1 $T=332690 53520 0 0 $X=332440 $Y=53280
X4259 2 digital_ldo_top_VIA1 $T=332690 58960 0 0 $X=332440 $Y=58720
X4260 2 digital_ldo_top_VIA1 $T=332690 64400 0 0 $X=332440 $Y=64160
X4261 2 digital_ldo_top_VIA1 $T=332690 69840 0 0 $X=332440 $Y=69600
X4262 2 digital_ldo_top_VIA1 $T=332690 75280 0 0 $X=332440 $Y=75040
X4263 2 digital_ldo_top_VIA1 $T=332690 80720 0 0 $X=332440 $Y=80480
X4264 2 digital_ldo_top_VIA1 $T=332690 86160 0 0 $X=332440 $Y=85920
X4265 2 digital_ldo_top_VIA1 $T=332690 91600 0 0 $X=332440 $Y=91360
X4266 2 digital_ldo_top_VIA1 $T=332690 97040 0 0 $X=332440 $Y=96800
X4267 2 digital_ldo_top_VIA1 $T=332690 102480 0 0 $X=332440 $Y=102240
X4268 2 digital_ldo_top_VIA1 $T=332690 107920 0 0 $X=332440 $Y=107680
X4269 2 digital_ldo_top_VIA1 $T=332690 113360 0 0 $X=332440 $Y=113120
X4270 2 digital_ldo_top_VIA1 $T=332690 118800 0 0 $X=332440 $Y=118560
X4271 2 digital_ldo_top_VIA1 $T=332690 124240 0 0 $X=332440 $Y=124000
X4272 2 digital_ldo_top_VIA1 $T=332690 129680 0 0 $X=332440 $Y=129440
X4273 3 digital_ldo_top_VIA1 $T=334990 12720 0 0 $X=334740 $Y=12480
X4274 3 digital_ldo_top_VIA1 $T=334990 50800 0 0 $X=334740 $Y=50560
X4275 3 digital_ldo_top_VIA1 $T=334990 56240 0 0 $X=334740 $Y=56000
X4276 3 digital_ldo_top_VIA1 $T=334990 61680 0 0 $X=334740 $Y=61440
X4277 3 digital_ldo_top_VIA1 $T=334990 67120 0 0 $X=334740 $Y=66880
X4278 3 digital_ldo_top_VIA1 $T=334990 72560 0 0 $X=334740 $Y=72320
X4279 3 digital_ldo_top_VIA1 $T=334990 78000 0 0 $X=334740 $Y=77760
X4280 3 digital_ldo_top_VIA1 $T=334990 83440 0 0 $X=334740 $Y=83200
X4281 3 digital_ldo_top_VIA1 $T=334990 88880 0 0 $X=334740 $Y=88640
X4282 3 digital_ldo_top_VIA1 $T=334990 94320 0 0 $X=334740 $Y=94080
X4283 3 digital_ldo_top_VIA1 $T=334990 99760 0 0 $X=334740 $Y=99520
X4284 3 digital_ldo_top_VIA1 $T=334990 105200 0 0 $X=334740 $Y=104960
X4285 3 digital_ldo_top_VIA1 $T=334990 110640 0 0 $X=334740 $Y=110400
X4286 3 digital_ldo_top_VIA1 $T=334990 116080 0 0 $X=334740 $Y=115840
X4287 3 digital_ldo_top_VIA1 $T=334990 121520 0 0 $X=334740 $Y=121280
X4288 3 digital_ldo_top_VIA1 $T=334990 126960 0 0 $X=334740 $Y=126720
X4289 2 digital_ldo_top_VIA1 $T=336370 53520 0 0 $X=336120 $Y=53280
X4290 2 digital_ldo_top_VIA1 $T=336370 58960 0 0 $X=336120 $Y=58720
X4291 2 digital_ldo_top_VIA1 $T=336370 64400 0 0 $X=336120 $Y=64160
X4292 2 digital_ldo_top_VIA1 $T=336370 69840 0 0 $X=336120 $Y=69600
X4293 2 digital_ldo_top_VIA1 $T=336370 75280 0 0 $X=336120 $Y=75040
X4294 2 digital_ldo_top_VIA1 $T=336370 80720 0 0 $X=336120 $Y=80480
X4295 2 digital_ldo_top_VIA1 $T=336370 86160 0 0 $X=336120 $Y=85920
X4296 2 digital_ldo_top_VIA1 $T=336370 91600 0 0 $X=336120 $Y=91360
X4297 2 digital_ldo_top_VIA1 $T=336370 97040 0 0 $X=336120 $Y=96800
X4298 2 digital_ldo_top_VIA1 $T=336370 102480 0 0 $X=336120 $Y=102240
X4299 2 digital_ldo_top_VIA1 $T=336370 107920 0 0 $X=336120 $Y=107680
X4300 2 digital_ldo_top_VIA1 $T=336370 113360 0 0 $X=336120 $Y=113120
X4301 2 digital_ldo_top_VIA1 $T=336370 118800 0 0 $X=336120 $Y=118560
X4302 2 digital_ldo_top_VIA1 $T=336370 124240 0 0 $X=336120 $Y=124000
X4303 2 digital_ldo_top_VIA1 $T=336370 129680 0 0 $X=336120 $Y=129440
X4304 3 digital_ldo_top_VIA1 $T=338670 12720 0 0 $X=338420 $Y=12480
X4305 3 digital_ldo_top_VIA1 $T=338670 50800 0 0 $X=338420 $Y=50560
X4306 3 digital_ldo_top_VIA1 $T=338670 56240 0 0 $X=338420 $Y=56000
X4307 3 digital_ldo_top_VIA1 $T=338670 61680 0 0 $X=338420 $Y=61440
X4308 3 digital_ldo_top_VIA1 $T=338670 67120 0 0 $X=338420 $Y=66880
X4309 3 digital_ldo_top_VIA1 $T=338670 72560 0 0 $X=338420 $Y=72320
X4310 3 digital_ldo_top_VIA1 $T=338670 78000 0 0 $X=338420 $Y=77760
X4311 3 digital_ldo_top_VIA1 $T=338670 83440 0 0 $X=338420 $Y=83200
X4312 3 digital_ldo_top_VIA1 $T=338670 88880 0 0 $X=338420 $Y=88640
X4313 3 digital_ldo_top_VIA1 $T=338670 94320 0 0 $X=338420 $Y=94080
X4314 3 digital_ldo_top_VIA1 $T=338670 99760 0 0 $X=338420 $Y=99520
X4315 3 digital_ldo_top_VIA1 $T=338670 105200 0 0 $X=338420 $Y=104960
X4316 3 digital_ldo_top_VIA1 $T=338670 110640 0 0 $X=338420 $Y=110400
X4317 3 digital_ldo_top_VIA1 $T=338670 116080 0 0 $X=338420 $Y=115840
X4318 3 digital_ldo_top_VIA1 $T=338670 121520 0 0 $X=338420 $Y=121280
X4319 3 digital_ldo_top_VIA1 $T=338670 126960 0 0 $X=338420 $Y=126720
X4320 2 digital_ldo_top_VIA1 $T=340050 53520 0 0 $X=339800 $Y=53280
X4321 2 digital_ldo_top_VIA1 $T=340050 58960 0 0 $X=339800 $Y=58720
X4322 2 digital_ldo_top_VIA1 $T=340050 64400 0 0 $X=339800 $Y=64160
X4323 2 digital_ldo_top_VIA1 $T=340050 69840 0 0 $X=339800 $Y=69600
X4324 2 digital_ldo_top_VIA1 $T=340050 75280 0 0 $X=339800 $Y=75040
X4325 2 digital_ldo_top_VIA1 $T=340050 80720 0 0 $X=339800 $Y=80480
X4326 2 digital_ldo_top_VIA1 $T=340050 86160 0 0 $X=339800 $Y=85920
X4327 2 digital_ldo_top_VIA1 $T=340050 91600 0 0 $X=339800 $Y=91360
X4328 2 digital_ldo_top_VIA1 $T=340050 97040 0 0 $X=339800 $Y=96800
X4329 2 digital_ldo_top_VIA1 $T=340050 102480 0 0 $X=339800 $Y=102240
X4330 2 digital_ldo_top_VIA1 $T=340050 107920 0 0 $X=339800 $Y=107680
X4331 2 digital_ldo_top_VIA1 $T=340050 113360 0 0 $X=339800 $Y=113120
X4332 2 digital_ldo_top_VIA1 $T=340050 118800 0 0 $X=339800 $Y=118560
X4333 2 digital_ldo_top_VIA1 $T=340050 124240 0 0 $X=339800 $Y=124000
X4334 2 digital_ldo_top_VIA1 $T=340050 129680 0 0 $X=339800 $Y=129440
X4335 3 digital_ldo_top_VIA1 $T=342350 12720 0 0 $X=342100 $Y=12480
X4336 3 digital_ldo_top_VIA1 $T=342350 50800 0 0 $X=342100 $Y=50560
X4337 3 digital_ldo_top_VIA1 $T=342350 56240 0 0 $X=342100 $Y=56000
X4338 3 digital_ldo_top_VIA1 $T=342350 61680 0 0 $X=342100 $Y=61440
X4339 3 digital_ldo_top_VIA1 $T=342350 67120 0 0 $X=342100 $Y=66880
X4340 3 digital_ldo_top_VIA1 $T=342350 72560 0 0 $X=342100 $Y=72320
X4341 3 digital_ldo_top_VIA1 $T=342350 78000 0 0 $X=342100 $Y=77760
X4342 3 digital_ldo_top_VIA1 $T=342350 83440 0 0 $X=342100 $Y=83200
X4343 3 digital_ldo_top_VIA1 $T=342350 88880 0 0 $X=342100 $Y=88640
X4344 3 digital_ldo_top_VIA1 $T=342350 94320 0 0 $X=342100 $Y=94080
X4345 3 digital_ldo_top_VIA1 $T=342350 99760 0 0 $X=342100 $Y=99520
X4346 3 digital_ldo_top_VIA1 $T=342350 105200 0 0 $X=342100 $Y=104960
X4347 3 digital_ldo_top_VIA1 $T=342350 110640 0 0 $X=342100 $Y=110400
X4348 3 digital_ldo_top_VIA1 $T=342350 116080 0 0 $X=342100 $Y=115840
X4349 3 digital_ldo_top_VIA1 $T=342350 121520 0 0 $X=342100 $Y=121280
X4350 3 digital_ldo_top_VIA1 $T=342350 126960 0 0 $X=342100 $Y=126720
X4351 2 digital_ldo_top_VIA1 $T=343730 53520 0 0 $X=343480 $Y=53280
X4352 2 digital_ldo_top_VIA1 $T=343730 58960 0 0 $X=343480 $Y=58720
X4353 2 digital_ldo_top_VIA1 $T=343730 64400 0 0 $X=343480 $Y=64160
X4354 2 digital_ldo_top_VIA1 $T=343730 69840 0 0 $X=343480 $Y=69600
X4355 2 digital_ldo_top_VIA1 $T=343730 75280 0 0 $X=343480 $Y=75040
X4356 2 digital_ldo_top_VIA1 $T=343730 80720 0 0 $X=343480 $Y=80480
X4357 2 digital_ldo_top_VIA1 $T=343730 86160 0 0 $X=343480 $Y=85920
X4358 2 digital_ldo_top_VIA1 $T=343730 91600 0 0 $X=343480 $Y=91360
X4359 2 digital_ldo_top_VIA1 $T=343730 97040 0 0 $X=343480 $Y=96800
X4360 2 digital_ldo_top_VIA1 $T=343730 102480 0 0 $X=343480 $Y=102240
X4361 2 digital_ldo_top_VIA1 $T=343730 107920 0 0 $X=343480 $Y=107680
X4362 2 digital_ldo_top_VIA1 $T=343730 113360 0 0 $X=343480 $Y=113120
X4363 2 digital_ldo_top_VIA1 $T=343730 118800 0 0 $X=343480 $Y=118560
X4364 2 digital_ldo_top_VIA1 $T=343730 124240 0 0 $X=343480 $Y=124000
X4365 2 digital_ldo_top_VIA1 $T=343730 129680 0 0 $X=343480 $Y=129440
X4366 3 digital_ldo_top_VIA1 $T=346030 12720 0 0 $X=345780 $Y=12480
X4367 3 digital_ldo_top_VIA1 $T=346030 50800 0 0 $X=345780 $Y=50560
X4368 3 digital_ldo_top_VIA1 $T=346030 56240 0 0 $X=345780 $Y=56000
X4369 3 digital_ldo_top_VIA1 $T=346030 61680 0 0 $X=345780 $Y=61440
X4370 3 digital_ldo_top_VIA1 $T=346030 67120 0 0 $X=345780 $Y=66880
X4371 3 digital_ldo_top_VIA1 $T=346030 72560 0 0 $X=345780 $Y=72320
X4372 3 digital_ldo_top_VIA1 $T=346030 78000 0 0 $X=345780 $Y=77760
X4373 3 digital_ldo_top_VIA1 $T=346030 83440 0 0 $X=345780 $Y=83200
X4374 3 digital_ldo_top_VIA1 $T=346030 88880 0 0 $X=345780 $Y=88640
X4375 3 digital_ldo_top_VIA1 $T=346030 94320 0 0 $X=345780 $Y=94080
X4376 3 digital_ldo_top_VIA1 $T=346030 99760 0 0 $X=345780 $Y=99520
X4377 3 digital_ldo_top_VIA1 $T=346030 105200 0 0 $X=345780 $Y=104960
X4378 3 digital_ldo_top_VIA1 $T=346030 110640 0 0 $X=345780 $Y=110400
X4379 3 digital_ldo_top_VIA1 $T=346030 116080 0 0 $X=345780 $Y=115840
X4380 3 digital_ldo_top_VIA1 $T=346030 121520 0 0 $X=345780 $Y=121280
X4381 3 digital_ldo_top_VIA1 $T=346030 126960 0 0 $X=345780 $Y=126720
X4382 2 digital_ldo_top_VIA1 $T=347410 53520 0 0 $X=347160 $Y=53280
X4383 2 digital_ldo_top_VIA1 $T=347410 58960 0 0 $X=347160 $Y=58720
X4384 2 digital_ldo_top_VIA1 $T=347410 64400 0 0 $X=347160 $Y=64160
X4385 2 digital_ldo_top_VIA1 $T=347410 69840 0 0 $X=347160 $Y=69600
X4386 2 digital_ldo_top_VIA1 $T=347410 75280 0 0 $X=347160 $Y=75040
X4387 2 digital_ldo_top_VIA1 $T=347410 80720 0 0 $X=347160 $Y=80480
X4388 2 digital_ldo_top_VIA1 $T=347410 86160 0 0 $X=347160 $Y=85920
X4389 2 digital_ldo_top_VIA1 $T=347410 91600 0 0 $X=347160 $Y=91360
X4390 2 digital_ldo_top_VIA1 $T=347410 97040 0 0 $X=347160 $Y=96800
X4391 2 digital_ldo_top_VIA1 $T=347410 102480 0 0 $X=347160 $Y=102240
X4392 2 digital_ldo_top_VIA1 $T=347410 107920 0 0 $X=347160 $Y=107680
X4393 2 digital_ldo_top_VIA1 $T=347410 113360 0 0 $X=347160 $Y=113120
X4394 2 digital_ldo_top_VIA1 $T=347410 118800 0 0 $X=347160 $Y=118560
X4395 2 digital_ldo_top_VIA1 $T=347410 124240 0 0 $X=347160 $Y=124000
X4396 2 digital_ldo_top_VIA1 $T=347410 129680 0 0 $X=347160 $Y=129440
X4397 3 digital_ldo_top_VIA1 $T=349710 12720 0 0 $X=349460 $Y=12480
X4398 3 digital_ldo_top_VIA1 $T=349710 50800 0 0 $X=349460 $Y=50560
X4399 3 digital_ldo_top_VIA1 $T=349710 56240 0 0 $X=349460 $Y=56000
X4400 3 digital_ldo_top_VIA1 $T=349710 61680 0 0 $X=349460 $Y=61440
X4401 3 digital_ldo_top_VIA1 $T=349710 67120 0 0 $X=349460 $Y=66880
X4402 3 digital_ldo_top_VIA1 $T=349710 72560 0 0 $X=349460 $Y=72320
X4403 3 digital_ldo_top_VIA1 $T=349710 78000 0 0 $X=349460 $Y=77760
X4404 3 digital_ldo_top_VIA1 $T=349710 83440 0 0 $X=349460 $Y=83200
X4405 3 digital_ldo_top_VIA1 $T=349710 88880 0 0 $X=349460 $Y=88640
X4406 3 digital_ldo_top_VIA1 $T=349710 94320 0 0 $X=349460 $Y=94080
X4407 3 digital_ldo_top_VIA1 $T=349710 99760 0 0 $X=349460 $Y=99520
X4408 3 digital_ldo_top_VIA1 $T=349710 105200 0 0 $X=349460 $Y=104960
X4409 3 digital_ldo_top_VIA1 $T=349710 110640 0 0 $X=349460 $Y=110400
X4410 3 digital_ldo_top_VIA1 $T=349710 116080 0 0 $X=349460 $Y=115840
X4411 3 digital_ldo_top_VIA1 $T=349710 121520 0 0 $X=349460 $Y=121280
X4412 3 digital_ldo_top_VIA1 $T=349710 126960 0 0 $X=349460 $Y=126720
X4413 2 digital_ldo_top_VIA1 $T=351090 15440 0 0 $X=350840 $Y=15200
X4414 2 digital_ldo_top_VIA1 $T=351090 20880 0 0 $X=350840 $Y=20640
X4415 2 digital_ldo_top_VIA1 $T=351090 26320 0 0 $X=350840 $Y=26080
X4416 2 digital_ldo_top_VIA1 $T=351090 31760 0 0 $X=350840 $Y=31520
X4417 2 digital_ldo_top_VIA1 $T=351090 37200 0 0 $X=350840 $Y=36960
X4418 2 digital_ldo_top_VIA1 $T=351090 42640 0 0 $X=350840 $Y=42400
X4419 2 digital_ldo_top_VIA1 $T=351090 48080 0 0 $X=350840 $Y=47840
X4420 2 digital_ldo_top_VIA1 $T=351090 53520 0 0 $X=350840 $Y=53280
X4421 2 digital_ldo_top_VIA1 $T=351090 58960 0 0 $X=350840 $Y=58720
X4422 2 digital_ldo_top_VIA1 $T=351090 64400 0 0 $X=350840 $Y=64160
X4423 2 digital_ldo_top_VIA1 $T=351090 69840 0 0 $X=350840 $Y=69600
X4424 2 digital_ldo_top_VIA1 $T=351090 75280 0 0 $X=350840 $Y=75040
X4425 2 digital_ldo_top_VIA1 $T=351090 80720 0 0 $X=350840 $Y=80480
X4426 2 digital_ldo_top_VIA1 $T=351090 86160 0 0 $X=350840 $Y=85920
X4427 2 digital_ldo_top_VIA1 $T=351090 91600 0 0 $X=350840 $Y=91360
X4428 2 digital_ldo_top_VIA1 $T=351090 97040 0 0 $X=350840 $Y=96800
X4429 2 digital_ldo_top_VIA1 $T=351090 102480 0 0 $X=350840 $Y=102240
X4430 2 digital_ldo_top_VIA1 $T=351090 107920 0 0 $X=350840 $Y=107680
X4431 2 digital_ldo_top_VIA1 $T=351090 113360 0 0 $X=350840 $Y=113120
X4432 2 digital_ldo_top_VIA1 $T=351090 118800 0 0 $X=350840 $Y=118560
X4433 2 digital_ldo_top_VIA1 $T=351090 124240 0 0 $X=350840 $Y=124000
X4434 2 digital_ldo_top_VIA1 $T=351090 129680 0 0 $X=350840 $Y=129440
X4435 3 digital_ldo_top_VIA1 $T=353390 12720 0 0 $X=353140 $Y=12480
X4436 3 digital_ldo_top_VIA1 $T=353390 18160 0 0 $X=353140 $Y=17920
X4437 3 digital_ldo_top_VIA1 $T=353390 23600 0 0 $X=353140 $Y=23360
X4438 3 digital_ldo_top_VIA1 $T=353390 29040 0 0 $X=353140 $Y=28800
X4439 3 digital_ldo_top_VIA1 $T=353390 34480 0 0 $X=353140 $Y=34240
X4440 3 digital_ldo_top_VIA1 $T=353390 39920 0 0 $X=353140 $Y=39680
X4441 3 digital_ldo_top_VIA1 $T=353390 45360 0 0 $X=353140 $Y=45120
X4442 3 digital_ldo_top_VIA1 $T=353390 50800 0 0 $X=353140 $Y=50560
X4443 3 digital_ldo_top_VIA1 $T=353390 56240 0 0 $X=353140 $Y=56000
X4444 3 digital_ldo_top_VIA1 $T=353390 61680 0 0 $X=353140 $Y=61440
X4445 3 digital_ldo_top_VIA1 $T=353390 67120 0 0 $X=353140 $Y=66880
X4446 3 digital_ldo_top_VIA1 $T=353390 72560 0 0 $X=353140 $Y=72320
X4447 3 digital_ldo_top_VIA1 $T=353390 78000 0 0 $X=353140 $Y=77760
X4448 3 digital_ldo_top_VIA1 $T=353390 83440 0 0 $X=353140 $Y=83200
X4449 3 digital_ldo_top_VIA1 $T=353390 88880 0 0 $X=353140 $Y=88640
X4450 3 digital_ldo_top_VIA1 $T=353390 94320 0 0 $X=353140 $Y=94080
X4451 3 digital_ldo_top_VIA1 $T=353390 99760 0 0 $X=353140 $Y=99520
X4452 3 digital_ldo_top_VIA1 $T=353390 105200 0 0 $X=353140 $Y=104960
X4453 3 digital_ldo_top_VIA1 $T=353390 110640 0 0 $X=353140 $Y=110400
X4454 3 digital_ldo_top_VIA1 $T=353390 116080 0 0 $X=353140 $Y=115840
X4455 3 digital_ldo_top_VIA1 $T=353390 121520 0 0 $X=353140 $Y=121280
X4456 3 digital_ldo_top_VIA1 $T=353390 126960 0 0 $X=353140 $Y=126720
X4457 2 digital_ldo_top_VIA1 $T=354770 15440 0 0 $X=354520 $Y=15200
X4458 2 digital_ldo_top_VIA1 $T=354770 20880 0 0 $X=354520 $Y=20640
X4459 2 digital_ldo_top_VIA1 $T=354770 26320 0 0 $X=354520 $Y=26080
X4460 2 digital_ldo_top_VIA1 $T=354770 31760 0 0 $X=354520 $Y=31520
X4461 2 digital_ldo_top_VIA1 $T=354770 37200 0 0 $X=354520 $Y=36960
X4462 2 digital_ldo_top_VIA1 $T=354770 42640 0 0 $X=354520 $Y=42400
X4463 2 digital_ldo_top_VIA1 $T=354770 48080 0 0 $X=354520 $Y=47840
X4464 2 digital_ldo_top_VIA1 $T=354770 53520 0 0 $X=354520 $Y=53280
X4465 2 digital_ldo_top_VIA1 $T=354770 58960 0 0 $X=354520 $Y=58720
X4466 2 digital_ldo_top_VIA1 $T=354770 64400 0 0 $X=354520 $Y=64160
X4467 2 digital_ldo_top_VIA1 $T=354770 69840 0 0 $X=354520 $Y=69600
X4468 2 digital_ldo_top_VIA1 $T=354770 75280 0 0 $X=354520 $Y=75040
X4469 2 digital_ldo_top_VIA1 $T=354770 80720 0 0 $X=354520 $Y=80480
X4470 2 digital_ldo_top_VIA1 $T=354770 86160 0 0 $X=354520 $Y=85920
X4471 2 digital_ldo_top_VIA1 $T=354770 91600 0 0 $X=354520 $Y=91360
X4472 2 digital_ldo_top_VIA1 $T=354770 97040 0 0 $X=354520 $Y=96800
X4473 2 digital_ldo_top_VIA1 $T=354770 102480 0 0 $X=354520 $Y=102240
X4474 2 digital_ldo_top_VIA1 $T=354770 107920 0 0 $X=354520 $Y=107680
X4475 2 digital_ldo_top_VIA1 $T=354770 113360 0 0 $X=354520 $Y=113120
X4476 2 digital_ldo_top_VIA1 $T=354770 118800 0 0 $X=354520 $Y=118560
X4477 2 digital_ldo_top_VIA1 $T=354770 124240 0 0 $X=354520 $Y=124000
X4478 2 digital_ldo_top_VIA1 $T=354770 129680 0 0 $X=354520 $Y=129440
X4479 3 digital_ldo_top_VIA1 $T=357070 12720 0 0 $X=356820 $Y=12480
X4480 3 digital_ldo_top_VIA1 $T=357070 18160 0 0 $X=356820 $Y=17920
X4481 3 digital_ldo_top_VIA1 $T=357070 23600 0 0 $X=356820 $Y=23360
X4482 3 digital_ldo_top_VIA1 $T=357070 29040 0 0 $X=356820 $Y=28800
X4483 3 digital_ldo_top_VIA1 $T=357070 34480 0 0 $X=356820 $Y=34240
X4484 3 digital_ldo_top_VIA1 $T=357070 39920 0 0 $X=356820 $Y=39680
X4485 3 digital_ldo_top_VIA1 $T=357070 45360 0 0 $X=356820 $Y=45120
X4486 3 digital_ldo_top_VIA1 $T=357070 50800 0 0 $X=356820 $Y=50560
X4487 3 digital_ldo_top_VIA1 $T=357070 56240 0 0 $X=356820 $Y=56000
X4488 3 digital_ldo_top_VIA1 $T=357070 61680 0 0 $X=356820 $Y=61440
X4489 3 digital_ldo_top_VIA1 $T=357070 67120 0 0 $X=356820 $Y=66880
X4490 3 digital_ldo_top_VIA1 $T=357070 72560 0 0 $X=356820 $Y=72320
X4491 3 digital_ldo_top_VIA1 $T=357070 78000 0 0 $X=356820 $Y=77760
X4492 3 digital_ldo_top_VIA1 $T=357070 83440 0 0 $X=356820 $Y=83200
X4493 3 digital_ldo_top_VIA1 $T=357070 88880 0 0 $X=356820 $Y=88640
X4494 3 digital_ldo_top_VIA1 $T=357070 94320 0 0 $X=356820 $Y=94080
X4495 3 digital_ldo_top_VIA1 $T=357070 99760 0 0 $X=356820 $Y=99520
X4496 3 digital_ldo_top_VIA1 $T=357070 105200 0 0 $X=356820 $Y=104960
X4497 3 digital_ldo_top_VIA1 $T=357070 110640 0 0 $X=356820 $Y=110400
X4498 3 digital_ldo_top_VIA1 $T=357070 116080 0 0 $X=356820 $Y=115840
X4499 3 digital_ldo_top_VIA1 $T=357070 121520 0 0 $X=356820 $Y=121280
X4500 3 digital_ldo_top_VIA1 $T=357070 126960 0 0 $X=356820 $Y=126720
X4501 2 digital_ldo_top_VIA1 $T=358450 15440 0 0 $X=358200 $Y=15200
X4502 2 digital_ldo_top_VIA1 $T=358450 20880 0 0 $X=358200 $Y=20640
X4503 2 digital_ldo_top_VIA1 $T=358450 26320 0 0 $X=358200 $Y=26080
X4504 2 digital_ldo_top_VIA1 $T=358450 31760 0 0 $X=358200 $Y=31520
X4505 2 digital_ldo_top_VIA1 $T=358450 37200 0 0 $X=358200 $Y=36960
X4506 2 digital_ldo_top_VIA1 $T=358450 42640 0 0 $X=358200 $Y=42400
X4507 2 digital_ldo_top_VIA1 $T=358450 48080 0 0 $X=358200 $Y=47840
X4508 2 digital_ldo_top_VIA1 $T=358450 53520 0 0 $X=358200 $Y=53280
X4509 2 digital_ldo_top_VIA1 $T=358450 58960 0 0 $X=358200 $Y=58720
X4510 2 digital_ldo_top_VIA1 $T=358450 64400 0 0 $X=358200 $Y=64160
X4511 2 digital_ldo_top_VIA1 $T=358450 69840 0 0 $X=358200 $Y=69600
X4512 2 digital_ldo_top_VIA1 $T=358450 75280 0 0 $X=358200 $Y=75040
X4513 2 digital_ldo_top_VIA1 $T=358450 80720 0 0 $X=358200 $Y=80480
X4514 2 digital_ldo_top_VIA1 $T=358450 86160 0 0 $X=358200 $Y=85920
X4515 2 digital_ldo_top_VIA1 $T=358450 91600 0 0 $X=358200 $Y=91360
X4516 2 digital_ldo_top_VIA1 $T=358450 97040 0 0 $X=358200 $Y=96800
X4517 2 digital_ldo_top_VIA1 $T=358450 102480 0 0 $X=358200 $Y=102240
X4518 2 digital_ldo_top_VIA1 $T=358450 107920 0 0 $X=358200 $Y=107680
X4519 2 digital_ldo_top_VIA1 $T=358450 113360 0 0 $X=358200 $Y=113120
X4520 2 digital_ldo_top_VIA1 $T=358450 118800 0 0 $X=358200 $Y=118560
X4521 2 digital_ldo_top_VIA1 $T=358450 124240 0 0 $X=358200 $Y=124000
X4522 2 digital_ldo_top_VIA1 $T=358450 129680 0 0 $X=358200 $Y=129440
X4523 3 digital_ldo_top_VIA1 $T=360750 12720 0 0 $X=360500 $Y=12480
X4524 3 digital_ldo_top_VIA1 $T=360750 18160 0 0 $X=360500 $Y=17920
X4525 3 digital_ldo_top_VIA1 $T=360750 23600 0 0 $X=360500 $Y=23360
X4526 3 digital_ldo_top_VIA1 $T=360750 29040 0 0 $X=360500 $Y=28800
X4527 3 digital_ldo_top_VIA1 $T=360750 34480 0 0 $X=360500 $Y=34240
X4528 3 digital_ldo_top_VIA1 $T=360750 39920 0 0 $X=360500 $Y=39680
X4529 3 digital_ldo_top_VIA1 $T=360750 45360 0 0 $X=360500 $Y=45120
X4530 3 digital_ldo_top_VIA1 $T=360750 50800 0 0 $X=360500 $Y=50560
X4531 3 digital_ldo_top_VIA1 $T=360750 56240 0 0 $X=360500 $Y=56000
X4532 3 digital_ldo_top_VIA1 $T=360750 61680 0 0 $X=360500 $Y=61440
X4533 3 digital_ldo_top_VIA1 $T=360750 67120 0 0 $X=360500 $Y=66880
X4534 3 digital_ldo_top_VIA1 $T=360750 72560 0 0 $X=360500 $Y=72320
X4535 3 digital_ldo_top_VIA1 $T=360750 78000 0 0 $X=360500 $Y=77760
X4536 3 digital_ldo_top_VIA1 $T=360750 83440 0 0 $X=360500 $Y=83200
X4537 3 digital_ldo_top_VIA1 $T=360750 88880 0 0 $X=360500 $Y=88640
X4538 3 digital_ldo_top_VIA1 $T=360750 94320 0 0 $X=360500 $Y=94080
X4539 3 digital_ldo_top_VIA1 $T=360750 99760 0 0 $X=360500 $Y=99520
X4540 3 digital_ldo_top_VIA1 $T=360750 105200 0 0 $X=360500 $Y=104960
X4541 3 digital_ldo_top_VIA1 $T=360750 110640 0 0 $X=360500 $Y=110400
X4542 3 digital_ldo_top_VIA1 $T=360750 116080 0 0 $X=360500 $Y=115840
X4543 3 digital_ldo_top_VIA1 $T=360750 121520 0 0 $X=360500 $Y=121280
X4544 3 digital_ldo_top_VIA1 $T=360750 126960 0 0 $X=360500 $Y=126720
X4545 2 digital_ldo_top_VIA1 $T=362130 15440 0 0 $X=361880 $Y=15200
X4546 2 digital_ldo_top_VIA1 $T=362130 20880 0 0 $X=361880 $Y=20640
X4547 2 digital_ldo_top_VIA1 $T=362130 26320 0 0 $X=361880 $Y=26080
X4548 2 digital_ldo_top_VIA1 $T=362130 31760 0 0 $X=361880 $Y=31520
X4549 2 digital_ldo_top_VIA1 $T=362130 37200 0 0 $X=361880 $Y=36960
X4550 2 digital_ldo_top_VIA1 $T=362130 42640 0 0 $X=361880 $Y=42400
X4551 2 digital_ldo_top_VIA1 $T=362130 48080 0 0 $X=361880 $Y=47840
X4552 2 digital_ldo_top_VIA1 $T=362130 53520 0 0 $X=361880 $Y=53280
X4553 2 digital_ldo_top_VIA1 $T=362130 58960 0 0 $X=361880 $Y=58720
X4554 2 digital_ldo_top_VIA1 $T=362130 64400 0 0 $X=361880 $Y=64160
X4555 2 digital_ldo_top_VIA1 $T=362130 69840 0 0 $X=361880 $Y=69600
X4556 2 digital_ldo_top_VIA1 $T=362130 75280 0 0 $X=361880 $Y=75040
X4557 2 digital_ldo_top_VIA1 $T=362130 80720 0 0 $X=361880 $Y=80480
X4558 2 digital_ldo_top_VIA1 $T=362130 86160 0 0 $X=361880 $Y=85920
X4559 2 digital_ldo_top_VIA1 $T=362130 91600 0 0 $X=361880 $Y=91360
X4560 2 digital_ldo_top_VIA1 $T=362130 97040 0 0 $X=361880 $Y=96800
X4561 2 digital_ldo_top_VIA1 $T=362130 102480 0 0 $X=361880 $Y=102240
X4562 2 digital_ldo_top_VIA1 $T=362130 107920 0 0 $X=361880 $Y=107680
X4563 2 digital_ldo_top_VIA1 $T=362130 113360 0 0 $X=361880 $Y=113120
X4564 2 digital_ldo_top_VIA1 $T=362130 118800 0 0 $X=361880 $Y=118560
X4565 2 digital_ldo_top_VIA1 $T=362130 124240 0 0 $X=361880 $Y=124000
X4566 2 digital_ldo_top_VIA1 $T=362130 129680 0 0 $X=361880 $Y=129440
X4567 3 digital_ldo_top_VIA1 $T=364430 12720 0 0 $X=364180 $Y=12480
X4568 3 digital_ldo_top_VIA1 $T=364430 18160 0 0 $X=364180 $Y=17920
X4569 3 digital_ldo_top_VIA1 $T=364430 23600 0 0 $X=364180 $Y=23360
X4570 3 digital_ldo_top_VIA1 $T=364430 29040 0 0 $X=364180 $Y=28800
X4571 3 digital_ldo_top_VIA1 $T=364430 34480 0 0 $X=364180 $Y=34240
X4572 3 digital_ldo_top_VIA1 $T=364430 39920 0 0 $X=364180 $Y=39680
X4573 3 digital_ldo_top_VIA1 $T=364430 45360 0 0 $X=364180 $Y=45120
X4574 3 digital_ldo_top_VIA1 $T=364430 50800 0 0 $X=364180 $Y=50560
X4575 3 digital_ldo_top_VIA1 $T=364430 56240 0 0 $X=364180 $Y=56000
X4576 3 digital_ldo_top_VIA1 $T=364430 61680 0 0 $X=364180 $Y=61440
X4577 3 digital_ldo_top_VIA1 $T=364430 67120 0 0 $X=364180 $Y=66880
X4578 3 digital_ldo_top_VIA1 $T=364430 72560 0 0 $X=364180 $Y=72320
X4579 3 digital_ldo_top_VIA1 $T=364430 78000 0 0 $X=364180 $Y=77760
X4580 3 digital_ldo_top_VIA1 $T=364430 83440 0 0 $X=364180 $Y=83200
X4581 3 digital_ldo_top_VIA1 $T=364430 88880 0 0 $X=364180 $Y=88640
X4582 3 digital_ldo_top_VIA1 $T=364430 94320 0 0 $X=364180 $Y=94080
X4583 3 digital_ldo_top_VIA1 $T=364430 99760 0 0 $X=364180 $Y=99520
X4584 3 digital_ldo_top_VIA1 $T=364430 105200 0 0 $X=364180 $Y=104960
X4585 3 digital_ldo_top_VIA1 $T=364430 110640 0 0 $X=364180 $Y=110400
X4586 3 digital_ldo_top_VIA1 $T=364430 116080 0 0 $X=364180 $Y=115840
X4587 3 digital_ldo_top_VIA1 $T=364430 121520 0 0 $X=364180 $Y=121280
X4588 3 digital_ldo_top_VIA1 $T=364430 126960 0 0 $X=364180 $Y=126720
X4589 2 digital_ldo_top_VIA1 $T=365810 15440 0 0 $X=365560 $Y=15200
X4590 2 digital_ldo_top_VIA1 $T=365810 20880 0 0 $X=365560 $Y=20640
X4591 2 digital_ldo_top_VIA1 $T=365810 26320 0 0 $X=365560 $Y=26080
X4592 2 digital_ldo_top_VIA1 $T=365810 31760 0 0 $X=365560 $Y=31520
X4593 2 digital_ldo_top_VIA1 $T=365810 37200 0 0 $X=365560 $Y=36960
X4594 2 digital_ldo_top_VIA1 $T=365810 42640 0 0 $X=365560 $Y=42400
X4595 2 digital_ldo_top_VIA1 $T=365810 48080 0 0 $X=365560 $Y=47840
X4596 2 digital_ldo_top_VIA1 $T=365810 53520 0 0 $X=365560 $Y=53280
X4597 2 digital_ldo_top_VIA1 $T=365810 58960 0 0 $X=365560 $Y=58720
X4598 2 digital_ldo_top_VIA1 $T=365810 64400 0 0 $X=365560 $Y=64160
X4599 2 digital_ldo_top_VIA1 $T=365810 69840 0 0 $X=365560 $Y=69600
X4600 2 digital_ldo_top_VIA1 $T=365810 75280 0 0 $X=365560 $Y=75040
X4601 2 digital_ldo_top_VIA1 $T=365810 80720 0 0 $X=365560 $Y=80480
X4602 2 digital_ldo_top_VIA1 $T=365810 86160 0 0 $X=365560 $Y=85920
X4603 2 digital_ldo_top_VIA1 $T=365810 91600 0 0 $X=365560 $Y=91360
X4604 2 digital_ldo_top_VIA1 $T=365810 97040 0 0 $X=365560 $Y=96800
X4605 2 digital_ldo_top_VIA1 $T=365810 102480 0 0 $X=365560 $Y=102240
X4606 2 digital_ldo_top_VIA1 $T=365810 107920 0 0 $X=365560 $Y=107680
X4607 2 digital_ldo_top_VIA1 $T=365810 113360 0 0 $X=365560 $Y=113120
X4608 2 digital_ldo_top_VIA1 $T=365810 118800 0 0 $X=365560 $Y=118560
X4609 2 digital_ldo_top_VIA1 $T=365810 124240 0 0 $X=365560 $Y=124000
X4610 2 digital_ldo_top_VIA1 $T=365810 129680 0 0 $X=365560 $Y=129440
X4611 3 digital_ldo_top_VIA1 $T=368110 12720 0 0 $X=367860 $Y=12480
X4612 3 digital_ldo_top_VIA1 $T=368110 18160 0 0 $X=367860 $Y=17920
X4613 3 digital_ldo_top_VIA1 $T=368110 23600 0 0 $X=367860 $Y=23360
X4614 3 digital_ldo_top_VIA1 $T=368110 29040 0 0 $X=367860 $Y=28800
X4615 3 digital_ldo_top_VIA1 $T=368110 34480 0 0 $X=367860 $Y=34240
X4616 3 digital_ldo_top_VIA1 $T=368110 39920 0 0 $X=367860 $Y=39680
X4617 3 digital_ldo_top_VIA1 $T=368110 45360 0 0 $X=367860 $Y=45120
X4618 3 digital_ldo_top_VIA1 $T=368110 50800 0 0 $X=367860 $Y=50560
X4619 3 digital_ldo_top_VIA1 $T=368110 56240 0 0 $X=367860 $Y=56000
X4620 3 digital_ldo_top_VIA1 $T=368110 61680 0 0 $X=367860 $Y=61440
X4621 3 digital_ldo_top_VIA1 $T=368110 67120 0 0 $X=367860 $Y=66880
X4622 3 digital_ldo_top_VIA1 $T=368110 72560 0 0 $X=367860 $Y=72320
X4623 3 digital_ldo_top_VIA1 $T=368110 78000 0 0 $X=367860 $Y=77760
X4624 3 digital_ldo_top_VIA1 $T=368110 83440 0 0 $X=367860 $Y=83200
X4625 3 digital_ldo_top_VIA1 $T=368110 88880 0 0 $X=367860 $Y=88640
X4626 3 digital_ldo_top_VIA1 $T=368110 94320 0 0 $X=367860 $Y=94080
X4627 3 digital_ldo_top_VIA1 $T=368110 99760 0 0 $X=367860 $Y=99520
X4628 3 digital_ldo_top_VIA1 $T=368110 105200 0 0 $X=367860 $Y=104960
X4629 3 digital_ldo_top_VIA1 $T=368110 110640 0 0 $X=367860 $Y=110400
X4630 3 digital_ldo_top_VIA1 $T=368110 116080 0 0 $X=367860 $Y=115840
X4631 3 digital_ldo_top_VIA1 $T=368110 121520 0 0 $X=367860 $Y=121280
X4632 3 digital_ldo_top_VIA1 $T=368110 126960 0 0 $X=367860 $Y=126720
X4633 2 digital_ldo_top_VIA1 $T=369490 15440 0 0 $X=369240 $Y=15200
X4634 2 digital_ldo_top_VIA1 $T=369490 20880 0 0 $X=369240 $Y=20640
X4635 2 digital_ldo_top_VIA1 $T=369490 26320 0 0 $X=369240 $Y=26080
X4636 2 digital_ldo_top_VIA1 $T=369490 31760 0 0 $X=369240 $Y=31520
X4637 2 digital_ldo_top_VIA1 $T=369490 37200 0 0 $X=369240 $Y=36960
X4638 2 digital_ldo_top_VIA1 $T=369490 42640 0 0 $X=369240 $Y=42400
X4639 2 digital_ldo_top_VIA1 $T=369490 48080 0 0 $X=369240 $Y=47840
X4640 2 digital_ldo_top_VIA1 $T=369490 53520 0 0 $X=369240 $Y=53280
X4641 2 digital_ldo_top_VIA1 $T=369490 58960 0 0 $X=369240 $Y=58720
X4642 2 digital_ldo_top_VIA1 $T=369490 64400 0 0 $X=369240 $Y=64160
X4643 2 digital_ldo_top_VIA1 $T=369490 69840 0 0 $X=369240 $Y=69600
X4644 2 digital_ldo_top_VIA1 $T=369490 75280 0 0 $X=369240 $Y=75040
X4645 2 digital_ldo_top_VIA1 $T=369490 80720 0 0 $X=369240 $Y=80480
X4646 2 digital_ldo_top_VIA1 $T=369490 86160 0 0 $X=369240 $Y=85920
X4647 2 digital_ldo_top_VIA1 $T=369490 91600 0 0 $X=369240 $Y=91360
X4648 2 digital_ldo_top_VIA1 $T=369490 97040 0 0 $X=369240 $Y=96800
X4649 2 digital_ldo_top_VIA1 $T=369490 102480 0 0 $X=369240 $Y=102240
X4650 2 digital_ldo_top_VIA1 $T=369490 107920 0 0 $X=369240 $Y=107680
X4651 2 digital_ldo_top_VIA1 $T=369490 113360 0 0 $X=369240 $Y=113120
X4652 2 digital_ldo_top_VIA1 $T=369490 118800 0 0 $X=369240 $Y=118560
X4653 2 digital_ldo_top_VIA1 $T=369490 124240 0 0 $X=369240 $Y=124000
X4654 2 digital_ldo_top_VIA1 $T=369490 129680 0 0 $X=369240 $Y=129440
X4655 3 digital_ldo_top_VIA1 $T=371790 12720 0 0 $X=371540 $Y=12480
X4656 3 digital_ldo_top_VIA1 $T=371790 18160 0 0 $X=371540 $Y=17920
X4657 3 digital_ldo_top_VIA1 $T=371790 23600 0 0 $X=371540 $Y=23360
X4658 3 digital_ldo_top_VIA1 $T=371790 29040 0 0 $X=371540 $Y=28800
X4659 3 digital_ldo_top_VIA1 $T=371790 34480 0 0 $X=371540 $Y=34240
X4660 3 digital_ldo_top_VIA1 $T=371790 39920 0 0 $X=371540 $Y=39680
X4661 3 digital_ldo_top_VIA1 $T=371790 45360 0 0 $X=371540 $Y=45120
X4662 3 digital_ldo_top_VIA1 $T=371790 50800 0 0 $X=371540 $Y=50560
X4663 3 digital_ldo_top_VIA1 $T=371790 56240 0 0 $X=371540 $Y=56000
X4664 3 digital_ldo_top_VIA1 $T=371790 61680 0 0 $X=371540 $Y=61440
X4665 3 digital_ldo_top_VIA1 $T=371790 67120 0 0 $X=371540 $Y=66880
X4666 3 digital_ldo_top_VIA1 $T=371790 72560 0 0 $X=371540 $Y=72320
X4667 3 digital_ldo_top_VIA1 $T=371790 78000 0 0 $X=371540 $Y=77760
X4668 3 digital_ldo_top_VIA1 $T=371790 83440 0 0 $X=371540 $Y=83200
X4669 3 digital_ldo_top_VIA1 $T=371790 88880 0 0 $X=371540 $Y=88640
X4670 3 digital_ldo_top_VIA1 $T=371790 94320 0 0 $X=371540 $Y=94080
X4671 3 digital_ldo_top_VIA1 $T=371790 99760 0 0 $X=371540 $Y=99520
X4672 3 digital_ldo_top_VIA1 $T=371790 105200 0 0 $X=371540 $Y=104960
X4673 3 digital_ldo_top_VIA1 $T=371790 110640 0 0 $X=371540 $Y=110400
X4674 3 digital_ldo_top_VIA1 $T=371790 116080 0 0 $X=371540 $Y=115840
X4675 3 digital_ldo_top_VIA1 $T=371790 121520 0 0 $X=371540 $Y=121280
X4676 3 digital_ldo_top_VIA1 $T=371790 126960 0 0 $X=371540 $Y=126720
X4677 2 digital_ldo_top_VIA1 $T=373170 15440 0 0 $X=372920 $Y=15200
X4678 2 digital_ldo_top_VIA1 $T=373170 20880 0 0 $X=372920 $Y=20640
X4679 2 digital_ldo_top_VIA1 $T=373170 26320 0 0 $X=372920 $Y=26080
X4680 2 digital_ldo_top_VIA1 $T=373170 31760 0 0 $X=372920 $Y=31520
X4681 2 digital_ldo_top_VIA1 $T=373170 37200 0 0 $X=372920 $Y=36960
X4682 2 digital_ldo_top_VIA1 $T=373170 42640 0 0 $X=372920 $Y=42400
X4683 2 digital_ldo_top_VIA1 $T=373170 48080 0 0 $X=372920 $Y=47840
X4684 2 digital_ldo_top_VIA1 $T=373170 53520 0 0 $X=372920 $Y=53280
X4685 2 digital_ldo_top_VIA1 $T=373170 58960 0 0 $X=372920 $Y=58720
X4686 2 digital_ldo_top_VIA1 $T=373170 64400 0 0 $X=372920 $Y=64160
X4687 2 digital_ldo_top_VIA1 $T=373170 69840 0 0 $X=372920 $Y=69600
X4688 2 digital_ldo_top_VIA1 $T=373170 75280 0 0 $X=372920 $Y=75040
X4689 2 digital_ldo_top_VIA1 $T=373170 80720 0 0 $X=372920 $Y=80480
X4690 2 digital_ldo_top_VIA1 $T=373170 86160 0 0 $X=372920 $Y=85920
X4691 2 digital_ldo_top_VIA1 $T=373170 91600 0 0 $X=372920 $Y=91360
X4692 2 digital_ldo_top_VIA1 $T=373170 97040 0 0 $X=372920 $Y=96800
X4693 2 digital_ldo_top_VIA1 $T=373170 102480 0 0 $X=372920 $Y=102240
X4694 2 digital_ldo_top_VIA1 $T=373170 107920 0 0 $X=372920 $Y=107680
X4695 2 digital_ldo_top_VIA1 $T=373170 113360 0 0 $X=372920 $Y=113120
X4696 2 digital_ldo_top_VIA1 $T=373170 118800 0 0 $X=372920 $Y=118560
X4697 2 digital_ldo_top_VIA1 $T=373170 124240 0 0 $X=372920 $Y=124000
X4698 2 digital_ldo_top_VIA1 $T=373170 129680 0 0 $X=372920 $Y=129440
X4699 3 digital_ldo_top_VIA1 $T=375470 12720 0 0 $X=375220 $Y=12480
X4700 3 digital_ldo_top_VIA1 $T=375470 18160 0 0 $X=375220 $Y=17920
X4701 3 digital_ldo_top_VIA1 $T=375470 23600 0 0 $X=375220 $Y=23360
X4702 3 digital_ldo_top_VIA1 $T=375470 29040 0 0 $X=375220 $Y=28800
X4703 3 digital_ldo_top_VIA1 $T=375470 34480 0 0 $X=375220 $Y=34240
X4704 3 digital_ldo_top_VIA1 $T=375470 39920 0 0 $X=375220 $Y=39680
X4705 3 digital_ldo_top_VIA1 $T=375470 45360 0 0 $X=375220 $Y=45120
X4706 3 digital_ldo_top_VIA1 $T=375470 50800 0 0 $X=375220 $Y=50560
X4707 3 digital_ldo_top_VIA1 $T=375470 56240 0 0 $X=375220 $Y=56000
X4708 3 digital_ldo_top_VIA1 $T=375470 61680 0 0 $X=375220 $Y=61440
X4709 3 digital_ldo_top_VIA1 $T=375470 67120 0 0 $X=375220 $Y=66880
X4710 3 digital_ldo_top_VIA1 $T=375470 72560 0 0 $X=375220 $Y=72320
X4711 3 digital_ldo_top_VIA1 $T=375470 78000 0 0 $X=375220 $Y=77760
X4712 3 digital_ldo_top_VIA1 $T=375470 83440 0 0 $X=375220 $Y=83200
X4713 3 digital_ldo_top_VIA1 $T=375470 88880 0 0 $X=375220 $Y=88640
X4714 3 digital_ldo_top_VIA1 $T=375470 94320 0 0 $X=375220 $Y=94080
X4715 3 digital_ldo_top_VIA1 $T=375470 99760 0 0 $X=375220 $Y=99520
X4716 3 digital_ldo_top_VIA1 $T=375470 105200 0 0 $X=375220 $Y=104960
X4717 3 digital_ldo_top_VIA1 $T=375470 110640 0 0 $X=375220 $Y=110400
X4718 3 digital_ldo_top_VIA1 $T=375470 116080 0 0 $X=375220 $Y=115840
X4719 3 digital_ldo_top_VIA1 $T=375470 121520 0 0 $X=375220 $Y=121280
X4720 3 digital_ldo_top_VIA1 $T=375470 126960 0 0 $X=375220 $Y=126720
X4721 2 digital_ldo_top_VIA1 $T=376850 15440 0 0 $X=376600 $Y=15200
X4722 2 digital_ldo_top_VIA1 $T=376850 20880 0 0 $X=376600 $Y=20640
X4723 2 digital_ldo_top_VIA1 $T=376850 26320 0 0 $X=376600 $Y=26080
X4724 2 digital_ldo_top_VIA1 $T=376850 31760 0 0 $X=376600 $Y=31520
X4725 2 digital_ldo_top_VIA1 $T=376850 37200 0 0 $X=376600 $Y=36960
X4726 2 digital_ldo_top_VIA1 $T=376850 42640 0 0 $X=376600 $Y=42400
X4727 2 digital_ldo_top_VIA1 $T=376850 48080 0 0 $X=376600 $Y=47840
X4728 2 digital_ldo_top_VIA1 $T=376850 53520 0 0 $X=376600 $Y=53280
X4729 2 digital_ldo_top_VIA1 $T=376850 58960 0 0 $X=376600 $Y=58720
X4730 2 digital_ldo_top_VIA1 $T=376850 64400 0 0 $X=376600 $Y=64160
X4731 2 digital_ldo_top_VIA1 $T=376850 69840 0 0 $X=376600 $Y=69600
X4732 2 digital_ldo_top_VIA1 $T=376850 75280 0 0 $X=376600 $Y=75040
X4733 2 digital_ldo_top_VIA1 $T=376850 80720 0 0 $X=376600 $Y=80480
X4734 2 digital_ldo_top_VIA1 $T=376850 86160 0 0 $X=376600 $Y=85920
X4735 2 digital_ldo_top_VIA1 $T=376850 91600 0 0 $X=376600 $Y=91360
X4736 2 digital_ldo_top_VIA1 $T=376850 97040 0 0 $X=376600 $Y=96800
X4737 2 digital_ldo_top_VIA1 $T=376850 102480 0 0 $X=376600 $Y=102240
X4738 2 digital_ldo_top_VIA1 $T=376850 107920 0 0 $X=376600 $Y=107680
X4739 2 digital_ldo_top_VIA1 $T=376850 113360 0 0 $X=376600 $Y=113120
X4740 2 digital_ldo_top_VIA1 $T=376850 118800 0 0 $X=376600 $Y=118560
X4741 2 digital_ldo_top_VIA1 $T=376850 124240 0 0 $X=376600 $Y=124000
X4742 2 digital_ldo_top_VIA1 $T=376850 129680 0 0 $X=376600 $Y=129440
X4743 3 digital_ldo_top_VIA1 $T=379150 12720 0 0 $X=378900 $Y=12480
X4744 3 digital_ldo_top_VIA1 $T=379150 18160 0 0 $X=378900 $Y=17920
X4745 3 digital_ldo_top_VIA1 $T=379150 23600 0 0 $X=378900 $Y=23360
X4746 3 digital_ldo_top_VIA1 $T=379150 29040 0 0 $X=378900 $Y=28800
X4747 3 digital_ldo_top_VIA1 $T=379150 34480 0 0 $X=378900 $Y=34240
X4748 3 digital_ldo_top_VIA1 $T=379150 39920 0 0 $X=378900 $Y=39680
X4749 3 digital_ldo_top_VIA1 $T=379150 45360 0 0 $X=378900 $Y=45120
X4750 3 digital_ldo_top_VIA1 $T=379150 50800 0 0 $X=378900 $Y=50560
X4751 3 digital_ldo_top_VIA1 $T=379150 56240 0 0 $X=378900 $Y=56000
X4752 3 digital_ldo_top_VIA1 $T=379150 61680 0 0 $X=378900 $Y=61440
X4753 3 digital_ldo_top_VIA1 $T=379150 67120 0 0 $X=378900 $Y=66880
X4754 3 digital_ldo_top_VIA1 $T=379150 72560 0 0 $X=378900 $Y=72320
X4755 3 digital_ldo_top_VIA1 $T=379150 78000 0 0 $X=378900 $Y=77760
X4756 3 digital_ldo_top_VIA1 $T=379150 83440 0 0 $X=378900 $Y=83200
X4757 3 digital_ldo_top_VIA1 $T=379150 88880 0 0 $X=378900 $Y=88640
X4758 3 digital_ldo_top_VIA1 $T=379150 94320 0 0 $X=378900 $Y=94080
X4759 3 digital_ldo_top_VIA1 $T=379150 99760 0 0 $X=378900 $Y=99520
X4760 3 digital_ldo_top_VIA1 $T=379150 105200 0 0 $X=378900 $Y=104960
X4761 3 digital_ldo_top_VIA1 $T=379150 110640 0 0 $X=378900 $Y=110400
X4762 3 digital_ldo_top_VIA1 $T=379150 116080 0 0 $X=378900 $Y=115840
X4763 3 digital_ldo_top_VIA1 $T=379150 121520 0 0 $X=378900 $Y=121280
X4764 3 digital_ldo_top_VIA1 $T=379150 126960 0 0 $X=378900 $Y=126720
X4765 3 digital_ldo_top_VIA2 $T=40590 27710 0 0 $X=40340 $Y=27510
X4766 3 digital_ldo_top_VIA2 $T=40590 31490 0 0 $X=40340 $Y=31290
X4767 3 digital_ldo_top_VIA2 $T=40590 37970 0 0 $X=40340 $Y=37770
X4768 2 digital_ldo_top_VIA2 $T=41970 48230 0 0 $X=41720 $Y=48030
X4769 2 digital_ldo_top_VIA2 $T=41970 51470 0 0 $X=41720 $Y=51270
X4770 3 digital_ldo_top_VIA2 $T=44270 27710 0 0 $X=44020 $Y=27510
X4771 3 digital_ldo_top_VIA2 $T=47950 27710 0 0 $X=47700 $Y=27510
X4772 2 digital_ldo_top_VIA2 $T=49330 48230 0 0 $X=49080 $Y=48030
X4773 2 digital_ldo_top_VIA2 $T=49330 51470 0 0 $X=49080 $Y=51270
X4774 2 digital_ldo_top_VIA2 $T=49330 54170 0 0 $X=49080 $Y=53970
X4775 2 digital_ldo_top_VIA3 $T=53230 15440 0 0 $X=53100 $Y=15200
X4776 2 digital_ldo_top_VIA3 $T=53230 20880 0 0 $X=53100 $Y=20640
X4777 2 digital_ldo_top_VIA3 $T=53230 26320 0 0 $X=53100 $Y=26080
X4778 2 digital_ldo_top_VIA3 $T=53230 31760 0 0 $X=53100 $Y=31520
X4779 2 digital_ldo_top_VIA3 $T=53230 37200 0 0 $X=53100 $Y=36960
X4780 2 digital_ldo_top_VIA3 $T=53230 42640 0 0 $X=53100 $Y=42400
X4781 2 digital_ldo_top_VIA3 $T=53230 48080 0 0 $X=53100 $Y=47840
X4782 2 digital_ldo_top_VIA3 $T=53230 53520 0 0 $X=53100 $Y=53280
X4783 2 digital_ldo_top_VIA3 $T=53230 58960 0 0 $X=53100 $Y=58720
X4784 3 digital_ldo_top_VIA4 $T=11150 11700 0 0 $X=10900 $Y=11470
X4785 3 digital_ldo_top_VIA4 $T=11150 15780 0 0 $X=10900 $Y=15550
X4786 3 digital_ldo_top_VIA4 $T=11150 19860 0 0 $X=10900 $Y=19630
X4787 3 digital_ldo_top_VIA4 $T=11150 23940 0 0 $X=10900 $Y=23710
X4788 3 digital_ldo_top_VIA4 $T=11150 28020 0 0 $X=10900 $Y=27790
X4789 3 digital_ldo_top_VIA4 $T=11150 32100 0 0 $X=10900 $Y=31870
X4790 3 digital_ldo_top_VIA4 $T=11150 36180 0 0 $X=10900 $Y=35950
X4791 3 digital_ldo_top_VIA4 $T=11150 40260 0 0 $X=10900 $Y=40030
X4792 3 digital_ldo_top_VIA4 $T=11150 44340 0 0 $X=10900 $Y=44110
X4793 3 digital_ldo_top_VIA4 $T=11150 48420 0 0 $X=10900 $Y=48190
X4794 3 digital_ldo_top_VIA4 $T=11150 52500 0 0 $X=10900 $Y=52270
X4795 3 digital_ldo_top_VIA4 $T=11150 56580 0 0 $X=10900 $Y=56350
X4796 3 digital_ldo_top_VIA4 $T=11150 60660 0 0 $X=10900 $Y=60430
X4797 3 digital_ldo_top_VIA4 $T=11150 64740 0 0 $X=10900 $Y=64510
X4798 3 digital_ldo_top_VIA4 $T=11150 68820 0 0 $X=10900 $Y=68590
X4799 3 digital_ldo_top_VIA4 $T=11150 72900 0 0 $X=10900 $Y=72670
X4800 3 digital_ldo_top_VIA4 $T=11150 76980 0 0 $X=10900 $Y=76750
X4801 3 digital_ldo_top_VIA4 $T=11150 81060 0 0 $X=10900 $Y=80830
X4802 3 digital_ldo_top_VIA4 $T=11150 85140 0 0 $X=10900 $Y=84910
X4803 3 digital_ldo_top_VIA4 $T=11150 89220 0 0 $X=10900 $Y=88990
X4804 3 digital_ldo_top_VIA4 $T=11150 93300 0 0 $X=10900 $Y=93070
X4805 3 digital_ldo_top_VIA4 $T=11150 97380 0 0 $X=10900 $Y=97150
X4806 3 digital_ldo_top_VIA4 $T=11150 101460 0 0 $X=10900 $Y=101230
X4807 3 digital_ldo_top_VIA4 $T=11150 105540 0 0 $X=10900 $Y=105310
X4808 3 digital_ldo_top_VIA4 $T=11150 109620 0 0 $X=10900 $Y=109390
X4809 3 digital_ldo_top_VIA4 $T=11150 113700 0 0 $X=10900 $Y=113470
X4810 3 digital_ldo_top_VIA4 $T=11150 117780 0 0 $X=10900 $Y=117550
X4811 3 digital_ldo_top_VIA4 $T=11150 121860 0 0 $X=10900 $Y=121630
X4812 3 digital_ldo_top_VIA4 $T=11150 125940 0 0 $X=10900 $Y=125710
X4813 2 digital_ldo_top_VIA4 $T=12530 13060 0 0 $X=12280 $Y=12830
X4814 2 digital_ldo_top_VIA4 $T=12530 17140 0 0 $X=12280 $Y=16910
X4815 2 digital_ldo_top_VIA4 $T=12530 21220 0 0 $X=12280 $Y=20990
X4816 2 digital_ldo_top_VIA4 $T=12530 25300 0 0 $X=12280 $Y=25070
X4817 2 digital_ldo_top_VIA4 $T=12530 29380 0 0 $X=12280 $Y=29150
X4818 2 digital_ldo_top_VIA4 $T=12530 33460 0 0 $X=12280 $Y=33230
X4819 2 digital_ldo_top_VIA4 $T=12530 37540 0 0 $X=12280 $Y=37310
X4820 2 digital_ldo_top_VIA4 $T=12530 41620 0 0 $X=12280 $Y=41390
X4821 2 digital_ldo_top_VIA4 $T=12530 45700 0 0 $X=12280 $Y=45470
X4822 2 digital_ldo_top_VIA4 $T=12530 49780 0 0 $X=12280 $Y=49550
X4823 2 digital_ldo_top_VIA4 $T=12530 53860 0 0 $X=12280 $Y=53630
X4824 2 digital_ldo_top_VIA4 $T=12530 57940 0 0 $X=12280 $Y=57710
X4825 2 digital_ldo_top_VIA4 $T=12530 62020 0 0 $X=12280 $Y=61790
X4826 2 digital_ldo_top_VIA4 $T=12530 66100 0 0 $X=12280 $Y=65870
X4827 2 digital_ldo_top_VIA4 $T=12530 70180 0 0 $X=12280 $Y=69950
X4828 2 digital_ldo_top_VIA4 $T=12530 74260 0 0 $X=12280 $Y=74030
X4829 2 digital_ldo_top_VIA4 $T=12530 78340 0 0 $X=12280 $Y=78110
X4830 2 digital_ldo_top_VIA4 $T=12530 82420 0 0 $X=12280 $Y=82190
X4831 2 digital_ldo_top_VIA4 $T=12530 86500 0 0 $X=12280 $Y=86270
X4832 2 digital_ldo_top_VIA4 $T=12530 90580 0 0 $X=12280 $Y=90350
X4833 2 digital_ldo_top_VIA4 $T=12530 94660 0 0 $X=12280 $Y=94430
X4834 2 digital_ldo_top_VIA4 $T=12530 98740 0 0 $X=12280 $Y=98510
X4835 2 digital_ldo_top_VIA4 $T=12530 102820 0 0 $X=12280 $Y=102590
X4836 2 digital_ldo_top_VIA4 $T=12530 106900 0 0 $X=12280 $Y=106670
X4837 2 digital_ldo_top_VIA4 $T=12530 110980 0 0 $X=12280 $Y=110750
X4838 2 digital_ldo_top_VIA4 $T=12530 115060 0 0 $X=12280 $Y=114830
X4839 2 digital_ldo_top_VIA4 $T=12530 119140 0 0 $X=12280 $Y=118910
X4840 2 digital_ldo_top_VIA4 $T=12530 123220 0 0 $X=12280 $Y=122990
X4841 2 digital_ldo_top_VIA4 $T=12530 127300 0 0 $X=12280 $Y=127070
X4842 3 digital_ldo_top_VIA4 $T=14830 11700 0 0 $X=14580 $Y=11470
X4843 3 digital_ldo_top_VIA4 $T=14830 15780 0 0 $X=14580 $Y=15550
X4844 3 digital_ldo_top_VIA4 $T=14830 19860 0 0 $X=14580 $Y=19630
X4845 3 digital_ldo_top_VIA4 $T=14830 23940 0 0 $X=14580 $Y=23710
X4846 3 digital_ldo_top_VIA4 $T=14830 28020 0 0 $X=14580 $Y=27790
X4847 3 digital_ldo_top_VIA4 $T=14830 32100 0 0 $X=14580 $Y=31870
X4848 3 digital_ldo_top_VIA4 $T=14830 36180 0 0 $X=14580 $Y=35950
X4849 3 digital_ldo_top_VIA4 $T=14830 40260 0 0 $X=14580 $Y=40030
X4850 3 digital_ldo_top_VIA4 $T=14830 44340 0 0 $X=14580 $Y=44110
X4851 3 digital_ldo_top_VIA4 $T=14830 48420 0 0 $X=14580 $Y=48190
X4852 3 digital_ldo_top_VIA4 $T=14830 52500 0 0 $X=14580 $Y=52270
X4853 3 digital_ldo_top_VIA4 $T=14830 56580 0 0 $X=14580 $Y=56350
X4854 3 digital_ldo_top_VIA4 $T=14830 60660 0 0 $X=14580 $Y=60430
X4855 3 digital_ldo_top_VIA4 $T=14830 64740 0 0 $X=14580 $Y=64510
X4856 3 digital_ldo_top_VIA4 $T=14830 68820 0 0 $X=14580 $Y=68590
X4857 3 digital_ldo_top_VIA4 $T=14830 72900 0 0 $X=14580 $Y=72670
X4858 3 digital_ldo_top_VIA4 $T=14830 76980 0 0 $X=14580 $Y=76750
X4859 3 digital_ldo_top_VIA4 $T=14830 81060 0 0 $X=14580 $Y=80830
X4860 3 digital_ldo_top_VIA4 $T=14830 85140 0 0 $X=14580 $Y=84910
X4861 3 digital_ldo_top_VIA4 $T=14830 89220 0 0 $X=14580 $Y=88990
X4862 3 digital_ldo_top_VIA4 $T=14830 93300 0 0 $X=14580 $Y=93070
X4863 3 digital_ldo_top_VIA4 $T=14830 97380 0 0 $X=14580 $Y=97150
X4864 3 digital_ldo_top_VIA4 $T=14830 101460 0 0 $X=14580 $Y=101230
X4865 3 digital_ldo_top_VIA4 $T=14830 105540 0 0 $X=14580 $Y=105310
X4866 3 digital_ldo_top_VIA4 $T=14830 109620 0 0 $X=14580 $Y=109390
X4867 3 digital_ldo_top_VIA4 $T=14830 113700 0 0 $X=14580 $Y=113470
X4868 3 digital_ldo_top_VIA4 $T=14830 117780 0 0 $X=14580 $Y=117550
X4869 3 digital_ldo_top_VIA4 $T=14830 121860 0 0 $X=14580 $Y=121630
X4870 3 digital_ldo_top_VIA4 $T=14830 125940 0 0 $X=14580 $Y=125710
X4871 2 digital_ldo_top_VIA4 $T=16210 13060 0 0 $X=15960 $Y=12830
X4872 2 digital_ldo_top_VIA4 $T=16210 17140 0 0 $X=15960 $Y=16910
X4873 2 digital_ldo_top_VIA4 $T=16210 21220 0 0 $X=15960 $Y=20990
X4874 2 digital_ldo_top_VIA4 $T=16210 25300 0 0 $X=15960 $Y=25070
X4875 2 digital_ldo_top_VIA4 $T=16210 29380 0 0 $X=15960 $Y=29150
X4876 2 digital_ldo_top_VIA4 $T=16210 33460 0 0 $X=15960 $Y=33230
X4877 2 digital_ldo_top_VIA4 $T=16210 37540 0 0 $X=15960 $Y=37310
X4878 2 digital_ldo_top_VIA4 $T=16210 41620 0 0 $X=15960 $Y=41390
X4879 2 digital_ldo_top_VIA4 $T=16210 45700 0 0 $X=15960 $Y=45470
X4880 2 digital_ldo_top_VIA4 $T=16210 49780 0 0 $X=15960 $Y=49550
X4881 2 digital_ldo_top_VIA4 $T=16210 53860 0 0 $X=15960 $Y=53630
X4882 2 digital_ldo_top_VIA4 $T=16210 57940 0 0 $X=15960 $Y=57710
X4883 2 digital_ldo_top_VIA4 $T=16210 62020 0 0 $X=15960 $Y=61790
X4884 2 digital_ldo_top_VIA4 $T=16210 66100 0 0 $X=15960 $Y=65870
X4885 2 digital_ldo_top_VIA4 $T=16210 70180 0 0 $X=15960 $Y=69950
X4886 2 digital_ldo_top_VIA4 $T=16210 74260 0 0 $X=15960 $Y=74030
X4887 2 digital_ldo_top_VIA4 $T=16210 78340 0 0 $X=15960 $Y=78110
X4888 2 digital_ldo_top_VIA4 $T=16210 82420 0 0 $X=15960 $Y=82190
X4889 2 digital_ldo_top_VIA4 $T=16210 86500 0 0 $X=15960 $Y=86270
X4890 2 digital_ldo_top_VIA4 $T=16210 90580 0 0 $X=15960 $Y=90350
X4891 2 digital_ldo_top_VIA4 $T=16210 94660 0 0 $X=15960 $Y=94430
X4892 2 digital_ldo_top_VIA4 $T=16210 98740 0 0 $X=15960 $Y=98510
X4893 2 digital_ldo_top_VIA4 $T=16210 102820 0 0 $X=15960 $Y=102590
X4894 2 digital_ldo_top_VIA4 $T=16210 106900 0 0 $X=15960 $Y=106670
X4895 2 digital_ldo_top_VIA4 $T=16210 110980 0 0 $X=15960 $Y=110750
X4896 2 digital_ldo_top_VIA4 $T=16210 115060 0 0 $X=15960 $Y=114830
X4897 2 digital_ldo_top_VIA4 $T=16210 119140 0 0 $X=15960 $Y=118910
X4898 2 digital_ldo_top_VIA4 $T=16210 123220 0 0 $X=15960 $Y=122990
X4899 2 digital_ldo_top_VIA4 $T=16210 127300 0 0 $X=15960 $Y=127070
X4900 3 digital_ldo_top_VIA4 $T=18510 11700 0 0 $X=18260 $Y=11470
X4901 3 digital_ldo_top_VIA4 $T=18510 36180 0 0 $X=18260 $Y=35950
X4902 3 digital_ldo_top_VIA4 $T=18510 40260 0 0 $X=18260 $Y=40030
X4903 3 digital_ldo_top_VIA4 $T=18510 44340 0 0 $X=18260 $Y=44110
X4904 3 digital_ldo_top_VIA4 $T=18510 48420 0 0 $X=18260 $Y=48190
X4905 3 digital_ldo_top_VIA4 $T=18510 52500 0 0 $X=18260 $Y=52270
X4906 3 digital_ldo_top_VIA4 $T=18510 56580 0 0 $X=18260 $Y=56350
X4907 3 digital_ldo_top_VIA4 $T=18510 60660 0 0 $X=18260 $Y=60430
X4908 3 digital_ldo_top_VIA4 $T=18510 64740 0 0 $X=18260 $Y=64510
X4909 3 digital_ldo_top_VIA4 $T=18510 68820 0 0 $X=18260 $Y=68590
X4910 3 digital_ldo_top_VIA4 $T=18510 72900 0 0 $X=18260 $Y=72670
X4911 3 digital_ldo_top_VIA4 $T=18510 76980 0 0 $X=18260 $Y=76750
X4912 3 digital_ldo_top_VIA4 $T=18510 81060 0 0 $X=18260 $Y=80830
X4913 3 digital_ldo_top_VIA4 $T=18510 85140 0 0 $X=18260 $Y=84910
X4914 3 digital_ldo_top_VIA4 $T=18510 89220 0 0 $X=18260 $Y=88990
X4915 3 digital_ldo_top_VIA4 $T=18510 93300 0 0 $X=18260 $Y=93070
X4916 3 digital_ldo_top_VIA4 $T=18510 97380 0 0 $X=18260 $Y=97150
X4917 3 digital_ldo_top_VIA4 $T=18510 101460 0 0 $X=18260 $Y=101230
X4918 3 digital_ldo_top_VIA4 $T=18510 105540 0 0 $X=18260 $Y=105310
X4919 3 digital_ldo_top_VIA4 $T=18510 109620 0 0 $X=18260 $Y=109390
X4920 3 digital_ldo_top_VIA4 $T=18510 113700 0 0 $X=18260 $Y=113470
X4921 3 digital_ldo_top_VIA4 $T=18510 117780 0 0 $X=18260 $Y=117550
X4922 3 digital_ldo_top_VIA4 $T=18510 121860 0 0 $X=18260 $Y=121630
X4923 3 digital_ldo_top_VIA4 $T=18510 125940 0 0 $X=18260 $Y=125710
X4924 2 digital_ldo_top_VIA4 $T=19890 13060 0 0 $X=19640 $Y=12830
X4925 2 digital_ldo_top_VIA4 $T=19890 33460 0 0 $X=19640 $Y=33230
X4926 2 digital_ldo_top_VIA4 $T=19890 37540 0 0 $X=19640 $Y=37310
X4927 2 digital_ldo_top_VIA4 $T=19890 41620 0 0 $X=19640 $Y=41390
X4928 2 digital_ldo_top_VIA4 $T=19890 45700 0 0 $X=19640 $Y=45470
X4929 2 digital_ldo_top_VIA4 $T=19890 49780 0 0 $X=19640 $Y=49550
X4930 2 digital_ldo_top_VIA4 $T=19890 53860 0 0 $X=19640 $Y=53630
X4931 2 digital_ldo_top_VIA4 $T=19890 57940 0 0 $X=19640 $Y=57710
X4932 2 digital_ldo_top_VIA4 $T=19890 62020 0 0 $X=19640 $Y=61790
X4933 2 digital_ldo_top_VIA4 $T=19890 66100 0 0 $X=19640 $Y=65870
X4934 2 digital_ldo_top_VIA4 $T=19890 70180 0 0 $X=19640 $Y=69950
X4935 2 digital_ldo_top_VIA4 $T=19890 74260 0 0 $X=19640 $Y=74030
X4936 2 digital_ldo_top_VIA4 $T=19890 78340 0 0 $X=19640 $Y=78110
X4937 2 digital_ldo_top_VIA4 $T=19890 82420 0 0 $X=19640 $Y=82190
X4938 2 digital_ldo_top_VIA4 $T=19890 86500 0 0 $X=19640 $Y=86270
X4939 2 digital_ldo_top_VIA4 $T=19890 90580 0 0 $X=19640 $Y=90350
X4940 2 digital_ldo_top_VIA4 $T=19890 94660 0 0 $X=19640 $Y=94430
X4941 2 digital_ldo_top_VIA4 $T=19890 98740 0 0 $X=19640 $Y=98510
X4942 2 digital_ldo_top_VIA4 $T=19890 102820 0 0 $X=19640 $Y=102590
X4943 2 digital_ldo_top_VIA4 $T=19890 106900 0 0 $X=19640 $Y=106670
X4944 2 digital_ldo_top_VIA4 $T=19890 110980 0 0 $X=19640 $Y=110750
X4945 2 digital_ldo_top_VIA4 $T=19890 115060 0 0 $X=19640 $Y=114830
X4946 2 digital_ldo_top_VIA4 $T=19890 119140 0 0 $X=19640 $Y=118910
X4947 2 digital_ldo_top_VIA4 $T=19890 123220 0 0 $X=19640 $Y=122990
X4948 2 digital_ldo_top_VIA4 $T=19890 127300 0 0 $X=19640 $Y=127070
X4949 3 digital_ldo_top_VIA4 $T=22190 11700 0 0 $X=21940 $Y=11470
X4950 3 digital_ldo_top_VIA4 $T=22190 36180 0 0 $X=21940 $Y=35950
X4951 3 digital_ldo_top_VIA4 $T=22190 40260 0 0 $X=21940 $Y=40030
X4952 3 digital_ldo_top_VIA4 $T=22190 44340 0 0 $X=21940 $Y=44110
X4953 3 digital_ldo_top_VIA4 $T=22190 48420 0 0 $X=21940 $Y=48190
X4954 3 digital_ldo_top_VIA4 $T=22190 52500 0 0 $X=21940 $Y=52270
X4955 3 digital_ldo_top_VIA4 $T=22190 56580 0 0 $X=21940 $Y=56350
X4956 3 digital_ldo_top_VIA4 $T=22190 60660 0 0 $X=21940 $Y=60430
X4957 3 digital_ldo_top_VIA4 $T=22190 64740 0 0 $X=21940 $Y=64510
X4958 3 digital_ldo_top_VIA4 $T=22190 68820 0 0 $X=21940 $Y=68590
X4959 3 digital_ldo_top_VIA4 $T=22190 72900 0 0 $X=21940 $Y=72670
X4960 3 digital_ldo_top_VIA4 $T=22190 76980 0 0 $X=21940 $Y=76750
X4961 3 digital_ldo_top_VIA4 $T=22190 81060 0 0 $X=21940 $Y=80830
X4962 3 digital_ldo_top_VIA4 $T=22190 85140 0 0 $X=21940 $Y=84910
X4963 3 digital_ldo_top_VIA4 $T=22190 89220 0 0 $X=21940 $Y=88990
X4964 3 digital_ldo_top_VIA4 $T=22190 93300 0 0 $X=21940 $Y=93070
X4965 3 digital_ldo_top_VIA4 $T=22190 97380 0 0 $X=21940 $Y=97150
X4966 3 digital_ldo_top_VIA4 $T=22190 101460 0 0 $X=21940 $Y=101230
X4967 3 digital_ldo_top_VIA4 $T=22190 105540 0 0 $X=21940 $Y=105310
X4968 3 digital_ldo_top_VIA4 $T=22190 109620 0 0 $X=21940 $Y=109390
X4969 3 digital_ldo_top_VIA4 $T=22190 113700 0 0 $X=21940 $Y=113470
X4970 3 digital_ldo_top_VIA4 $T=22190 117780 0 0 $X=21940 $Y=117550
X4971 3 digital_ldo_top_VIA4 $T=22190 121860 0 0 $X=21940 $Y=121630
X4972 3 digital_ldo_top_VIA4 $T=22190 125940 0 0 $X=21940 $Y=125710
X4973 2 digital_ldo_top_VIA4 $T=23570 13060 0 0 $X=23320 $Y=12830
X4974 2 digital_ldo_top_VIA4 $T=23570 33460 0 0 $X=23320 $Y=33230
X4975 2 digital_ldo_top_VIA4 $T=23570 37540 0 0 $X=23320 $Y=37310
X4976 2 digital_ldo_top_VIA4 $T=23570 41620 0 0 $X=23320 $Y=41390
X4977 2 digital_ldo_top_VIA4 $T=23570 45700 0 0 $X=23320 $Y=45470
X4978 2 digital_ldo_top_VIA4 $T=23570 49780 0 0 $X=23320 $Y=49550
X4979 2 digital_ldo_top_VIA4 $T=23570 53860 0 0 $X=23320 $Y=53630
X4980 2 digital_ldo_top_VIA4 $T=23570 57940 0 0 $X=23320 $Y=57710
X4981 2 digital_ldo_top_VIA4 $T=23570 62020 0 0 $X=23320 $Y=61790
X4982 2 digital_ldo_top_VIA4 $T=23570 66100 0 0 $X=23320 $Y=65870
X4983 2 digital_ldo_top_VIA4 $T=23570 70180 0 0 $X=23320 $Y=69950
X4984 2 digital_ldo_top_VIA4 $T=23570 74260 0 0 $X=23320 $Y=74030
X4985 2 digital_ldo_top_VIA4 $T=23570 78340 0 0 $X=23320 $Y=78110
X4986 2 digital_ldo_top_VIA4 $T=23570 82420 0 0 $X=23320 $Y=82190
X4987 2 digital_ldo_top_VIA4 $T=23570 86500 0 0 $X=23320 $Y=86270
X4988 2 digital_ldo_top_VIA4 $T=23570 90580 0 0 $X=23320 $Y=90350
X4989 2 digital_ldo_top_VIA4 $T=23570 94660 0 0 $X=23320 $Y=94430
X4990 2 digital_ldo_top_VIA4 $T=23570 98740 0 0 $X=23320 $Y=98510
X4991 2 digital_ldo_top_VIA4 $T=23570 102820 0 0 $X=23320 $Y=102590
X4992 2 digital_ldo_top_VIA4 $T=23570 106900 0 0 $X=23320 $Y=106670
X4993 2 digital_ldo_top_VIA4 $T=23570 110980 0 0 $X=23320 $Y=110750
X4994 2 digital_ldo_top_VIA4 $T=23570 115060 0 0 $X=23320 $Y=114830
X4995 2 digital_ldo_top_VIA4 $T=23570 119140 0 0 $X=23320 $Y=118910
X4996 2 digital_ldo_top_VIA4 $T=23570 123220 0 0 $X=23320 $Y=122990
X4997 2 digital_ldo_top_VIA4 $T=23570 127300 0 0 $X=23320 $Y=127070
X4998 3 digital_ldo_top_VIA4 $T=25870 11700 0 0 $X=25620 $Y=11470
X4999 3 digital_ldo_top_VIA4 $T=25870 36180 0 0 $X=25620 $Y=35950
X5000 3 digital_ldo_top_VIA4 $T=25870 40260 0 0 $X=25620 $Y=40030
X5001 3 digital_ldo_top_VIA4 $T=25870 44340 0 0 $X=25620 $Y=44110
X5002 3 digital_ldo_top_VIA4 $T=25870 48420 0 0 $X=25620 $Y=48190
X5003 3 digital_ldo_top_VIA4 $T=25870 52500 0 0 $X=25620 $Y=52270
X5004 3 digital_ldo_top_VIA4 $T=25870 56580 0 0 $X=25620 $Y=56350
X5005 3 digital_ldo_top_VIA4 $T=25870 60660 0 0 $X=25620 $Y=60430
X5006 3 digital_ldo_top_VIA4 $T=25870 64740 0 0 $X=25620 $Y=64510
X5007 3 digital_ldo_top_VIA4 $T=25870 68820 0 0 $X=25620 $Y=68590
X5008 3 digital_ldo_top_VIA4 $T=25870 72900 0 0 $X=25620 $Y=72670
X5009 3 digital_ldo_top_VIA4 $T=25870 76980 0 0 $X=25620 $Y=76750
X5010 3 digital_ldo_top_VIA4 $T=25870 81060 0 0 $X=25620 $Y=80830
X5011 3 digital_ldo_top_VIA4 $T=25870 85140 0 0 $X=25620 $Y=84910
X5012 3 digital_ldo_top_VIA4 $T=25870 89220 0 0 $X=25620 $Y=88990
X5013 3 digital_ldo_top_VIA4 $T=25870 93300 0 0 $X=25620 $Y=93070
X5014 3 digital_ldo_top_VIA4 $T=25870 97380 0 0 $X=25620 $Y=97150
X5015 3 digital_ldo_top_VIA4 $T=25870 101460 0 0 $X=25620 $Y=101230
X5016 3 digital_ldo_top_VIA4 $T=25870 105540 0 0 $X=25620 $Y=105310
X5017 3 digital_ldo_top_VIA4 $T=25870 109620 0 0 $X=25620 $Y=109390
X5018 3 digital_ldo_top_VIA4 $T=25870 113700 0 0 $X=25620 $Y=113470
X5019 3 digital_ldo_top_VIA4 $T=25870 117780 0 0 $X=25620 $Y=117550
X5020 3 digital_ldo_top_VIA4 $T=25870 121860 0 0 $X=25620 $Y=121630
X5021 3 digital_ldo_top_VIA4 $T=25870 125940 0 0 $X=25620 $Y=125710
X5022 2 digital_ldo_top_VIA4 $T=27250 13060 0 0 $X=27000 $Y=12830
X5023 2 digital_ldo_top_VIA4 $T=27250 33460 0 0 $X=27000 $Y=33230
X5024 2 digital_ldo_top_VIA4 $T=27250 37540 0 0 $X=27000 $Y=37310
X5025 2 digital_ldo_top_VIA4 $T=27250 41620 0 0 $X=27000 $Y=41390
X5026 2 digital_ldo_top_VIA4 $T=27250 45700 0 0 $X=27000 $Y=45470
X5027 2 digital_ldo_top_VIA4 $T=27250 49780 0 0 $X=27000 $Y=49550
X5028 2 digital_ldo_top_VIA4 $T=27250 53860 0 0 $X=27000 $Y=53630
X5029 2 digital_ldo_top_VIA4 $T=27250 57940 0 0 $X=27000 $Y=57710
X5030 2 digital_ldo_top_VIA4 $T=27250 62020 0 0 $X=27000 $Y=61790
X5031 2 digital_ldo_top_VIA4 $T=27250 66100 0 0 $X=27000 $Y=65870
X5032 2 digital_ldo_top_VIA4 $T=27250 70180 0 0 $X=27000 $Y=69950
X5033 2 digital_ldo_top_VIA4 $T=27250 74260 0 0 $X=27000 $Y=74030
X5034 2 digital_ldo_top_VIA4 $T=27250 78340 0 0 $X=27000 $Y=78110
X5035 2 digital_ldo_top_VIA4 $T=27250 82420 0 0 $X=27000 $Y=82190
X5036 2 digital_ldo_top_VIA4 $T=27250 86500 0 0 $X=27000 $Y=86270
X5037 2 digital_ldo_top_VIA4 $T=27250 90580 0 0 $X=27000 $Y=90350
X5038 2 digital_ldo_top_VIA4 $T=27250 94660 0 0 $X=27000 $Y=94430
X5039 2 digital_ldo_top_VIA4 $T=27250 98740 0 0 $X=27000 $Y=98510
X5040 2 digital_ldo_top_VIA4 $T=27250 102820 0 0 $X=27000 $Y=102590
X5041 2 digital_ldo_top_VIA4 $T=27250 106900 0 0 $X=27000 $Y=106670
X5042 2 digital_ldo_top_VIA4 $T=27250 110980 0 0 $X=27000 $Y=110750
X5043 2 digital_ldo_top_VIA4 $T=27250 115060 0 0 $X=27000 $Y=114830
X5044 2 digital_ldo_top_VIA4 $T=27250 119140 0 0 $X=27000 $Y=118910
X5045 2 digital_ldo_top_VIA4 $T=27250 123220 0 0 $X=27000 $Y=122990
X5046 2 digital_ldo_top_VIA4 $T=27250 127300 0 0 $X=27000 $Y=127070
X5047 3 digital_ldo_top_VIA4 $T=29550 11700 0 0 $X=29300 $Y=11470
X5048 3 digital_ldo_top_VIA4 $T=29550 36180 0 0 $X=29300 $Y=35950
X5049 3 digital_ldo_top_VIA4 $T=29550 40260 0 0 $X=29300 $Y=40030
X5050 3 digital_ldo_top_VIA4 $T=29550 44340 0 0 $X=29300 $Y=44110
X5051 3 digital_ldo_top_VIA4 $T=29550 48420 0 0 $X=29300 $Y=48190
X5052 3 digital_ldo_top_VIA4 $T=29550 52500 0 0 $X=29300 $Y=52270
X5053 3 digital_ldo_top_VIA4 $T=29550 56580 0 0 $X=29300 $Y=56350
X5054 3 digital_ldo_top_VIA4 $T=29550 60660 0 0 $X=29300 $Y=60430
X5055 3 digital_ldo_top_VIA4 $T=29550 64740 0 0 $X=29300 $Y=64510
X5056 3 digital_ldo_top_VIA4 $T=29550 68820 0 0 $X=29300 $Y=68590
X5057 3 digital_ldo_top_VIA4 $T=29550 72900 0 0 $X=29300 $Y=72670
X5058 3 digital_ldo_top_VIA4 $T=29550 76980 0 0 $X=29300 $Y=76750
X5059 3 digital_ldo_top_VIA4 $T=29550 81060 0 0 $X=29300 $Y=80830
X5060 3 digital_ldo_top_VIA4 $T=29550 85140 0 0 $X=29300 $Y=84910
X5061 3 digital_ldo_top_VIA4 $T=29550 89220 0 0 $X=29300 $Y=88990
X5062 3 digital_ldo_top_VIA4 $T=29550 93300 0 0 $X=29300 $Y=93070
X5063 3 digital_ldo_top_VIA4 $T=29550 97380 0 0 $X=29300 $Y=97150
X5064 3 digital_ldo_top_VIA4 $T=29550 101460 0 0 $X=29300 $Y=101230
X5065 3 digital_ldo_top_VIA4 $T=29550 105540 0 0 $X=29300 $Y=105310
X5066 3 digital_ldo_top_VIA4 $T=29550 109620 0 0 $X=29300 $Y=109390
X5067 3 digital_ldo_top_VIA4 $T=29550 113700 0 0 $X=29300 $Y=113470
X5068 3 digital_ldo_top_VIA4 $T=29550 117780 0 0 $X=29300 $Y=117550
X5069 3 digital_ldo_top_VIA4 $T=29550 121860 0 0 $X=29300 $Y=121630
X5070 3 digital_ldo_top_VIA4 $T=29550 125940 0 0 $X=29300 $Y=125710
X5071 2 digital_ldo_top_VIA4 $T=30930 13060 0 0 $X=30680 $Y=12830
X5072 2 digital_ldo_top_VIA4 $T=30930 17140 0 0 $X=30680 $Y=16910
X5073 2 digital_ldo_top_VIA4 $T=30930 21220 0 0 $X=30680 $Y=20990
X5074 2 digital_ldo_top_VIA4 $T=30930 25300 0 0 $X=30680 $Y=25070
X5075 2 digital_ldo_top_VIA4 $T=30930 29380 0 0 $X=30680 $Y=29150
X5076 2 digital_ldo_top_VIA4 $T=30930 33460 0 0 $X=30680 $Y=33230
X5077 2 digital_ldo_top_VIA4 $T=30930 37540 0 0 $X=30680 $Y=37310
X5078 2 digital_ldo_top_VIA4 $T=30930 41620 0 0 $X=30680 $Y=41390
X5079 2 digital_ldo_top_VIA4 $T=30930 45700 0 0 $X=30680 $Y=45470
X5080 2 digital_ldo_top_VIA4 $T=30930 49780 0 0 $X=30680 $Y=49550
X5081 2 digital_ldo_top_VIA4 $T=30930 53860 0 0 $X=30680 $Y=53630
X5082 2 digital_ldo_top_VIA4 $T=30930 57940 0 0 $X=30680 $Y=57710
X5083 2 digital_ldo_top_VIA4 $T=30930 62020 0 0 $X=30680 $Y=61790
X5084 2 digital_ldo_top_VIA4 $T=30930 66100 0 0 $X=30680 $Y=65870
X5085 2 digital_ldo_top_VIA4 $T=30930 70180 0 0 $X=30680 $Y=69950
X5086 2 digital_ldo_top_VIA4 $T=30930 74260 0 0 $X=30680 $Y=74030
X5087 2 digital_ldo_top_VIA4 $T=30930 78340 0 0 $X=30680 $Y=78110
X5088 2 digital_ldo_top_VIA4 $T=30930 82420 0 0 $X=30680 $Y=82190
X5089 2 digital_ldo_top_VIA4 $T=30930 86500 0 0 $X=30680 $Y=86270
X5090 2 digital_ldo_top_VIA4 $T=30930 90580 0 0 $X=30680 $Y=90350
X5091 2 digital_ldo_top_VIA4 $T=30930 94660 0 0 $X=30680 $Y=94430
X5092 2 digital_ldo_top_VIA4 $T=30930 98740 0 0 $X=30680 $Y=98510
X5093 2 digital_ldo_top_VIA4 $T=30930 102820 0 0 $X=30680 $Y=102590
X5094 2 digital_ldo_top_VIA4 $T=30930 106900 0 0 $X=30680 $Y=106670
X5095 2 digital_ldo_top_VIA4 $T=30930 110980 0 0 $X=30680 $Y=110750
X5096 2 digital_ldo_top_VIA4 $T=30930 115060 0 0 $X=30680 $Y=114830
X5097 2 digital_ldo_top_VIA4 $T=30930 119140 0 0 $X=30680 $Y=118910
X5098 2 digital_ldo_top_VIA4 $T=30930 123220 0 0 $X=30680 $Y=122990
X5099 2 digital_ldo_top_VIA4 $T=30930 127300 0 0 $X=30680 $Y=127070
X5100 3 digital_ldo_top_VIA4 $T=33230 11700 0 0 $X=32980 $Y=11470
X5101 3 digital_ldo_top_VIA4 $T=33230 15780 0 0 $X=32980 $Y=15550
X5102 3 digital_ldo_top_VIA4 $T=33230 19860 0 0 $X=32980 $Y=19630
X5103 3 digital_ldo_top_VIA4 $T=33230 23940 0 0 $X=32980 $Y=23710
X5104 3 digital_ldo_top_VIA4 $T=33230 28020 0 0 $X=32980 $Y=27790
X5105 3 digital_ldo_top_VIA4 $T=33230 32100 0 0 $X=32980 $Y=31870
X5106 3 digital_ldo_top_VIA4 $T=33230 36180 0 0 $X=32980 $Y=35950
X5107 3 digital_ldo_top_VIA4 $T=33230 40260 0 0 $X=32980 $Y=40030
X5108 3 digital_ldo_top_VIA4 $T=33230 44340 0 0 $X=32980 $Y=44110
X5109 3 digital_ldo_top_VIA4 $T=33230 48420 0 0 $X=32980 $Y=48190
X5110 3 digital_ldo_top_VIA4 $T=33230 52500 0 0 $X=32980 $Y=52270
X5111 3 digital_ldo_top_VIA4 $T=33230 56580 0 0 $X=32980 $Y=56350
X5112 3 digital_ldo_top_VIA4 $T=33230 60660 0 0 $X=32980 $Y=60430
X5113 3 digital_ldo_top_VIA4 $T=33230 64740 0 0 $X=32980 $Y=64510
X5114 3 digital_ldo_top_VIA4 $T=33230 68820 0 0 $X=32980 $Y=68590
X5115 3 digital_ldo_top_VIA4 $T=33230 72900 0 0 $X=32980 $Y=72670
X5116 3 digital_ldo_top_VIA4 $T=33230 76980 0 0 $X=32980 $Y=76750
X5117 3 digital_ldo_top_VIA4 $T=33230 81060 0 0 $X=32980 $Y=80830
X5118 3 digital_ldo_top_VIA4 $T=33230 85140 0 0 $X=32980 $Y=84910
X5119 3 digital_ldo_top_VIA4 $T=33230 89220 0 0 $X=32980 $Y=88990
X5120 3 digital_ldo_top_VIA4 $T=33230 93300 0 0 $X=32980 $Y=93070
X5121 3 digital_ldo_top_VIA4 $T=33230 97380 0 0 $X=32980 $Y=97150
X5122 3 digital_ldo_top_VIA4 $T=33230 101460 0 0 $X=32980 $Y=101230
X5123 3 digital_ldo_top_VIA4 $T=33230 105540 0 0 $X=32980 $Y=105310
X5124 3 digital_ldo_top_VIA4 $T=33230 109620 0 0 $X=32980 $Y=109390
X5125 3 digital_ldo_top_VIA4 $T=33230 113700 0 0 $X=32980 $Y=113470
X5126 3 digital_ldo_top_VIA4 $T=33230 117780 0 0 $X=32980 $Y=117550
X5127 3 digital_ldo_top_VIA4 $T=33230 121860 0 0 $X=32980 $Y=121630
X5128 3 digital_ldo_top_VIA4 $T=33230 125940 0 0 $X=32980 $Y=125710
X5129 2 digital_ldo_top_VIA4 $T=34610 13060 0 0 $X=34360 $Y=12830
X5130 2 digital_ldo_top_VIA4 $T=34610 17140 0 0 $X=34360 $Y=16910
X5131 2 digital_ldo_top_VIA4 $T=34610 21220 0 0 $X=34360 $Y=20990
X5132 2 digital_ldo_top_VIA4 $T=34610 25300 0 0 $X=34360 $Y=25070
X5133 2 digital_ldo_top_VIA4 $T=34610 29380 0 0 $X=34360 $Y=29150
X5134 2 digital_ldo_top_VIA4 $T=34610 33460 0 0 $X=34360 $Y=33230
X5135 2 digital_ldo_top_VIA4 $T=34610 37540 0 0 $X=34360 $Y=37310
X5136 2 digital_ldo_top_VIA4 $T=34610 41620 0 0 $X=34360 $Y=41390
X5137 2 digital_ldo_top_VIA4 $T=34610 45700 0 0 $X=34360 $Y=45470
X5138 2 digital_ldo_top_VIA4 $T=34610 49780 0 0 $X=34360 $Y=49550
X5139 2 digital_ldo_top_VIA4 $T=34610 53860 0 0 $X=34360 $Y=53630
X5140 2 digital_ldo_top_VIA4 $T=34610 57940 0 0 $X=34360 $Y=57710
X5141 2 digital_ldo_top_VIA4 $T=34610 62020 0 0 $X=34360 $Y=61790
X5142 2 digital_ldo_top_VIA4 $T=34610 66100 0 0 $X=34360 $Y=65870
X5143 2 digital_ldo_top_VIA4 $T=34610 70180 0 0 $X=34360 $Y=69950
X5144 2 digital_ldo_top_VIA4 $T=34610 74260 0 0 $X=34360 $Y=74030
X5145 2 digital_ldo_top_VIA4 $T=34610 78340 0 0 $X=34360 $Y=78110
X5146 2 digital_ldo_top_VIA4 $T=34610 82420 0 0 $X=34360 $Y=82190
X5147 2 digital_ldo_top_VIA4 $T=34610 86500 0 0 $X=34360 $Y=86270
X5148 2 digital_ldo_top_VIA4 $T=34610 90580 0 0 $X=34360 $Y=90350
X5149 2 digital_ldo_top_VIA4 $T=34610 94660 0 0 $X=34360 $Y=94430
X5150 2 digital_ldo_top_VIA4 $T=34610 98740 0 0 $X=34360 $Y=98510
X5151 2 digital_ldo_top_VIA4 $T=34610 102820 0 0 $X=34360 $Y=102590
X5152 2 digital_ldo_top_VIA4 $T=34610 106900 0 0 $X=34360 $Y=106670
X5153 2 digital_ldo_top_VIA4 $T=34610 110980 0 0 $X=34360 $Y=110750
X5154 2 digital_ldo_top_VIA4 $T=34610 115060 0 0 $X=34360 $Y=114830
X5155 2 digital_ldo_top_VIA4 $T=34610 119140 0 0 $X=34360 $Y=118910
X5156 2 digital_ldo_top_VIA4 $T=34610 123220 0 0 $X=34360 $Y=122990
X5157 2 digital_ldo_top_VIA4 $T=34610 127300 0 0 $X=34360 $Y=127070
X5158 3 digital_ldo_top_VIA4 $T=36910 11700 0 0 $X=36660 $Y=11470
X5159 3 digital_ldo_top_VIA4 $T=36910 15780 0 0 $X=36660 $Y=15550
X5160 3 digital_ldo_top_VIA4 $T=36910 19860 0 0 $X=36660 $Y=19630
X5161 3 digital_ldo_top_VIA4 $T=36910 23940 0 0 $X=36660 $Y=23710
X5162 3 digital_ldo_top_VIA4 $T=36910 28020 0 0 $X=36660 $Y=27790
X5163 3 digital_ldo_top_VIA4 $T=36910 32100 0 0 $X=36660 $Y=31870
X5164 3 digital_ldo_top_VIA4 $T=36910 36180 0 0 $X=36660 $Y=35950
X5165 3 digital_ldo_top_VIA4 $T=36910 40260 0 0 $X=36660 $Y=40030
X5166 3 digital_ldo_top_VIA4 $T=36910 44340 0 0 $X=36660 $Y=44110
X5167 3 digital_ldo_top_VIA4 $T=36910 48420 0 0 $X=36660 $Y=48190
X5168 3 digital_ldo_top_VIA4 $T=36910 52500 0 0 $X=36660 $Y=52270
X5169 3 digital_ldo_top_VIA4 $T=36910 56580 0 0 $X=36660 $Y=56350
X5170 3 digital_ldo_top_VIA4 $T=36910 60660 0 0 $X=36660 $Y=60430
X5171 3 digital_ldo_top_VIA4 $T=36910 64740 0 0 $X=36660 $Y=64510
X5172 3 digital_ldo_top_VIA4 $T=36910 68820 0 0 $X=36660 $Y=68590
X5173 3 digital_ldo_top_VIA4 $T=36910 72900 0 0 $X=36660 $Y=72670
X5174 3 digital_ldo_top_VIA4 $T=36910 76980 0 0 $X=36660 $Y=76750
X5175 3 digital_ldo_top_VIA4 $T=36910 81060 0 0 $X=36660 $Y=80830
X5176 3 digital_ldo_top_VIA4 $T=36910 85140 0 0 $X=36660 $Y=84910
X5177 3 digital_ldo_top_VIA4 $T=36910 89220 0 0 $X=36660 $Y=88990
X5178 3 digital_ldo_top_VIA4 $T=36910 93300 0 0 $X=36660 $Y=93070
X5179 3 digital_ldo_top_VIA4 $T=36910 97380 0 0 $X=36660 $Y=97150
X5180 3 digital_ldo_top_VIA4 $T=36910 101460 0 0 $X=36660 $Y=101230
X5181 3 digital_ldo_top_VIA4 $T=36910 105540 0 0 $X=36660 $Y=105310
X5182 3 digital_ldo_top_VIA4 $T=36910 109620 0 0 $X=36660 $Y=109390
X5183 3 digital_ldo_top_VIA4 $T=36910 113700 0 0 $X=36660 $Y=113470
X5184 3 digital_ldo_top_VIA4 $T=36910 117780 0 0 $X=36660 $Y=117550
X5185 3 digital_ldo_top_VIA4 $T=36910 121860 0 0 $X=36660 $Y=121630
X5186 3 digital_ldo_top_VIA4 $T=36910 125940 0 0 $X=36660 $Y=125710
X5187 2 digital_ldo_top_VIA4 $T=38290 13060 0 0 $X=38040 $Y=12830
X5188 2 digital_ldo_top_VIA4 $T=38290 17140 0 0 $X=38040 $Y=16910
X5189 2 digital_ldo_top_VIA4 $T=38290 21220 0 0 $X=38040 $Y=20990
X5190 2 digital_ldo_top_VIA4 $T=38290 25300 0 0 $X=38040 $Y=25070
X5191 2 digital_ldo_top_VIA4 $T=38290 29380 0 0 $X=38040 $Y=29150
X5192 2 digital_ldo_top_VIA4 $T=38290 33460 0 0 $X=38040 $Y=33230
X5193 2 digital_ldo_top_VIA4 $T=38290 37540 0 0 $X=38040 $Y=37310
X5194 2 digital_ldo_top_VIA4 $T=38290 41620 0 0 $X=38040 $Y=41390
X5195 2 digital_ldo_top_VIA4 $T=38290 45700 0 0 $X=38040 $Y=45470
X5196 2 digital_ldo_top_VIA4 $T=38290 49780 0 0 $X=38040 $Y=49550
X5197 2 digital_ldo_top_VIA4 $T=38290 53860 0 0 $X=38040 $Y=53630
X5198 2 digital_ldo_top_VIA4 $T=38290 57940 0 0 $X=38040 $Y=57710
X5199 2 digital_ldo_top_VIA4 $T=38290 62020 0 0 $X=38040 $Y=61790
X5200 2 digital_ldo_top_VIA4 $T=38290 66100 0 0 $X=38040 $Y=65870
X5201 2 digital_ldo_top_VIA4 $T=38290 70180 0 0 $X=38040 $Y=69950
X5202 2 digital_ldo_top_VIA4 $T=38290 74260 0 0 $X=38040 $Y=74030
X5203 2 digital_ldo_top_VIA4 $T=38290 78340 0 0 $X=38040 $Y=78110
X5204 2 digital_ldo_top_VIA4 $T=38290 82420 0 0 $X=38040 $Y=82190
X5205 2 digital_ldo_top_VIA4 $T=38290 86500 0 0 $X=38040 $Y=86270
X5206 2 digital_ldo_top_VIA4 $T=38290 90580 0 0 $X=38040 $Y=90350
X5207 2 digital_ldo_top_VIA4 $T=38290 94660 0 0 $X=38040 $Y=94430
X5208 2 digital_ldo_top_VIA4 $T=38290 98740 0 0 $X=38040 $Y=98510
X5209 2 digital_ldo_top_VIA4 $T=38290 102820 0 0 $X=38040 $Y=102590
X5210 2 digital_ldo_top_VIA4 $T=38290 106900 0 0 $X=38040 $Y=106670
X5211 2 digital_ldo_top_VIA4 $T=38290 110980 0 0 $X=38040 $Y=110750
X5212 2 digital_ldo_top_VIA4 $T=38290 115060 0 0 $X=38040 $Y=114830
X5213 2 digital_ldo_top_VIA4 $T=38290 119140 0 0 $X=38040 $Y=118910
X5214 2 digital_ldo_top_VIA4 $T=38290 123220 0 0 $X=38040 $Y=122990
X5215 2 digital_ldo_top_VIA4 $T=38290 127300 0 0 $X=38040 $Y=127070
X5216 3 digital_ldo_top_VIA4 $T=40590 11700 0 0 $X=40340 $Y=11470
X5217 3 digital_ldo_top_VIA4 $T=40590 15780 0 0 $X=40340 $Y=15550
X5218 3 digital_ldo_top_VIA4 $T=40590 19860 0 0 $X=40340 $Y=19630
X5219 3 digital_ldo_top_VIA4 $T=40590 23940 0 0 $X=40340 $Y=23710
X5220 3 digital_ldo_top_VIA4 $T=40590 28020 0 0 $X=40340 $Y=27790
X5221 3 digital_ldo_top_VIA4 $T=40590 32100 0 0 $X=40340 $Y=31870
X5222 3 digital_ldo_top_VIA4 $T=40590 36180 0 0 $X=40340 $Y=35950
X5223 3 digital_ldo_top_VIA4 $T=40590 40260 0 0 $X=40340 $Y=40030
X5224 3 digital_ldo_top_VIA4 $T=40590 44340 0 0 $X=40340 $Y=44110
X5225 3 digital_ldo_top_VIA4 $T=40590 48420 0 0 $X=40340 $Y=48190
X5226 3 digital_ldo_top_VIA4 $T=40590 52500 0 0 $X=40340 $Y=52270
X5227 3 digital_ldo_top_VIA4 $T=40590 56580 0 0 $X=40340 $Y=56350
X5228 3 digital_ldo_top_VIA4 $T=40590 60660 0 0 $X=40340 $Y=60430
X5229 3 digital_ldo_top_VIA4 $T=40590 64740 0 0 $X=40340 $Y=64510
X5230 3 digital_ldo_top_VIA4 $T=40590 68820 0 0 $X=40340 $Y=68590
X5231 3 digital_ldo_top_VIA4 $T=40590 72900 0 0 $X=40340 $Y=72670
X5232 3 digital_ldo_top_VIA4 $T=40590 76980 0 0 $X=40340 $Y=76750
X5233 3 digital_ldo_top_VIA4 $T=40590 81060 0 0 $X=40340 $Y=80830
X5234 3 digital_ldo_top_VIA4 $T=40590 85140 0 0 $X=40340 $Y=84910
X5235 3 digital_ldo_top_VIA4 $T=40590 89220 0 0 $X=40340 $Y=88990
X5236 3 digital_ldo_top_VIA4 $T=40590 93300 0 0 $X=40340 $Y=93070
X5237 3 digital_ldo_top_VIA4 $T=40590 97380 0 0 $X=40340 $Y=97150
X5238 3 digital_ldo_top_VIA4 $T=40590 101460 0 0 $X=40340 $Y=101230
X5239 3 digital_ldo_top_VIA4 $T=40590 105540 0 0 $X=40340 $Y=105310
X5240 3 digital_ldo_top_VIA4 $T=40590 109620 0 0 $X=40340 $Y=109390
X5241 3 digital_ldo_top_VIA4 $T=40590 113700 0 0 $X=40340 $Y=113470
X5242 3 digital_ldo_top_VIA4 $T=40590 117780 0 0 $X=40340 $Y=117550
X5243 3 digital_ldo_top_VIA4 $T=40590 121860 0 0 $X=40340 $Y=121630
X5244 3 digital_ldo_top_VIA4 $T=40590 125940 0 0 $X=40340 $Y=125710
X5245 2 digital_ldo_top_VIA4 $T=41970 13060 0 0 $X=41720 $Y=12830
X5246 2 digital_ldo_top_VIA4 $T=41970 17140 0 0 $X=41720 $Y=16910
X5247 2 digital_ldo_top_VIA4 $T=41970 21220 0 0 $X=41720 $Y=20990
X5248 2 digital_ldo_top_VIA4 $T=41970 25300 0 0 $X=41720 $Y=25070
X5249 2 digital_ldo_top_VIA4 $T=41970 29380 0 0 $X=41720 $Y=29150
X5250 2 digital_ldo_top_VIA4 $T=41970 33460 0 0 $X=41720 $Y=33230
X5251 2 digital_ldo_top_VIA4 $T=41970 37540 0 0 $X=41720 $Y=37310
X5252 2 digital_ldo_top_VIA4 $T=41970 41620 0 0 $X=41720 $Y=41390
X5253 2 digital_ldo_top_VIA4 $T=41970 45700 0 0 $X=41720 $Y=45470
X5254 2 digital_ldo_top_VIA4 $T=41970 49780 0 0 $X=41720 $Y=49550
X5255 2 digital_ldo_top_VIA4 $T=41970 53860 0 0 $X=41720 $Y=53630
X5256 2 digital_ldo_top_VIA4 $T=41970 57940 0 0 $X=41720 $Y=57710
X5257 2 digital_ldo_top_VIA4 $T=41970 62020 0 0 $X=41720 $Y=61790
X5258 2 digital_ldo_top_VIA4 $T=41970 66100 0 0 $X=41720 $Y=65870
X5259 2 digital_ldo_top_VIA4 $T=41970 70180 0 0 $X=41720 $Y=69950
X5260 2 digital_ldo_top_VIA4 $T=41970 74260 0 0 $X=41720 $Y=74030
X5261 2 digital_ldo_top_VIA4 $T=41970 78340 0 0 $X=41720 $Y=78110
X5262 2 digital_ldo_top_VIA4 $T=41970 82420 0 0 $X=41720 $Y=82190
X5263 2 digital_ldo_top_VIA4 $T=41970 86500 0 0 $X=41720 $Y=86270
X5264 2 digital_ldo_top_VIA4 $T=41970 90580 0 0 $X=41720 $Y=90350
X5265 2 digital_ldo_top_VIA4 $T=41970 94660 0 0 $X=41720 $Y=94430
X5266 2 digital_ldo_top_VIA4 $T=41970 98740 0 0 $X=41720 $Y=98510
X5267 2 digital_ldo_top_VIA4 $T=41970 102820 0 0 $X=41720 $Y=102590
X5268 2 digital_ldo_top_VIA4 $T=41970 106900 0 0 $X=41720 $Y=106670
X5269 2 digital_ldo_top_VIA4 $T=41970 110980 0 0 $X=41720 $Y=110750
X5270 2 digital_ldo_top_VIA4 $T=41970 115060 0 0 $X=41720 $Y=114830
X5271 2 digital_ldo_top_VIA4 $T=41970 119140 0 0 $X=41720 $Y=118910
X5272 2 digital_ldo_top_VIA4 $T=41970 123220 0 0 $X=41720 $Y=122990
X5273 2 digital_ldo_top_VIA4 $T=41970 127300 0 0 $X=41720 $Y=127070
X5274 3 digital_ldo_top_VIA4 $T=44270 11700 0 0 $X=44020 $Y=11470
X5275 3 digital_ldo_top_VIA4 $T=44270 15780 0 0 $X=44020 $Y=15550
X5276 3 digital_ldo_top_VIA4 $T=44270 19860 0 0 $X=44020 $Y=19630
X5277 3 digital_ldo_top_VIA4 $T=44270 23940 0 0 $X=44020 $Y=23710
X5278 3 digital_ldo_top_VIA4 $T=44270 28020 0 0 $X=44020 $Y=27790
X5279 3 digital_ldo_top_VIA4 $T=44270 32100 0 0 $X=44020 $Y=31870
X5280 3 digital_ldo_top_VIA4 $T=44270 64740 0 0 $X=44020 $Y=64510
X5281 3 digital_ldo_top_VIA4 $T=44270 68820 0 0 $X=44020 $Y=68590
X5282 3 digital_ldo_top_VIA4 $T=44270 72900 0 0 $X=44020 $Y=72670
X5283 3 digital_ldo_top_VIA4 $T=44270 76980 0 0 $X=44020 $Y=76750
X5284 3 digital_ldo_top_VIA4 $T=44270 81060 0 0 $X=44020 $Y=80830
X5285 3 digital_ldo_top_VIA4 $T=44270 85140 0 0 $X=44020 $Y=84910
X5286 3 digital_ldo_top_VIA4 $T=44270 89220 0 0 $X=44020 $Y=88990
X5287 3 digital_ldo_top_VIA4 $T=44270 93300 0 0 $X=44020 $Y=93070
X5288 3 digital_ldo_top_VIA4 $T=44270 97380 0 0 $X=44020 $Y=97150
X5289 3 digital_ldo_top_VIA4 $T=44270 101460 0 0 $X=44020 $Y=101230
X5290 3 digital_ldo_top_VIA4 $T=44270 105540 0 0 $X=44020 $Y=105310
X5291 3 digital_ldo_top_VIA4 $T=44270 109620 0 0 $X=44020 $Y=109390
X5292 3 digital_ldo_top_VIA4 $T=44270 113700 0 0 $X=44020 $Y=113470
X5293 3 digital_ldo_top_VIA4 $T=44270 117780 0 0 $X=44020 $Y=117550
X5294 3 digital_ldo_top_VIA4 $T=44270 121860 0 0 $X=44020 $Y=121630
X5295 3 digital_ldo_top_VIA4 $T=44270 125940 0 0 $X=44020 $Y=125710
X5296 2 digital_ldo_top_VIA4 $T=45650 13060 0 0 $X=45400 $Y=12830
X5297 2 digital_ldo_top_VIA4 $T=45650 66100 0 0 $X=45400 $Y=65870
X5298 2 digital_ldo_top_VIA4 $T=45650 70180 0 0 $X=45400 $Y=69950
X5299 2 digital_ldo_top_VIA4 $T=45650 74260 0 0 $X=45400 $Y=74030
X5300 2 digital_ldo_top_VIA4 $T=45650 78340 0 0 $X=45400 $Y=78110
X5301 2 digital_ldo_top_VIA4 $T=45650 82420 0 0 $X=45400 $Y=82190
X5302 2 digital_ldo_top_VIA4 $T=45650 86500 0 0 $X=45400 $Y=86270
X5303 2 digital_ldo_top_VIA4 $T=45650 90580 0 0 $X=45400 $Y=90350
X5304 2 digital_ldo_top_VIA4 $T=45650 94660 0 0 $X=45400 $Y=94430
X5305 2 digital_ldo_top_VIA4 $T=45650 98740 0 0 $X=45400 $Y=98510
X5306 2 digital_ldo_top_VIA4 $T=45650 102820 0 0 $X=45400 $Y=102590
X5307 2 digital_ldo_top_VIA4 $T=45650 106900 0 0 $X=45400 $Y=106670
X5308 2 digital_ldo_top_VIA4 $T=45650 110980 0 0 $X=45400 $Y=110750
X5309 2 digital_ldo_top_VIA4 $T=45650 115060 0 0 $X=45400 $Y=114830
X5310 2 digital_ldo_top_VIA4 $T=45650 119140 0 0 $X=45400 $Y=118910
X5311 2 digital_ldo_top_VIA4 $T=45650 123220 0 0 $X=45400 $Y=122990
X5312 2 digital_ldo_top_VIA4 $T=45650 127300 0 0 $X=45400 $Y=127070
X5313 3 digital_ldo_top_VIA4 $T=47950 11700 0 0 $X=47700 $Y=11470
X5314 3 digital_ldo_top_VIA4 $T=47950 15780 0 0 $X=47700 $Y=15550
X5315 3 digital_ldo_top_VIA4 $T=47950 19860 0 0 $X=47700 $Y=19630
X5316 3 digital_ldo_top_VIA4 $T=47950 23940 0 0 $X=47700 $Y=23710
X5317 3 digital_ldo_top_VIA4 $T=47950 28020 0 0 $X=47700 $Y=27790
X5318 3 digital_ldo_top_VIA4 $T=47950 32100 0 0 $X=47700 $Y=31870
X5319 3 digital_ldo_top_VIA4 $T=47950 64740 0 0 $X=47700 $Y=64510
X5320 3 digital_ldo_top_VIA4 $T=47950 68820 0 0 $X=47700 $Y=68590
X5321 3 digital_ldo_top_VIA4 $T=47950 72900 0 0 $X=47700 $Y=72670
X5322 3 digital_ldo_top_VIA4 $T=47950 76980 0 0 $X=47700 $Y=76750
X5323 3 digital_ldo_top_VIA4 $T=47950 81060 0 0 $X=47700 $Y=80830
X5324 3 digital_ldo_top_VIA4 $T=47950 85140 0 0 $X=47700 $Y=84910
X5325 3 digital_ldo_top_VIA4 $T=47950 89220 0 0 $X=47700 $Y=88990
X5326 3 digital_ldo_top_VIA4 $T=47950 93300 0 0 $X=47700 $Y=93070
X5327 3 digital_ldo_top_VIA4 $T=47950 97380 0 0 $X=47700 $Y=97150
X5328 3 digital_ldo_top_VIA4 $T=47950 101460 0 0 $X=47700 $Y=101230
X5329 3 digital_ldo_top_VIA4 $T=47950 105540 0 0 $X=47700 $Y=105310
X5330 3 digital_ldo_top_VIA4 $T=47950 109620 0 0 $X=47700 $Y=109390
X5331 3 digital_ldo_top_VIA4 $T=47950 113700 0 0 $X=47700 $Y=113470
X5332 3 digital_ldo_top_VIA4 $T=47950 117780 0 0 $X=47700 $Y=117550
X5333 3 digital_ldo_top_VIA4 $T=47950 121860 0 0 $X=47700 $Y=121630
X5334 3 digital_ldo_top_VIA4 $T=47950 125940 0 0 $X=47700 $Y=125710
X5335 2 digital_ldo_top_VIA4 $T=49330 13060 0 0 $X=49080 $Y=12830
X5336 2 digital_ldo_top_VIA4 $T=49330 17140 0 0 $X=49080 $Y=16910
X5337 2 digital_ldo_top_VIA4 $T=49330 21220 0 0 $X=49080 $Y=20990
X5338 2 digital_ldo_top_VIA4 $T=49330 25300 0 0 $X=49080 $Y=25070
X5339 2 digital_ldo_top_VIA4 $T=49330 29380 0 0 $X=49080 $Y=29150
X5340 2 digital_ldo_top_VIA4 $T=49330 33460 0 0 $X=49080 $Y=33230
X5341 2 digital_ldo_top_VIA4 $T=49330 37540 0 0 $X=49080 $Y=37310
X5342 2 digital_ldo_top_VIA4 $T=49330 41620 0 0 $X=49080 $Y=41390
X5343 2 digital_ldo_top_VIA4 $T=49330 45700 0 0 $X=49080 $Y=45470
X5344 2 digital_ldo_top_VIA4 $T=49330 49780 0 0 $X=49080 $Y=49550
X5345 2 digital_ldo_top_VIA4 $T=49330 53860 0 0 $X=49080 $Y=53630
X5346 2 digital_ldo_top_VIA4 $T=49330 57940 0 0 $X=49080 $Y=57710
X5347 2 digital_ldo_top_VIA4 $T=49330 62020 0 0 $X=49080 $Y=61790
X5348 2 digital_ldo_top_VIA4 $T=49330 66100 0 0 $X=49080 $Y=65870
X5349 2 digital_ldo_top_VIA4 $T=49330 70180 0 0 $X=49080 $Y=69950
X5350 2 digital_ldo_top_VIA4 $T=49330 74260 0 0 $X=49080 $Y=74030
X5351 2 digital_ldo_top_VIA4 $T=49330 78340 0 0 $X=49080 $Y=78110
X5352 2 digital_ldo_top_VIA4 $T=49330 82420 0 0 $X=49080 $Y=82190
X5353 2 digital_ldo_top_VIA4 $T=49330 86500 0 0 $X=49080 $Y=86270
X5354 2 digital_ldo_top_VIA4 $T=49330 90580 0 0 $X=49080 $Y=90350
X5355 2 digital_ldo_top_VIA4 $T=49330 94660 0 0 $X=49080 $Y=94430
X5356 2 digital_ldo_top_VIA4 $T=49330 98740 0 0 $X=49080 $Y=98510
X5357 2 digital_ldo_top_VIA4 $T=49330 102820 0 0 $X=49080 $Y=102590
X5358 2 digital_ldo_top_VIA4 $T=49330 106900 0 0 $X=49080 $Y=106670
X5359 2 digital_ldo_top_VIA4 $T=49330 110980 0 0 $X=49080 $Y=110750
X5360 2 digital_ldo_top_VIA4 $T=49330 115060 0 0 $X=49080 $Y=114830
X5361 2 digital_ldo_top_VIA4 $T=49330 119140 0 0 $X=49080 $Y=118910
X5362 2 digital_ldo_top_VIA4 $T=49330 123220 0 0 $X=49080 $Y=122990
X5363 2 digital_ldo_top_VIA4 $T=49330 127300 0 0 $X=49080 $Y=127070
X5364 3 digital_ldo_top_VIA4 $T=51630 11700 0 0 $X=51380 $Y=11470
X5365 3 digital_ldo_top_VIA4 $T=51630 15780 0 0 $X=51380 $Y=15550
X5366 3 digital_ldo_top_VIA4 $T=51630 19860 0 0 $X=51380 $Y=19630
X5367 3 digital_ldo_top_VIA4 $T=51630 23940 0 0 $X=51380 $Y=23710
X5368 3 digital_ldo_top_VIA4 $T=51630 28020 0 0 $X=51380 $Y=27790
X5369 3 digital_ldo_top_VIA4 $T=51630 32100 0 0 $X=51380 $Y=31870
X5370 3 digital_ldo_top_VIA4 $T=51630 36180 0 0 $X=51380 $Y=35950
X5371 3 digital_ldo_top_VIA4 $T=51630 40260 0 0 $X=51380 $Y=40030
X5372 3 digital_ldo_top_VIA4 $T=51630 44340 0 0 $X=51380 $Y=44110
X5373 3 digital_ldo_top_VIA4 $T=51630 48420 0 0 $X=51380 $Y=48190
X5374 3 digital_ldo_top_VIA4 $T=51630 52500 0 0 $X=51380 $Y=52270
X5375 3 digital_ldo_top_VIA4 $T=51630 56580 0 0 $X=51380 $Y=56350
X5376 3 digital_ldo_top_VIA4 $T=51630 60660 0 0 $X=51380 $Y=60430
X5377 3 digital_ldo_top_VIA4 $T=51630 64740 0 0 $X=51380 $Y=64510
X5378 3 digital_ldo_top_VIA4 $T=51630 68820 0 0 $X=51380 $Y=68590
X5379 3 digital_ldo_top_VIA4 $T=51630 72900 0 0 $X=51380 $Y=72670
X5380 3 digital_ldo_top_VIA4 $T=51630 76980 0 0 $X=51380 $Y=76750
X5381 3 digital_ldo_top_VIA4 $T=51630 81060 0 0 $X=51380 $Y=80830
X5382 3 digital_ldo_top_VIA4 $T=51630 85140 0 0 $X=51380 $Y=84910
X5383 3 digital_ldo_top_VIA4 $T=51630 89220 0 0 $X=51380 $Y=88990
X5384 3 digital_ldo_top_VIA4 $T=51630 93300 0 0 $X=51380 $Y=93070
X5385 3 digital_ldo_top_VIA4 $T=51630 97380 0 0 $X=51380 $Y=97150
X5386 3 digital_ldo_top_VIA4 $T=51630 101460 0 0 $X=51380 $Y=101230
X5387 3 digital_ldo_top_VIA4 $T=51630 105540 0 0 $X=51380 $Y=105310
X5388 3 digital_ldo_top_VIA4 $T=51630 109620 0 0 $X=51380 $Y=109390
X5389 3 digital_ldo_top_VIA4 $T=51630 113700 0 0 $X=51380 $Y=113470
X5390 3 digital_ldo_top_VIA4 $T=51630 117780 0 0 $X=51380 $Y=117550
X5391 3 digital_ldo_top_VIA4 $T=51630 121860 0 0 $X=51380 $Y=121630
X5392 3 digital_ldo_top_VIA4 $T=51630 125940 0 0 $X=51380 $Y=125710
X5393 2 digital_ldo_top_VIA4 $T=53010 13060 0 0 $X=52760 $Y=12830
X5394 2 digital_ldo_top_VIA4 $T=53010 17140 0 0 $X=52760 $Y=16910
X5395 2 digital_ldo_top_VIA4 $T=53010 21220 0 0 $X=52760 $Y=20990
X5396 2 digital_ldo_top_VIA4 $T=53010 25300 0 0 $X=52760 $Y=25070
X5397 2 digital_ldo_top_VIA4 $T=53010 29380 0 0 $X=52760 $Y=29150
X5398 2 digital_ldo_top_VIA4 $T=53010 33460 0 0 $X=52760 $Y=33230
X5399 2 digital_ldo_top_VIA4 $T=53010 37540 0 0 $X=52760 $Y=37310
X5400 2 digital_ldo_top_VIA4 $T=53010 41620 0 0 $X=52760 $Y=41390
X5401 2 digital_ldo_top_VIA4 $T=53010 45700 0 0 $X=52760 $Y=45470
X5402 2 digital_ldo_top_VIA4 $T=53010 49780 0 0 $X=52760 $Y=49550
X5403 2 digital_ldo_top_VIA4 $T=53010 53860 0 0 $X=52760 $Y=53630
X5404 2 digital_ldo_top_VIA4 $T=53010 57940 0 0 $X=52760 $Y=57710
X5405 2 digital_ldo_top_VIA4 $T=53010 62020 0 0 $X=52760 $Y=61790
X5406 2 digital_ldo_top_VIA4 $T=53010 66100 0 0 $X=52760 $Y=65870
X5407 2 digital_ldo_top_VIA4 $T=53010 70180 0 0 $X=52760 $Y=69950
X5408 2 digital_ldo_top_VIA4 $T=53010 74260 0 0 $X=52760 $Y=74030
X5409 2 digital_ldo_top_VIA4 $T=53010 78340 0 0 $X=52760 $Y=78110
X5410 2 digital_ldo_top_VIA4 $T=53010 82420 0 0 $X=52760 $Y=82190
X5411 2 digital_ldo_top_VIA4 $T=53010 86500 0 0 $X=52760 $Y=86270
X5412 2 digital_ldo_top_VIA4 $T=53010 90580 0 0 $X=52760 $Y=90350
X5413 2 digital_ldo_top_VIA4 $T=53010 94660 0 0 $X=52760 $Y=94430
X5414 2 digital_ldo_top_VIA4 $T=53010 98740 0 0 $X=52760 $Y=98510
X5415 2 digital_ldo_top_VIA4 $T=53010 102820 0 0 $X=52760 $Y=102590
X5416 2 digital_ldo_top_VIA4 $T=53010 106900 0 0 $X=52760 $Y=106670
X5417 2 digital_ldo_top_VIA4 $T=53010 110980 0 0 $X=52760 $Y=110750
X5418 2 digital_ldo_top_VIA4 $T=53010 115060 0 0 $X=52760 $Y=114830
X5419 2 digital_ldo_top_VIA4 $T=53010 119140 0 0 $X=52760 $Y=118910
X5420 2 digital_ldo_top_VIA4 $T=53010 123220 0 0 $X=52760 $Y=122990
X5421 2 digital_ldo_top_VIA4 $T=53010 127300 0 0 $X=52760 $Y=127070
X5422 3 digital_ldo_top_VIA4 $T=55310 11700 0 0 $X=55060 $Y=11470
X5423 3 digital_ldo_top_VIA4 $T=55310 15780 0 0 $X=55060 $Y=15550
X5424 3 digital_ldo_top_VIA4 $T=55310 19860 0 0 $X=55060 $Y=19630
X5425 3 digital_ldo_top_VIA4 $T=55310 23940 0 0 $X=55060 $Y=23710
X5426 3 digital_ldo_top_VIA4 $T=55310 28020 0 0 $X=55060 $Y=27790
X5427 3 digital_ldo_top_VIA4 $T=55310 32100 0 0 $X=55060 $Y=31870
X5428 3 digital_ldo_top_VIA4 $T=55310 36180 0 0 $X=55060 $Y=35950
X5429 3 digital_ldo_top_VIA4 $T=55310 40260 0 0 $X=55060 $Y=40030
X5430 3 digital_ldo_top_VIA4 $T=55310 44340 0 0 $X=55060 $Y=44110
X5431 3 digital_ldo_top_VIA4 $T=55310 48420 0 0 $X=55060 $Y=48190
X5432 3 digital_ldo_top_VIA4 $T=55310 52500 0 0 $X=55060 $Y=52270
X5433 3 digital_ldo_top_VIA4 $T=55310 56580 0 0 $X=55060 $Y=56350
X5434 3 digital_ldo_top_VIA4 $T=55310 60660 0 0 $X=55060 $Y=60430
X5435 3 digital_ldo_top_VIA4 $T=55310 64740 0 0 $X=55060 $Y=64510
X5436 3 digital_ldo_top_VIA4 $T=55310 68820 0 0 $X=55060 $Y=68590
X5437 3 digital_ldo_top_VIA4 $T=55310 72900 0 0 $X=55060 $Y=72670
X5438 3 digital_ldo_top_VIA4 $T=55310 76980 0 0 $X=55060 $Y=76750
X5439 3 digital_ldo_top_VIA4 $T=55310 81060 0 0 $X=55060 $Y=80830
X5440 3 digital_ldo_top_VIA4 $T=55310 85140 0 0 $X=55060 $Y=84910
X5441 3 digital_ldo_top_VIA4 $T=55310 89220 0 0 $X=55060 $Y=88990
X5442 3 digital_ldo_top_VIA4 $T=55310 93300 0 0 $X=55060 $Y=93070
X5443 3 digital_ldo_top_VIA4 $T=55310 97380 0 0 $X=55060 $Y=97150
X5444 3 digital_ldo_top_VIA4 $T=55310 101460 0 0 $X=55060 $Y=101230
X5445 3 digital_ldo_top_VIA4 $T=55310 105540 0 0 $X=55060 $Y=105310
X5446 3 digital_ldo_top_VIA4 $T=55310 109620 0 0 $X=55060 $Y=109390
X5447 3 digital_ldo_top_VIA4 $T=55310 113700 0 0 $X=55060 $Y=113470
X5448 3 digital_ldo_top_VIA4 $T=55310 117780 0 0 $X=55060 $Y=117550
X5449 3 digital_ldo_top_VIA4 $T=55310 121860 0 0 $X=55060 $Y=121630
X5450 3 digital_ldo_top_VIA4 $T=55310 125940 0 0 $X=55060 $Y=125710
X5451 2 digital_ldo_top_VIA4 $T=56690 13060 0 0 $X=56440 $Y=12830
X5452 2 digital_ldo_top_VIA4 $T=56690 17140 0 0 $X=56440 $Y=16910
X5453 2 digital_ldo_top_VIA4 $T=56690 21220 0 0 $X=56440 $Y=20990
X5454 2 digital_ldo_top_VIA4 $T=56690 25300 0 0 $X=56440 $Y=25070
X5455 2 digital_ldo_top_VIA4 $T=56690 29380 0 0 $X=56440 $Y=29150
X5456 2 digital_ldo_top_VIA4 $T=56690 33460 0 0 $X=56440 $Y=33230
X5457 2 digital_ldo_top_VIA4 $T=56690 37540 0 0 $X=56440 $Y=37310
X5458 2 digital_ldo_top_VIA4 $T=56690 41620 0 0 $X=56440 $Y=41390
X5459 2 digital_ldo_top_VIA4 $T=56690 45700 0 0 $X=56440 $Y=45470
X5460 2 digital_ldo_top_VIA4 $T=56690 49780 0 0 $X=56440 $Y=49550
X5461 2 digital_ldo_top_VIA4 $T=56690 53860 0 0 $X=56440 $Y=53630
X5462 2 digital_ldo_top_VIA4 $T=56690 57940 0 0 $X=56440 $Y=57710
X5463 2 digital_ldo_top_VIA4 $T=56690 62020 0 0 $X=56440 $Y=61790
X5464 2 digital_ldo_top_VIA4 $T=56690 66100 0 0 $X=56440 $Y=65870
X5465 2 digital_ldo_top_VIA4 $T=56690 70180 0 0 $X=56440 $Y=69950
X5466 2 digital_ldo_top_VIA4 $T=56690 74260 0 0 $X=56440 $Y=74030
X5467 2 digital_ldo_top_VIA4 $T=56690 78340 0 0 $X=56440 $Y=78110
X5468 2 digital_ldo_top_VIA4 $T=56690 82420 0 0 $X=56440 $Y=82190
X5469 2 digital_ldo_top_VIA4 $T=56690 86500 0 0 $X=56440 $Y=86270
X5470 2 digital_ldo_top_VIA4 $T=56690 90580 0 0 $X=56440 $Y=90350
X5471 2 digital_ldo_top_VIA4 $T=56690 94660 0 0 $X=56440 $Y=94430
X5472 2 digital_ldo_top_VIA4 $T=56690 98740 0 0 $X=56440 $Y=98510
X5473 2 digital_ldo_top_VIA4 $T=56690 102820 0 0 $X=56440 $Y=102590
X5474 2 digital_ldo_top_VIA4 $T=56690 106900 0 0 $X=56440 $Y=106670
X5475 2 digital_ldo_top_VIA4 $T=56690 110980 0 0 $X=56440 $Y=110750
X5476 2 digital_ldo_top_VIA4 $T=56690 115060 0 0 $X=56440 $Y=114830
X5477 2 digital_ldo_top_VIA4 $T=56690 119140 0 0 $X=56440 $Y=118910
X5478 2 digital_ldo_top_VIA4 $T=56690 123220 0 0 $X=56440 $Y=122990
X5479 2 digital_ldo_top_VIA4 $T=56690 127300 0 0 $X=56440 $Y=127070
X5480 3 digital_ldo_top_VIA4 $T=58990 11700 0 0 $X=58740 $Y=11470
X5481 3 digital_ldo_top_VIA4 $T=58990 36180 0 0 $X=58740 $Y=35950
X5482 3 digital_ldo_top_VIA4 $T=58990 40260 0 0 $X=58740 $Y=40030
X5483 3 digital_ldo_top_VIA4 $T=58990 44340 0 0 $X=58740 $Y=44110
X5484 3 digital_ldo_top_VIA4 $T=58990 48420 0 0 $X=58740 $Y=48190
X5485 3 digital_ldo_top_VIA4 $T=58990 52500 0 0 $X=58740 $Y=52270
X5486 3 digital_ldo_top_VIA4 $T=58990 56580 0 0 $X=58740 $Y=56350
X5487 3 digital_ldo_top_VIA4 $T=58990 60660 0 0 $X=58740 $Y=60430
X5488 3 digital_ldo_top_VIA4 $T=58990 64740 0 0 $X=58740 $Y=64510
X5489 3 digital_ldo_top_VIA4 $T=58990 68820 0 0 $X=58740 $Y=68590
X5490 3 digital_ldo_top_VIA4 $T=58990 72900 0 0 $X=58740 $Y=72670
X5491 3 digital_ldo_top_VIA4 $T=58990 76980 0 0 $X=58740 $Y=76750
X5492 3 digital_ldo_top_VIA4 $T=58990 81060 0 0 $X=58740 $Y=80830
X5493 3 digital_ldo_top_VIA4 $T=58990 85140 0 0 $X=58740 $Y=84910
X5494 3 digital_ldo_top_VIA4 $T=58990 89220 0 0 $X=58740 $Y=88990
X5495 3 digital_ldo_top_VIA4 $T=58990 93300 0 0 $X=58740 $Y=93070
X5496 3 digital_ldo_top_VIA4 $T=58990 97380 0 0 $X=58740 $Y=97150
X5497 3 digital_ldo_top_VIA4 $T=58990 101460 0 0 $X=58740 $Y=101230
X5498 3 digital_ldo_top_VIA4 $T=58990 105540 0 0 $X=58740 $Y=105310
X5499 3 digital_ldo_top_VIA4 $T=58990 109620 0 0 $X=58740 $Y=109390
X5500 3 digital_ldo_top_VIA4 $T=58990 113700 0 0 $X=58740 $Y=113470
X5501 3 digital_ldo_top_VIA4 $T=58990 117780 0 0 $X=58740 $Y=117550
X5502 3 digital_ldo_top_VIA4 $T=58990 121860 0 0 $X=58740 $Y=121630
X5503 3 digital_ldo_top_VIA4 $T=58990 125940 0 0 $X=58740 $Y=125710
X5504 2 digital_ldo_top_VIA4 $T=60370 13060 0 0 $X=60120 $Y=12830
X5505 2 digital_ldo_top_VIA4 $T=60370 33460 0 0 $X=60120 $Y=33230
X5506 2 digital_ldo_top_VIA4 $T=60370 37540 0 0 $X=60120 $Y=37310
X5507 2 digital_ldo_top_VIA4 $T=60370 41620 0 0 $X=60120 $Y=41390
X5508 2 digital_ldo_top_VIA4 $T=60370 45700 0 0 $X=60120 $Y=45470
X5509 2 digital_ldo_top_VIA4 $T=60370 49780 0 0 $X=60120 $Y=49550
X5510 2 digital_ldo_top_VIA4 $T=60370 53860 0 0 $X=60120 $Y=53630
X5511 2 digital_ldo_top_VIA4 $T=60370 57940 0 0 $X=60120 $Y=57710
X5512 2 digital_ldo_top_VIA4 $T=60370 62020 0 0 $X=60120 $Y=61790
X5513 2 digital_ldo_top_VIA4 $T=60370 66100 0 0 $X=60120 $Y=65870
X5514 2 digital_ldo_top_VIA4 $T=60370 70180 0 0 $X=60120 $Y=69950
X5515 2 digital_ldo_top_VIA4 $T=60370 74260 0 0 $X=60120 $Y=74030
X5516 2 digital_ldo_top_VIA4 $T=60370 78340 0 0 $X=60120 $Y=78110
X5517 2 digital_ldo_top_VIA4 $T=60370 82420 0 0 $X=60120 $Y=82190
X5518 2 digital_ldo_top_VIA4 $T=60370 86500 0 0 $X=60120 $Y=86270
X5519 2 digital_ldo_top_VIA4 $T=60370 90580 0 0 $X=60120 $Y=90350
X5520 2 digital_ldo_top_VIA4 $T=60370 94660 0 0 $X=60120 $Y=94430
X5521 2 digital_ldo_top_VIA4 $T=60370 98740 0 0 $X=60120 $Y=98510
X5522 2 digital_ldo_top_VIA4 $T=60370 102820 0 0 $X=60120 $Y=102590
X5523 2 digital_ldo_top_VIA4 $T=60370 106900 0 0 $X=60120 $Y=106670
X5524 2 digital_ldo_top_VIA4 $T=60370 110980 0 0 $X=60120 $Y=110750
X5525 2 digital_ldo_top_VIA4 $T=60370 115060 0 0 $X=60120 $Y=114830
X5526 2 digital_ldo_top_VIA4 $T=60370 119140 0 0 $X=60120 $Y=118910
X5527 2 digital_ldo_top_VIA4 $T=60370 123220 0 0 $X=60120 $Y=122990
X5528 2 digital_ldo_top_VIA4 $T=60370 127300 0 0 $X=60120 $Y=127070
X5529 3 digital_ldo_top_VIA4 $T=62670 11700 0 0 $X=62420 $Y=11470
X5530 3 digital_ldo_top_VIA4 $T=62670 36180 0 0 $X=62420 $Y=35950
X5531 3 digital_ldo_top_VIA4 $T=62670 40260 0 0 $X=62420 $Y=40030
X5532 3 digital_ldo_top_VIA4 $T=62670 44340 0 0 $X=62420 $Y=44110
X5533 3 digital_ldo_top_VIA4 $T=62670 48420 0 0 $X=62420 $Y=48190
X5534 3 digital_ldo_top_VIA4 $T=62670 52500 0 0 $X=62420 $Y=52270
X5535 3 digital_ldo_top_VIA4 $T=62670 56580 0 0 $X=62420 $Y=56350
X5536 3 digital_ldo_top_VIA4 $T=62670 60660 0 0 $X=62420 $Y=60430
X5537 3 digital_ldo_top_VIA4 $T=62670 64740 0 0 $X=62420 $Y=64510
X5538 3 digital_ldo_top_VIA4 $T=62670 68820 0 0 $X=62420 $Y=68590
X5539 3 digital_ldo_top_VIA4 $T=62670 72900 0 0 $X=62420 $Y=72670
X5540 3 digital_ldo_top_VIA4 $T=62670 76980 0 0 $X=62420 $Y=76750
X5541 3 digital_ldo_top_VIA4 $T=62670 81060 0 0 $X=62420 $Y=80830
X5542 3 digital_ldo_top_VIA4 $T=62670 85140 0 0 $X=62420 $Y=84910
X5543 3 digital_ldo_top_VIA4 $T=62670 89220 0 0 $X=62420 $Y=88990
X5544 3 digital_ldo_top_VIA4 $T=62670 93300 0 0 $X=62420 $Y=93070
X5545 3 digital_ldo_top_VIA4 $T=62670 97380 0 0 $X=62420 $Y=97150
X5546 3 digital_ldo_top_VIA4 $T=62670 101460 0 0 $X=62420 $Y=101230
X5547 3 digital_ldo_top_VIA4 $T=62670 105540 0 0 $X=62420 $Y=105310
X5548 3 digital_ldo_top_VIA4 $T=62670 109620 0 0 $X=62420 $Y=109390
X5549 3 digital_ldo_top_VIA4 $T=62670 113700 0 0 $X=62420 $Y=113470
X5550 3 digital_ldo_top_VIA4 $T=62670 117780 0 0 $X=62420 $Y=117550
X5551 3 digital_ldo_top_VIA4 $T=62670 121860 0 0 $X=62420 $Y=121630
X5552 3 digital_ldo_top_VIA4 $T=62670 125940 0 0 $X=62420 $Y=125710
X5553 2 digital_ldo_top_VIA4 $T=64050 13060 0 0 $X=63800 $Y=12830
X5554 2 digital_ldo_top_VIA4 $T=64050 33460 0 0 $X=63800 $Y=33230
X5555 2 digital_ldo_top_VIA4 $T=64050 37540 0 0 $X=63800 $Y=37310
X5556 2 digital_ldo_top_VIA4 $T=64050 41620 0 0 $X=63800 $Y=41390
X5557 2 digital_ldo_top_VIA4 $T=64050 45700 0 0 $X=63800 $Y=45470
X5558 2 digital_ldo_top_VIA4 $T=64050 49780 0 0 $X=63800 $Y=49550
X5559 2 digital_ldo_top_VIA4 $T=64050 53860 0 0 $X=63800 $Y=53630
X5560 2 digital_ldo_top_VIA4 $T=64050 57940 0 0 $X=63800 $Y=57710
X5561 2 digital_ldo_top_VIA4 $T=64050 62020 0 0 $X=63800 $Y=61790
X5562 2 digital_ldo_top_VIA4 $T=64050 66100 0 0 $X=63800 $Y=65870
X5563 2 digital_ldo_top_VIA4 $T=64050 70180 0 0 $X=63800 $Y=69950
X5564 2 digital_ldo_top_VIA4 $T=64050 74260 0 0 $X=63800 $Y=74030
X5565 2 digital_ldo_top_VIA4 $T=64050 78340 0 0 $X=63800 $Y=78110
X5566 2 digital_ldo_top_VIA4 $T=64050 82420 0 0 $X=63800 $Y=82190
X5567 2 digital_ldo_top_VIA4 $T=64050 86500 0 0 $X=63800 $Y=86270
X5568 2 digital_ldo_top_VIA4 $T=64050 90580 0 0 $X=63800 $Y=90350
X5569 2 digital_ldo_top_VIA4 $T=64050 94660 0 0 $X=63800 $Y=94430
X5570 2 digital_ldo_top_VIA4 $T=64050 98740 0 0 $X=63800 $Y=98510
X5571 2 digital_ldo_top_VIA4 $T=64050 102820 0 0 $X=63800 $Y=102590
X5572 2 digital_ldo_top_VIA4 $T=64050 106900 0 0 $X=63800 $Y=106670
X5573 2 digital_ldo_top_VIA4 $T=64050 110980 0 0 $X=63800 $Y=110750
X5574 2 digital_ldo_top_VIA4 $T=64050 115060 0 0 $X=63800 $Y=114830
X5575 2 digital_ldo_top_VIA4 $T=64050 119140 0 0 $X=63800 $Y=118910
X5576 2 digital_ldo_top_VIA4 $T=64050 123220 0 0 $X=63800 $Y=122990
X5577 2 digital_ldo_top_VIA4 $T=64050 127300 0 0 $X=63800 $Y=127070
X5578 3 digital_ldo_top_VIA4 $T=66350 11700 0 0 $X=66100 $Y=11470
X5579 3 digital_ldo_top_VIA4 $T=66350 36180 0 0 $X=66100 $Y=35950
X5580 3 digital_ldo_top_VIA4 $T=66350 40260 0 0 $X=66100 $Y=40030
X5581 3 digital_ldo_top_VIA4 $T=66350 44340 0 0 $X=66100 $Y=44110
X5582 3 digital_ldo_top_VIA4 $T=66350 48420 0 0 $X=66100 $Y=48190
X5583 3 digital_ldo_top_VIA4 $T=66350 52500 0 0 $X=66100 $Y=52270
X5584 3 digital_ldo_top_VIA4 $T=66350 56580 0 0 $X=66100 $Y=56350
X5585 3 digital_ldo_top_VIA4 $T=66350 60660 0 0 $X=66100 $Y=60430
X5586 3 digital_ldo_top_VIA4 $T=66350 64740 0 0 $X=66100 $Y=64510
X5587 3 digital_ldo_top_VIA4 $T=66350 68820 0 0 $X=66100 $Y=68590
X5588 3 digital_ldo_top_VIA4 $T=66350 72900 0 0 $X=66100 $Y=72670
X5589 3 digital_ldo_top_VIA4 $T=66350 76980 0 0 $X=66100 $Y=76750
X5590 3 digital_ldo_top_VIA4 $T=66350 81060 0 0 $X=66100 $Y=80830
X5591 3 digital_ldo_top_VIA4 $T=66350 85140 0 0 $X=66100 $Y=84910
X5592 3 digital_ldo_top_VIA4 $T=66350 89220 0 0 $X=66100 $Y=88990
X5593 3 digital_ldo_top_VIA4 $T=66350 93300 0 0 $X=66100 $Y=93070
X5594 3 digital_ldo_top_VIA4 $T=66350 97380 0 0 $X=66100 $Y=97150
X5595 3 digital_ldo_top_VIA4 $T=66350 101460 0 0 $X=66100 $Y=101230
X5596 3 digital_ldo_top_VIA4 $T=66350 105540 0 0 $X=66100 $Y=105310
X5597 3 digital_ldo_top_VIA4 $T=66350 109620 0 0 $X=66100 $Y=109390
X5598 3 digital_ldo_top_VIA4 $T=66350 113700 0 0 $X=66100 $Y=113470
X5599 3 digital_ldo_top_VIA4 $T=66350 117780 0 0 $X=66100 $Y=117550
X5600 3 digital_ldo_top_VIA4 $T=66350 121860 0 0 $X=66100 $Y=121630
X5601 3 digital_ldo_top_VIA4 $T=66350 125940 0 0 $X=66100 $Y=125710
X5602 2 digital_ldo_top_VIA4 $T=67730 13060 0 0 $X=67480 $Y=12830
X5603 2 digital_ldo_top_VIA4 $T=67730 33460 0 0 $X=67480 $Y=33230
X5604 2 digital_ldo_top_VIA4 $T=67730 37540 0 0 $X=67480 $Y=37310
X5605 2 digital_ldo_top_VIA4 $T=67730 41620 0 0 $X=67480 $Y=41390
X5606 2 digital_ldo_top_VIA4 $T=67730 45700 0 0 $X=67480 $Y=45470
X5607 2 digital_ldo_top_VIA4 $T=67730 49780 0 0 $X=67480 $Y=49550
X5608 2 digital_ldo_top_VIA4 $T=67730 53860 0 0 $X=67480 $Y=53630
X5609 2 digital_ldo_top_VIA4 $T=67730 57940 0 0 $X=67480 $Y=57710
X5610 2 digital_ldo_top_VIA4 $T=67730 62020 0 0 $X=67480 $Y=61790
X5611 2 digital_ldo_top_VIA4 $T=67730 66100 0 0 $X=67480 $Y=65870
X5612 2 digital_ldo_top_VIA4 $T=67730 70180 0 0 $X=67480 $Y=69950
X5613 2 digital_ldo_top_VIA4 $T=67730 74260 0 0 $X=67480 $Y=74030
X5614 2 digital_ldo_top_VIA4 $T=67730 78340 0 0 $X=67480 $Y=78110
X5615 2 digital_ldo_top_VIA4 $T=67730 82420 0 0 $X=67480 $Y=82190
X5616 2 digital_ldo_top_VIA4 $T=67730 86500 0 0 $X=67480 $Y=86270
X5617 2 digital_ldo_top_VIA4 $T=67730 90580 0 0 $X=67480 $Y=90350
X5618 2 digital_ldo_top_VIA4 $T=67730 94660 0 0 $X=67480 $Y=94430
X5619 2 digital_ldo_top_VIA4 $T=67730 98740 0 0 $X=67480 $Y=98510
X5620 2 digital_ldo_top_VIA4 $T=67730 102820 0 0 $X=67480 $Y=102590
X5621 2 digital_ldo_top_VIA4 $T=67730 106900 0 0 $X=67480 $Y=106670
X5622 2 digital_ldo_top_VIA4 $T=67730 110980 0 0 $X=67480 $Y=110750
X5623 2 digital_ldo_top_VIA4 $T=67730 115060 0 0 $X=67480 $Y=114830
X5624 2 digital_ldo_top_VIA4 $T=67730 119140 0 0 $X=67480 $Y=118910
X5625 2 digital_ldo_top_VIA4 $T=67730 123220 0 0 $X=67480 $Y=122990
X5626 2 digital_ldo_top_VIA4 $T=67730 127300 0 0 $X=67480 $Y=127070
X5627 3 digital_ldo_top_VIA4 $T=70030 11700 0 0 $X=69780 $Y=11470
X5628 3 digital_ldo_top_VIA4 $T=70030 36180 0 0 $X=69780 $Y=35950
X5629 3 digital_ldo_top_VIA4 $T=70030 40260 0 0 $X=69780 $Y=40030
X5630 3 digital_ldo_top_VIA4 $T=70030 44340 0 0 $X=69780 $Y=44110
X5631 3 digital_ldo_top_VIA4 $T=70030 48420 0 0 $X=69780 $Y=48190
X5632 3 digital_ldo_top_VIA4 $T=70030 52500 0 0 $X=69780 $Y=52270
X5633 3 digital_ldo_top_VIA4 $T=70030 56580 0 0 $X=69780 $Y=56350
X5634 3 digital_ldo_top_VIA4 $T=70030 60660 0 0 $X=69780 $Y=60430
X5635 3 digital_ldo_top_VIA4 $T=70030 64740 0 0 $X=69780 $Y=64510
X5636 3 digital_ldo_top_VIA4 $T=70030 68820 0 0 $X=69780 $Y=68590
X5637 3 digital_ldo_top_VIA4 $T=70030 72900 0 0 $X=69780 $Y=72670
X5638 3 digital_ldo_top_VIA4 $T=70030 76980 0 0 $X=69780 $Y=76750
X5639 3 digital_ldo_top_VIA4 $T=70030 81060 0 0 $X=69780 $Y=80830
X5640 3 digital_ldo_top_VIA4 $T=70030 85140 0 0 $X=69780 $Y=84910
X5641 3 digital_ldo_top_VIA4 $T=70030 89220 0 0 $X=69780 $Y=88990
X5642 3 digital_ldo_top_VIA4 $T=70030 93300 0 0 $X=69780 $Y=93070
X5643 3 digital_ldo_top_VIA4 $T=70030 97380 0 0 $X=69780 $Y=97150
X5644 3 digital_ldo_top_VIA4 $T=70030 101460 0 0 $X=69780 $Y=101230
X5645 3 digital_ldo_top_VIA4 $T=70030 105540 0 0 $X=69780 $Y=105310
X5646 3 digital_ldo_top_VIA4 $T=70030 109620 0 0 $X=69780 $Y=109390
X5647 3 digital_ldo_top_VIA4 $T=70030 113700 0 0 $X=69780 $Y=113470
X5648 3 digital_ldo_top_VIA4 $T=70030 117780 0 0 $X=69780 $Y=117550
X5649 3 digital_ldo_top_VIA4 $T=70030 121860 0 0 $X=69780 $Y=121630
X5650 3 digital_ldo_top_VIA4 $T=70030 125940 0 0 $X=69780 $Y=125710
X5651 2 digital_ldo_top_VIA4 $T=71410 13060 0 0 $X=71160 $Y=12830
X5652 2 digital_ldo_top_VIA4 $T=71410 33460 0 0 $X=71160 $Y=33230
X5653 2 digital_ldo_top_VIA4 $T=71410 37540 0 0 $X=71160 $Y=37310
X5654 2 digital_ldo_top_VIA4 $T=71410 41620 0 0 $X=71160 $Y=41390
X5655 2 digital_ldo_top_VIA4 $T=71410 45700 0 0 $X=71160 $Y=45470
X5656 2 digital_ldo_top_VIA4 $T=71410 49780 0 0 $X=71160 $Y=49550
X5657 2 digital_ldo_top_VIA4 $T=71410 53860 0 0 $X=71160 $Y=53630
X5658 2 digital_ldo_top_VIA4 $T=71410 57940 0 0 $X=71160 $Y=57710
X5659 2 digital_ldo_top_VIA4 $T=71410 62020 0 0 $X=71160 $Y=61790
X5660 2 digital_ldo_top_VIA4 $T=71410 66100 0 0 $X=71160 $Y=65870
X5661 2 digital_ldo_top_VIA4 $T=71410 70180 0 0 $X=71160 $Y=69950
X5662 2 digital_ldo_top_VIA4 $T=71410 74260 0 0 $X=71160 $Y=74030
X5663 2 digital_ldo_top_VIA4 $T=71410 78340 0 0 $X=71160 $Y=78110
X5664 2 digital_ldo_top_VIA4 $T=71410 82420 0 0 $X=71160 $Y=82190
X5665 2 digital_ldo_top_VIA4 $T=71410 86500 0 0 $X=71160 $Y=86270
X5666 2 digital_ldo_top_VIA4 $T=71410 90580 0 0 $X=71160 $Y=90350
X5667 2 digital_ldo_top_VIA4 $T=71410 94660 0 0 $X=71160 $Y=94430
X5668 2 digital_ldo_top_VIA4 $T=71410 98740 0 0 $X=71160 $Y=98510
X5669 2 digital_ldo_top_VIA4 $T=71410 102820 0 0 $X=71160 $Y=102590
X5670 2 digital_ldo_top_VIA4 $T=71410 106900 0 0 $X=71160 $Y=106670
X5671 2 digital_ldo_top_VIA4 $T=71410 110980 0 0 $X=71160 $Y=110750
X5672 2 digital_ldo_top_VIA4 $T=71410 115060 0 0 $X=71160 $Y=114830
X5673 2 digital_ldo_top_VIA4 $T=71410 119140 0 0 $X=71160 $Y=118910
X5674 2 digital_ldo_top_VIA4 $T=71410 123220 0 0 $X=71160 $Y=122990
X5675 2 digital_ldo_top_VIA4 $T=71410 127300 0 0 $X=71160 $Y=127070
X5676 3 digital_ldo_top_VIA4 $T=73710 11700 0 0 $X=73460 $Y=11470
X5677 3 digital_ldo_top_VIA4 $T=73710 36180 0 0 $X=73460 $Y=35950
X5678 3 digital_ldo_top_VIA4 $T=73710 40260 0 0 $X=73460 $Y=40030
X5679 3 digital_ldo_top_VIA4 $T=73710 44340 0 0 $X=73460 $Y=44110
X5680 3 digital_ldo_top_VIA4 $T=73710 48420 0 0 $X=73460 $Y=48190
X5681 3 digital_ldo_top_VIA4 $T=73710 52500 0 0 $X=73460 $Y=52270
X5682 3 digital_ldo_top_VIA4 $T=73710 56580 0 0 $X=73460 $Y=56350
X5683 3 digital_ldo_top_VIA4 $T=73710 60660 0 0 $X=73460 $Y=60430
X5684 3 digital_ldo_top_VIA4 $T=73710 64740 0 0 $X=73460 $Y=64510
X5685 3 digital_ldo_top_VIA4 $T=73710 68820 0 0 $X=73460 $Y=68590
X5686 3 digital_ldo_top_VIA4 $T=73710 72900 0 0 $X=73460 $Y=72670
X5687 3 digital_ldo_top_VIA4 $T=73710 76980 0 0 $X=73460 $Y=76750
X5688 3 digital_ldo_top_VIA4 $T=73710 81060 0 0 $X=73460 $Y=80830
X5689 3 digital_ldo_top_VIA4 $T=73710 85140 0 0 $X=73460 $Y=84910
X5690 3 digital_ldo_top_VIA4 $T=73710 89220 0 0 $X=73460 $Y=88990
X5691 3 digital_ldo_top_VIA4 $T=73710 93300 0 0 $X=73460 $Y=93070
X5692 3 digital_ldo_top_VIA4 $T=73710 97380 0 0 $X=73460 $Y=97150
X5693 3 digital_ldo_top_VIA4 $T=73710 101460 0 0 $X=73460 $Y=101230
X5694 3 digital_ldo_top_VIA4 $T=73710 105540 0 0 $X=73460 $Y=105310
X5695 3 digital_ldo_top_VIA4 $T=73710 109620 0 0 $X=73460 $Y=109390
X5696 3 digital_ldo_top_VIA4 $T=73710 113700 0 0 $X=73460 $Y=113470
X5697 3 digital_ldo_top_VIA4 $T=73710 117780 0 0 $X=73460 $Y=117550
X5698 3 digital_ldo_top_VIA4 $T=73710 121860 0 0 $X=73460 $Y=121630
X5699 3 digital_ldo_top_VIA4 $T=73710 125940 0 0 $X=73460 $Y=125710
X5700 2 digital_ldo_top_VIA4 $T=75090 13060 0 0 $X=74840 $Y=12830
X5701 2 digital_ldo_top_VIA4 $T=75090 33460 0 0 $X=74840 $Y=33230
X5702 2 digital_ldo_top_VIA4 $T=75090 37540 0 0 $X=74840 $Y=37310
X5703 2 digital_ldo_top_VIA4 $T=75090 41620 0 0 $X=74840 $Y=41390
X5704 2 digital_ldo_top_VIA4 $T=75090 45700 0 0 $X=74840 $Y=45470
X5705 2 digital_ldo_top_VIA4 $T=75090 49780 0 0 $X=74840 $Y=49550
X5706 2 digital_ldo_top_VIA4 $T=75090 53860 0 0 $X=74840 $Y=53630
X5707 2 digital_ldo_top_VIA4 $T=75090 57940 0 0 $X=74840 $Y=57710
X5708 2 digital_ldo_top_VIA4 $T=75090 62020 0 0 $X=74840 $Y=61790
X5709 2 digital_ldo_top_VIA4 $T=75090 66100 0 0 $X=74840 $Y=65870
X5710 2 digital_ldo_top_VIA4 $T=75090 70180 0 0 $X=74840 $Y=69950
X5711 2 digital_ldo_top_VIA4 $T=75090 74260 0 0 $X=74840 $Y=74030
X5712 2 digital_ldo_top_VIA4 $T=75090 78340 0 0 $X=74840 $Y=78110
X5713 2 digital_ldo_top_VIA4 $T=75090 82420 0 0 $X=74840 $Y=82190
X5714 2 digital_ldo_top_VIA4 $T=75090 86500 0 0 $X=74840 $Y=86270
X5715 2 digital_ldo_top_VIA4 $T=75090 90580 0 0 $X=74840 $Y=90350
X5716 2 digital_ldo_top_VIA4 $T=75090 94660 0 0 $X=74840 $Y=94430
X5717 2 digital_ldo_top_VIA4 $T=75090 98740 0 0 $X=74840 $Y=98510
X5718 2 digital_ldo_top_VIA4 $T=75090 102820 0 0 $X=74840 $Y=102590
X5719 2 digital_ldo_top_VIA4 $T=75090 106900 0 0 $X=74840 $Y=106670
X5720 2 digital_ldo_top_VIA4 $T=75090 110980 0 0 $X=74840 $Y=110750
X5721 2 digital_ldo_top_VIA4 $T=75090 115060 0 0 $X=74840 $Y=114830
X5722 2 digital_ldo_top_VIA4 $T=75090 119140 0 0 $X=74840 $Y=118910
X5723 2 digital_ldo_top_VIA4 $T=75090 123220 0 0 $X=74840 $Y=122990
X5724 2 digital_ldo_top_VIA4 $T=75090 127300 0 0 $X=74840 $Y=127070
X5725 3 digital_ldo_top_VIA4 $T=77390 11700 0 0 $X=77140 $Y=11470
X5726 3 digital_ldo_top_VIA4 $T=77390 44340 0 0 $X=77140 $Y=44110
X5727 3 digital_ldo_top_VIA4 $T=77390 48420 0 0 $X=77140 $Y=48190
X5728 3 digital_ldo_top_VIA4 $T=77390 52500 0 0 $X=77140 $Y=52270
X5729 3 digital_ldo_top_VIA4 $T=77390 56580 0 0 $X=77140 $Y=56350
X5730 3 digital_ldo_top_VIA4 $T=77390 60660 0 0 $X=77140 $Y=60430
X5731 3 digital_ldo_top_VIA4 $T=77390 64740 0 0 $X=77140 $Y=64510
X5732 3 digital_ldo_top_VIA4 $T=77390 68820 0 0 $X=77140 $Y=68590
X5733 3 digital_ldo_top_VIA4 $T=77390 72900 0 0 $X=77140 $Y=72670
X5734 3 digital_ldo_top_VIA4 $T=77390 76980 0 0 $X=77140 $Y=76750
X5735 3 digital_ldo_top_VIA4 $T=77390 81060 0 0 $X=77140 $Y=80830
X5736 3 digital_ldo_top_VIA4 $T=77390 85140 0 0 $X=77140 $Y=84910
X5737 3 digital_ldo_top_VIA4 $T=77390 89220 0 0 $X=77140 $Y=88990
X5738 3 digital_ldo_top_VIA4 $T=77390 93300 0 0 $X=77140 $Y=93070
X5739 3 digital_ldo_top_VIA4 $T=77390 97380 0 0 $X=77140 $Y=97150
X5740 3 digital_ldo_top_VIA4 $T=77390 101460 0 0 $X=77140 $Y=101230
X5741 3 digital_ldo_top_VIA4 $T=77390 105540 0 0 $X=77140 $Y=105310
X5742 3 digital_ldo_top_VIA4 $T=77390 109620 0 0 $X=77140 $Y=109390
X5743 3 digital_ldo_top_VIA4 $T=77390 113700 0 0 $X=77140 $Y=113470
X5744 3 digital_ldo_top_VIA4 $T=77390 117780 0 0 $X=77140 $Y=117550
X5745 3 digital_ldo_top_VIA4 $T=77390 121860 0 0 $X=77140 $Y=121630
X5746 3 digital_ldo_top_VIA4 $T=77390 125940 0 0 $X=77140 $Y=125710
X5747 2 digital_ldo_top_VIA4 $T=78770 13060 0 0 $X=78520 $Y=12830
X5748 2 digital_ldo_top_VIA4 $T=78770 45700 0 0 $X=78520 $Y=45470
X5749 2 digital_ldo_top_VIA4 $T=78770 49780 0 0 $X=78520 $Y=49550
X5750 2 digital_ldo_top_VIA4 $T=78770 53860 0 0 $X=78520 $Y=53630
X5751 2 digital_ldo_top_VIA4 $T=78770 57940 0 0 $X=78520 $Y=57710
X5752 2 digital_ldo_top_VIA4 $T=78770 62020 0 0 $X=78520 $Y=61790
X5753 2 digital_ldo_top_VIA4 $T=78770 66100 0 0 $X=78520 $Y=65870
X5754 2 digital_ldo_top_VIA4 $T=78770 70180 0 0 $X=78520 $Y=69950
X5755 2 digital_ldo_top_VIA4 $T=78770 74260 0 0 $X=78520 $Y=74030
X5756 2 digital_ldo_top_VIA4 $T=78770 78340 0 0 $X=78520 $Y=78110
X5757 2 digital_ldo_top_VIA4 $T=78770 82420 0 0 $X=78520 $Y=82190
X5758 2 digital_ldo_top_VIA4 $T=78770 86500 0 0 $X=78520 $Y=86270
X5759 2 digital_ldo_top_VIA4 $T=78770 90580 0 0 $X=78520 $Y=90350
X5760 2 digital_ldo_top_VIA4 $T=78770 94660 0 0 $X=78520 $Y=94430
X5761 2 digital_ldo_top_VIA4 $T=78770 98740 0 0 $X=78520 $Y=98510
X5762 2 digital_ldo_top_VIA4 $T=78770 102820 0 0 $X=78520 $Y=102590
X5763 2 digital_ldo_top_VIA4 $T=78770 106900 0 0 $X=78520 $Y=106670
X5764 2 digital_ldo_top_VIA4 $T=78770 110980 0 0 $X=78520 $Y=110750
X5765 2 digital_ldo_top_VIA4 $T=78770 115060 0 0 $X=78520 $Y=114830
X5766 2 digital_ldo_top_VIA4 $T=78770 119140 0 0 $X=78520 $Y=118910
X5767 2 digital_ldo_top_VIA4 $T=78770 123220 0 0 $X=78520 $Y=122990
X5768 2 digital_ldo_top_VIA4 $T=78770 127300 0 0 $X=78520 $Y=127070
X5769 3 digital_ldo_top_VIA4 $T=81070 11700 0 0 $X=80820 $Y=11470
X5770 3 digital_ldo_top_VIA4 $T=81070 44340 0 0 $X=80820 $Y=44110
X5771 3 digital_ldo_top_VIA4 $T=81070 48420 0 0 $X=80820 $Y=48190
X5772 3 digital_ldo_top_VIA4 $T=81070 52500 0 0 $X=80820 $Y=52270
X5773 3 digital_ldo_top_VIA4 $T=81070 56580 0 0 $X=80820 $Y=56350
X5774 3 digital_ldo_top_VIA4 $T=81070 60660 0 0 $X=80820 $Y=60430
X5775 3 digital_ldo_top_VIA4 $T=81070 64740 0 0 $X=80820 $Y=64510
X5776 3 digital_ldo_top_VIA4 $T=81070 68820 0 0 $X=80820 $Y=68590
X5777 3 digital_ldo_top_VIA4 $T=81070 72900 0 0 $X=80820 $Y=72670
X5778 3 digital_ldo_top_VIA4 $T=81070 76980 0 0 $X=80820 $Y=76750
X5779 3 digital_ldo_top_VIA4 $T=81070 81060 0 0 $X=80820 $Y=80830
X5780 3 digital_ldo_top_VIA4 $T=81070 85140 0 0 $X=80820 $Y=84910
X5781 3 digital_ldo_top_VIA4 $T=81070 89220 0 0 $X=80820 $Y=88990
X5782 3 digital_ldo_top_VIA4 $T=81070 93300 0 0 $X=80820 $Y=93070
X5783 3 digital_ldo_top_VIA4 $T=81070 97380 0 0 $X=80820 $Y=97150
X5784 3 digital_ldo_top_VIA4 $T=81070 101460 0 0 $X=80820 $Y=101230
X5785 3 digital_ldo_top_VIA4 $T=81070 105540 0 0 $X=80820 $Y=105310
X5786 3 digital_ldo_top_VIA4 $T=81070 109620 0 0 $X=80820 $Y=109390
X5787 3 digital_ldo_top_VIA4 $T=81070 113700 0 0 $X=80820 $Y=113470
X5788 3 digital_ldo_top_VIA4 $T=81070 117780 0 0 $X=80820 $Y=117550
X5789 3 digital_ldo_top_VIA4 $T=81070 121860 0 0 $X=80820 $Y=121630
X5790 3 digital_ldo_top_VIA4 $T=81070 125940 0 0 $X=80820 $Y=125710
X5791 2 digital_ldo_top_VIA4 $T=82450 13060 0 0 $X=82200 $Y=12830
X5792 2 digital_ldo_top_VIA4 $T=82450 45700 0 0 $X=82200 $Y=45470
X5793 2 digital_ldo_top_VIA4 $T=82450 49780 0 0 $X=82200 $Y=49550
X5794 2 digital_ldo_top_VIA4 $T=82450 53860 0 0 $X=82200 $Y=53630
X5795 2 digital_ldo_top_VIA4 $T=82450 57940 0 0 $X=82200 $Y=57710
X5796 2 digital_ldo_top_VIA4 $T=82450 62020 0 0 $X=82200 $Y=61790
X5797 2 digital_ldo_top_VIA4 $T=82450 66100 0 0 $X=82200 $Y=65870
X5798 2 digital_ldo_top_VIA4 $T=82450 70180 0 0 $X=82200 $Y=69950
X5799 2 digital_ldo_top_VIA4 $T=82450 74260 0 0 $X=82200 $Y=74030
X5800 2 digital_ldo_top_VIA4 $T=82450 78340 0 0 $X=82200 $Y=78110
X5801 2 digital_ldo_top_VIA4 $T=82450 82420 0 0 $X=82200 $Y=82190
X5802 2 digital_ldo_top_VIA4 $T=82450 86500 0 0 $X=82200 $Y=86270
X5803 2 digital_ldo_top_VIA4 $T=82450 90580 0 0 $X=82200 $Y=90350
X5804 2 digital_ldo_top_VIA4 $T=82450 94660 0 0 $X=82200 $Y=94430
X5805 2 digital_ldo_top_VIA4 $T=82450 98740 0 0 $X=82200 $Y=98510
X5806 2 digital_ldo_top_VIA4 $T=82450 102820 0 0 $X=82200 $Y=102590
X5807 2 digital_ldo_top_VIA4 $T=82450 106900 0 0 $X=82200 $Y=106670
X5808 2 digital_ldo_top_VIA4 $T=82450 110980 0 0 $X=82200 $Y=110750
X5809 2 digital_ldo_top_VIA4 $T=82450 115060 0 0 $X=82200 $Y=114830
X5810 2 digital_ldo_top_VIA4 $T=82450 119140 0 0 $X=82200 $Y=118910
X5811 2 digital_ldo_top_VIA4 $T=82450 123220 0 0 $X=82200 $Y=122990
X5812 2 digital_ldo_top_VIA4 $T=82450 127300 0 0 $X=82200 $Y=127070
X5813 3 digital_ldo_top_VIA4 $T=84750 11700 0 0 $X=84500 $Y=11470
X5814 3 digital_ldo_top_VIA4 $T=84750 44340 0 0 $X=84500 $Y=44110
X5815 3 digital_ldo_top_VIA4 $T=84750 48420 0 0 $X=84500 $Y=48190
X5816 3 digital_ldo_top_VIA4 $T=84750 52500 0 0 $X=84500 $Y=52270
X5817 3 digital_ldo_top_VIA4 $T=84750 56580 0 0 $X=84500 $Y=56350
X5818 3 digital_ldo_top_VIA4 $T=84750 60660 0 0 $X=84500 $Y=60430
X5819 3 digital_ldo_top_VIA4 $T=84750 64740 0 0 $X=84500 $Y=64510
X5820 3 digital_ldo_top_VIA4 $T=84750 68820 0 0 $X=84500 $Y=68590
X5821 3 digital_ldo_top_VIA4 $T=84750 72900 0 0 $X=84500 $Y=72670
X5822 3 digital_ldo_top_VIA4 $T=84750 76980 0 0 $X=84500 $Y=76750
X5823 3 digital_ldo_top_VIA4 $T=84750 81060 0 0 $X=84500 $Y=80830
X5824 3 digital_ldo_top_VIA4 $T=84750 85140 0 0 $X=84500 $Y=84910
X5825 3 digital_ldo_top_VIA4 $T=84750 89220 0 0 $X=84500 $Y=88990
X5826 3 digital_ldo_top_VIA4 $T=84750 93300 0 0 $X=84500 $Y=93070
X5827 3 digital_ldo_top_VIA4 $T=84750 97380 0 0 $X=84500 $Y=97150
X5828 3 digital_ldo_top_VIA4 $T=84750 101460 0 0 $X=84500 $Y=101230
X5829 3 digital_ldo_top_VIA4 $T=84750 105540 0 0 $X=84500 $Y=105310
X5830 3 digital_ldo_top_VIA4 $T=84750 109620 0 0 $X=84500 $Y=109390
X5831 3 digital_ldo_top_VIA4 $T=84750 113700 0 0 $X=84500 $Y=113470
X5832 3 digital_ldo_top_VIA4 $T=84750 117780 0 0 $X=84500 $Y=117550
X5833 3 digital_ldo_top_VIA4 $T=84750 121860 0 0 $X=84500 $Y=121630
X5834 3 digital_ldo_top_VIA4 $T=84750 125940 0 0 $X=84500 $Y=125710
X5835 2 digital_ldo_top_VIA4 $T=86130 13060 0 0 $X=85880 $Y=12830
X5836 2 digital_ldo_top_VIA4 $T=86130 45700 0 0 $X=85880 $Y=45470
X5837 2 digital_ldo_top_VIA4 $T=86130 49780 0 0 $X=85880 $Y=49550
X5838 2 digital_ldo_top_VIA4 $T=86130 53860 0 0 $X=85880 $Y=53630
X5839 2 digital_ldo_top_VIA4 $T=86130 57940 0 0 $X=85880 $Y=57710
X5840 2 digital_ldo_top_VIA4 $T=86130 62020 0 0 $X=85880 $Y=61790
X5841 2 digital_ldo_top_VIA4 $T=86130 66100 0 0 $X=85880 $Y=65870
X5842 2 digital_ldo_top_VIA4 $T=86130 70180 0 0 $X=85880 $Y=69950
X5843 2 digital_ldo_top_VIA4 $T=86130 74260 0 0 $X=85880 $Y=74030
X5844 2 digital_ldo_top_VIA4 $T=86130 78340 0 0 $X=85880 $Y=78110
X5845 2 digital_ldo_top_VIA4 $T=86130 82420 0 0 $X=85880 $Y=82190
X5846 2 digital_ldo_top_VIA4 $T=86130 86500 0 0 $X=85880 $Y=86270
X5847 2 digital_ldo_top_VIA4 $T=86130 90580 0 0 $X=85880 $Y=90350
X5848 2 digital_ldo_top_VIA4 $T=86130 94660 0 0 $X=85880 $Y=94430
X5849 2 digital_ldo_top_VIA4 $T=86130 98740 0 0 $X=85880 $Y=98510
X5850 2 digital_ldo_top_VIA4 $T=86130 102820 0 0 $X=85880 $Y=102590
X5851 2 digital_ldo_top_VIA4 $T=86130 106900 0 0 $X=85880 $Y=106670
X5852 2 digital_ldo_top_VIA4 $T=86130 110980 0 0 $X=85880 $Y=110750
X5853 2 digital_ldo_top_VIA4 $T=86130 115060 0 0 $X=85880 $Y=114830
X5854 2 digital_ldo_top_VIA4 $T=86130 119140 0 0 $X=85880 $Y=118910
X5855 2 digital_ldo_top_VIA4 $T=86130 123220 0 0 $X=85880 $Y=122990
X5856 2 digital_ldo_top_VIA4 $T=86130 127300 0 0 $X=85880 $Y=127070
X5857 3 digital_ldo_top_VIA4 $T=88430 11700 0 0 $X=88180 $Y=11470
X5858 3 digital_ldo_top_VIA4 $T=88430 44340 0 0 $X=88180 $Y=44110
X5859 3 digital_ldo_top_VIA4 $T=88430 48420 0 0 $X=88180 $Y=48190
X5860 3 digital_ldo_top_VIA4 $T=88430 52500 0 0 $X=88180 $Y=52270
X5861 3 digital_ldo_top_VIA4 $T=88430 56580 0 0 $X=88180 $Y=56350
X5862 3 digital_ldo_top_VIA4 $T=88430 60660 0 0 $X=88180 $Y=60430
X5863 3 digital_ldo_top_VIA4 $T=88430 64740 0 0 $X=88180 $Y=64510
X5864 3 digital_ldo_top_VIA4 $T=88430 68820 0 0 $X=88180 $Y=68590
X5865 3 digital_ldo_top_VIA4 $T=88430 72900 0 0 $X=88180 $Y=72670
X5866 3 digital_ldo_top_VIA4 $T=88430 76980 0 0 $X=88180 $Y=76750
X5867 3 digital_ldo_top_VIA4 $T=88430 81060 0 0 $X=88180 $Y=80830
X5868 3 digital_ldo_top_VIA4 $T=88430 85140 0 0 $X=88180 $Y=84910
X5869 3 digital_ldo_top_VIA4 $T=88430 89220 0 0 $X=88180 $Y=88990
X5870 3 digital_ldo_top_VIA4 $T=88430 93300 0 0 $X=88180 $Y=93070
X5871 3 digital_ldo_top_VIA4 $T=88430 97380 0 0 $X=88180 $Y=97150
X5872 3 digital_ldo_top_VIA4 $T=88430 101460 0 0 $X=88180 $Y=101230
X5873 3 digital_ldo_top_VIA4 $T=88430 105540 0 0 $X=88180 $Y=105310
X5874 3 digital_ldo_top_VIA4 $T=88430 109620 0 0 $X=88180 $Y=109390
X5875 3 digital_ldo_top_VIA4 $T=88430 113700 0 0 $X=88180 $Y=113470
X5876 3 digital_ldo_top_VIA4 $T=88430 117780 0 0 $X=88180 $Y=117550
X5877 3 digital_ldo_top_VIA4 $T=88430 121860 0 0 $X=88180 $Y=121630
X5878 3 digital_ldo_top_VIA4 $T=88430 125940 0 0 $X=88180 $Y=125710
X5879 2 digital_ldo_top_VIA4 $T=89810 13060 0 0 $X=89560 $Y=12830
X5880 2 digital_ldo_top_VIA4 $T=89810 45700 0 0 $X=89560 $Y=45470
X5881 2 digital_ldo_top_VIA4 $T=89810 49780 0 0 $X=89560 $Y=49550
X5882 2 digital_ldo_top_VIA4 $T=89810 53860 0 0 $X=89560 $Y=53630
X5883 2 digital_ldo_top_VIA4 $T=89810 57940 0 0 $X=89560 $Y=57710
X5884 2 digital_ldo_top_VIA4 $T=89810 62020 0 0 $X=89560 $Y=61790
X5885 2 digital_ldo_top_VIA4 $T=89810 66100 0 0 $X=89560 $Y=65870
X5886 2 digital_ldo_top_VIA4 $T=89810 70180 0 0 $X=89560 $Y=69950
X5887 2 digital_ldo_top_VIA4 $T=89810 74260 0 0 $X=89560 $Y=74030
X5888 2 digital_ldo_top_VIA4 $T=89810 78340 0 0 $X=89560 $Y=78110
X5889 2 digital_ldo_top_VIA4 $T=89810 82420 0 0 $X=89560 $Y=82190
X5890 2 digital_ldo_top_VIA4 $T=89810 86500 0 0 $X=89560 $Y=86270
X5891 2 digital_ldo_top_VIA4 $T=89810 90580 0 0 $X=89560 $Y=90350
X5892 2 digital_ldo_top_VIA4 $T=89810 94660 0 0 $X=89560 $Y=94430
X5893 2 digital_ldo_top_VIA4 $T=89810 98740 0 0 $X=89560 $Y=98510
X5894 2 digital_ldo_top_VIA4 $T=89810 102820 0 0 $X=89560 $Y=102590
X5895 2 digital_ldo_top_VIA4 $T=89810 106900 0 0 $X=89560 $Y=106670
X5896 2 digital_ldo_top_VIA4 $T=89810 110980 0 0 $X=89560 $Y=110750
X5897 2 digital_ldo_top_VIA4 $T=89810 115060 0 0 $X=89560 $Y=114830
X5898 2 digital_ldo_top_VIA4 $T=89810 119140 0 0 $X=89560 $Y=118910
X5899 2 digital_ldo_top_VIA4 $T=89810 123220 0 0 $X=89560 $Y=122990
X5900 2 digital_ldo_top_VIA4 $T=89810 127300 0 0 $X=89560 $Y=127070
X5901 3 digital_ldo_top_VIA4 $T=92110 11700 0 0 $X=91860 $Y=11470
X5902 3 digital_ldo_top_VIA4 $T=92110 15780 0 0 $X=91860 $Y=15550
X5903 3 digital_ldo_top_VIA4 $T=92110 19860 0 0 $X=91860 $Y=19630
X5904 3 digital_ldo_top_VIA4 $T=92110 23940 0 0 $X=91860 $Y=23710
X5905 3 digital_ldo_top_VIA4 $T=92110 28020 0 0 $X=91860 $Y=27790
X5906 3 digital_ldo_top_VIA4 $T=92110 32100 0 0 $X=91860 $Y=31870
X5907 3 digital_ldo_top_VIA4 $T=92110 36180 0 0 $X=91860 $Y=35950
X5908 3 digital_ldo_top_VIA4 $T=92110 40260 0 0 $X=91860 $Y=40030
X5909 3 digital_ldo_top_VIA4 $T=92110 44340 0 0 $X=91860 $Y=44110
X5910 3 digital_ldo_top_VIA4 $T=92110 48420 0 0 $X=91860 $Y=48190
X5911 3 digital_ldo_top_VIA4 $T=92110 52500 0 0 $X=91860 $Y=52270
X5912 3 digital_ldo_top_VIA4 $T=92110 56580 0 0 $X=91860 $Y=56350
X5913 3 digital_ldo_top_VIA4 $T=92110 60660 0 0 $X=91860 $Y=60430
X5914 3 digital_ldo_top_VIA4 $T=92110 64740 0 0 $X=91860 $Y=64510
X5915 3 digital_ldo_top_VIA4 $T=92110 68820 0 0 $X=91860 $Y=68590
X5916 3 digital_ldo_top_VIA4 $T=92110 72900 0 0 $X=91860 $Y=72670
X5917 3 digital_ldo_top_VIA4 $T=92110 76980 0 0 $X=91860 $Y=76750
X5918 3 digital_ldo_top_VIA4 $T=92110 81060 0 0 $X=91860 $Y=80830
X5919 3 digital_ldo_top_VIA4 $T=92110 85140 0 0 $X=91860 $Y=84910
X5920 3 digital_ldo_top_VIA4 $T=92110 89220 0 0 $X=91860 $Y=88990
X5921 3 digital_ldo_top_VIA4 $T=92110 93300 0 0 $X=91860 $Y=93070
X5922 3 digital_ldo_top_VIA4 $T=92110 97380 0 0 $X=91860 $Y=97150
X5923 3 digital_ldo_top_VIA4 $T=92110 101460 0 0 $X=91860 $Y=101230
X5924 3 digital_ldo_top_VIA4 $T=92110 105540 0 0 $X=91860 $Y=105310
X5925 3 digital_ldo_top_VIA4 $T=92110 109620 0 0 $X=91860 $Y=109390
X5926 3 digital_ldo_top_VIA4 $T=92110 113700 0 0 $X=91860 $Y=113470
X5927 3 digital_ldo_top_VIA4 $T=92110 117780 0 0 $X=91860 $Y=117550
X5928 3 digital_ldo_top_VIA4 $T=92110 121860 0 0 $X=91860 $Y=121630
X5929 3 digital_ldo_top_VIA4 $T=92110 125940 0 0 $X=91860 $Y=125710
X5930 2 digital_ldo_top_VIA4 $T=93490 13060 0 0 $X=93240 $Y=12830
X5931 2 digital_ldo_top_VIA4 $T=93490 17140 0 0 $X=93240 $Y=16910
X5932 2 digital_ldo_top_VIA4 $T=93490 21220 0 0 $X=93240 $Y=20990
X5933 2 digital_ldo_top_VIA4 $T=93490 25300 0 0 $X=93240 $Y=25070
X5934 2 digital_ldo_top_VIA4 $T=93490 29380 0 0 $X=93240 $Y=29150
X5935 2 digital_ldo_top_VIA4 $T=93490 33460 0 0 $X=93240 $Y=33230
X5936 2 digital_ldo_top_VIA4 $T=93490 37540 0 0 $X=93240 $Y=37310
X5937 2 digital_ldo_top_VIA4 $T=93490 41620 0 0 $X=93240 $Y=41390
X5938 2 digital_ldo_top_VIA4 $T=93490 45700 0 0 $X=93240 $Y=45470
X5939 2 digital_ldo_top_VIA4 $T=93490 49780 0 0 $X=93240 $Y=49550
X5940 2 digital_ldo_top_VIA4 $T=93490 53860 0 0 $X=93240 $Y=53630
X5941 2 digital_ldo_top_VIA4 $T=93490 57940 0 0 $X=93240 $Y=57710
X5942 2 digital_ldo_top_VIA4 $T=93490 62020 0 0 $X=93240 $Y=61790
X5943 2 digital_ldo_top_VIA4 $T=93490 66100 0 0 $X=93240 $Y=65870
X5944 2 digital_ldo_top_VIA4 $T=93490 70180 0 0 $X=93240 $Y=69950
X5945 2 digital_ldo_top_VIA4 $T=93490 74260 0 0 $X=93240 $Y=74030
X5946 2 digital_ldo_top_VIA4 $T=93490 78340 0 0 $X=93240 $Y=78110
X5947 2 digital_ldo_top_VIA4 $T=93490 82420 0 0 $X=93240 $Y=82190
X5948 2 digital_ldo_top_VIA4 $T=93490 86500 0 0 $X=93240 $Y=86270
X5949 2 digital_ldo_top_VIA4 $T=93490 90580 0 0 $X=93240 $Y=90350
X5950 2 digital_ldo_top_VIA4 $T=93490 94660 0 0 $X=93240 $Y=94430
X5951 2 digital_ldo_top_VIA4 $T=93490 98740 0 0 $X=93240 $Y=98510
X5952 2 digital_ldo_top_VIA4 $T=93490 102820 0 0 $X=93240 $Y=102590
X5953 2 digital_ldo_top_VIA4 $T=93490 106900 0 0 $X=93240 $Y=106670
X5954 2 digital_ldo_top_VIA4 $T=93490 110980 0 0 $X=93240 $Y=110750
X5955 2 digital_ldo_top_VIA4 $T=93490 115060 0 0 $X=93240 $Y=114830
X5956 2 digital_ldo_top_VIA4 $T=93490 119140 0 0 $X=93240 $Y=118910
X5957 2 digital_ldo_top_VIA4 $T=93490 123220 0 0 $X=93240 $Y=122990
X5958 2 digital_ldo_top_VIA4 $T=93490 127300 0 0 $X=93240 $Y=127070
X5959 3 digital_ldo_top_VIA4 $T=95790 11700 0 0 $X=95540 $Y=11470
X5960 3 digital_ldo_top_VIA4 $T=95790 15780 0 0 $X=95540 $Y=15550
X5961 3 digital_ldo_top_VIA4 $T=95790 19860 0 0 $X=95540 $Y=19630
X5962 3 digital_ldo_top_VIA4 $T=95790 23940 0 0 $X=95540 $Y=23710
X5963 3 digital_ldo_top_VIA4 $T=95790 28020 0 0 $X=95540 $Y=27790
X5964 3 digital_ldo_top_VIA4 $T=95790 32100 0 0 $X=95540 $Y=31870
X5965 3 digital_ldo_top_VIA4 $T=95790 36180 0 0 $X=95540 $Y=35950
X5966 3 digital_ldo_top_VIA4 $T=95790 40260 0 0 $X=95540 $Y=40030
X5967 3 digital_ldo_top_VIA4 $T=95790 44340 0 0 $X=95540 $Y=44110
X5968 3 digital_ldo_top_VIA4 $T=95790 48420 0 0 $X=95540 $Y=48190
X5969 3 digital_ldo_top_VIA4 $T=95790 52500 0 0 $X=95540 $Y=52270
X5970 3 digital_ldo_top_VIA4 $T=95790 56580 0 0 $X=95540 $Y=56350
X5971 3 digital_ldo_top_VIA4 $T=95790 60660 0 0 $X=95540 $Y=60430
X5972 3 digital_ldo_top_VIA4 $T=95790 64740 0 0 $X=95540 $Y=64510
X5973 3 digital_ldo_top_VIA4 $T=95790 68820 0 0 $X=95540 $Y=68590
X5974 3 digital_ldo_top_VIA4 $T=95790 72900 0 0 $X=95540 $Y=72670
X5975 3 digital_ldo_top_VIA4 $T=95790 76980 0 0 $X=95540 $Y=76750
X5976 3 digital_ldo_top_VIA4 $T=95790 81060 0 0 $X=95540 $Y=80830
X5977 3 digital_ldo_top_VIA4 $T=95790 85140 0 0 $X=95540 $Y=84910
X5978 3 digital_ldo_top_VIA4 $T=95790 89220 0 0 $X=95540 $Y=88990
X5979 3 digital_ldo_top_VIA4 $T=95790 93300 0 0 $X=95540 $Y=93070
X5980 3 digital_ldo_top_VIA4 $T=95790 97380 0 0 $X=95540 $Y=97150
X5981 3 digital_ldo_top_VIA4 $T=95790 101460 0 0 $X=95540 $Y=101230
X5982 3 digital_ldo_top_VIA4 $T=95790 105540 0 0 $X=95540 $Y=105310
X5983 3 digital_ldo_top_VIA4 $T=95790 109620 0 0 $X=95540 $Y=109390
X5984 3 digital_ldo_top_VIA4 $T=95790 113700 0 0 $X=95540 $Y=113470
X5985 3 digital_ldo_top_VIA4 $T=95790 117780 0 0 $X=95540 $Y=117550
X5986 3 digital_ldo_top_VIA4 $T=95790 121860 0 0 $X=95540 $Y=121630
X5987 3 digital_ldo_top_VIA4 $T=95790 125940 0 0 $X=95540 $Y=125710
X5988 2 digital_ldo_top_VIA4 $T=97170 13060 0 0 $X=96920 $Y=12830
X5989 2 digital_ldo_top_VIA4 $T=97170 17140 0 0 $X=96920 $Y=16910
X5990 2 digital_ldo_top_VIA4 $T=97170 21220 0 0 $X=96920 $Y=20990
X5991 2 digital_ldo_top_VIA4 $T=97170 25300 0 0 $X=96920 $Y=25070
X5992 2 digital_ldo_top_VIA4 $T=97170 29380 0 0 $X=96920 $Y=29150
X5993 2 digital_ldo_top_VIA4 $T=97170 33460 0 0 $X=96920 $Y=33230
X5994 2 digital_ldo_top_VIA4 $T=97170 37540 0 0 $X=96920 $Y=37310
X5995 2 digital_ldo_top_VIA4 $T=97170 41620 0 0 $X=96920 $Y=41390
X5996 2 digital_ldo_top_VIA4 $T=97170 45700 0 0 $X=96920 $Y=45470
X5997 2 digital_ldo_top_VIA4 $T=97170 49780 0 0 $X=96920 $Y=49550
X5998 2 digital_ldo_top_VIA4 $T=97170 53860 0 0 $X=96920 $Y=53630
X5999 2 digital_ldo_top_VIA4 $T=97170 57940 0 0 $X=96920 $Y=57710
X6000 2 digital_ldo_top_VIA4 $T=97170 62020 0 0 $X=96920 $Y=61790
X6001 2 digital_ldo_top_VIA4 $T=97170 66100 0 0 $X=96920 $Y=65870
X6002 2 digital_ldo_top_VIA4 $T=97170 70180 0 0 $X=96920 $Y=69950
X6003 2 digital_ldo_top_VIA4 $T=97170 74260 0 0 $X=96920 $Y=74030
X6004 2 digital_ldo_top_VIA4 $T=97170 78340 0 0 $X=96920 $Y=78110
X6005 2 digital_ldo_top_VIA4 $T=97170 82420 0 0 $X=96920 $Y=82190
X6006 2 digital_ldo_top_VIA4 $T=97170 86500 0 0 $X=96920 $Y=86270
X6007 2 digital_ldo_top_VIA4 $T=97170 90580 0 0 $X=96920 $Y=90350
X6008 2 digital_ldo_top_VIA4 $T=97170 94660 0 0 $X=96920 $Y=94430
X6009 2 digital_ldo_top_VIA4 $T=97170 98740 0 0 $X=96920 $Y=98510
X6010 2 digital_ldo_top_VIA4 $T=97170 102820 0 0 $X=96920 $Y=102590
X6011 2 digital_ldo_top_VIA4 $T=97170 106900 0 0 $X=96920 $Y=106670
X6012 2 digital_ldo_top_VIA4 $T=97170 110980 0 0 $X=96920 $Y=110750
X6013 2 digital_ldo_top_VIA4 $T=97170 115060 0 0 $X=96920 $Y=114830
X6014 2 digital_ldo_top_VIA4 $T=97170 119140 0 0 $X=96920 $Y=118910
X6015 2 digital_ldo_top_VIA4 $T=97170 123220 0 0 $X=96920 $Y=122990
X6016 2 digital_ldo_top_VIA4 $T=97170 127300 0 0 $X=96920 $Y=127070
X6017 3 digital_ldo_top_VIA4 $T=99470 11700 0 0 $X=99220 $Y=11470
X6018 3 digital_ldo_top_VIA4 $T=99470 15780 0 0 $X=99220 $Y=15550
X6019 3 digital_ldo_top_VIA4 $T=99470 19860 0 0 $X=99220 $Y=19630
X6020 3 digital_ldo_top_VIA4 $T=99470 23940 0 0 $X=99220 $Y=23710
X6021 3 digital_ldo_top_VIA4 $T=99470 28020 0 0 $X=99220 $Y=27790
X6022 3 digital_ldo_top_VIA4 $T=99470 32100 0 0 $X=99220 $Y=31870
X6023 3 digital_ldo_top_VIA4 $T=99470 36180 0 0 $X=99220 $Y=35950
X6024 3 digital_ldo_top_VIA4 $T=99470 40260 0 0 $X=99220 $Y=40030
X6025 3 digital_ldo_top_VIA4 $T=99470 44340 0 0 $X=99220 $Y=44110
X6026 3 digital_ldo_top_VIA4 $T=99470 48420 0 0 $X=99220 $Y=48190
X6027 3 digital_ldo_top_VIA4 $T=99470 52500 0 0 $X=99220 $Y=52270
X6028 3 digital_ldo_top_VIA4 $T=99470 56580 0 0 $X=99220 $Y=56350
X6029 3 digital_ldo_top_VIA4 $T=99470 60660 0 0 $X=99220 $Y=60430
X6030 3 digital_ldo_top_VIA4 $T=99470 64740 0 0 $X=99220 $Y=64510
X6031 3 digital_ldo_top_VIA4 $T=99470 68820 0 0 $X=99220 $Y=68590
X6032 3 digital_ldo_top_VIA4 $T=99470 72900 0 0 $X=99220 $Y=72670
X6033 3 digital_ldo_top_VIA4 $T=99470 76980 0 0 $X=99220 $Y=76750
X6034 3 digital_ldo_top_VIA4 $T=99470 81060 0 0 $X=99220 $Y=80830
X6035 3 digital_ldo_top_VIA4 $T=99470 85140 0 0 $X=99220 $Y=84910
X6036 3 digital_ldo_top_VIA4 $T=99470 89220 0 0 $X=99220 $Y=88990
X6037 3 digital_ldo_top_VIA4 $T=99470 93300 0 0 $X=99220 $Y=93070
X6038 3 digital_ldo_top_VIA4 $T=99470 97380 0 0 $X=99220 $Y=97150
X6039 3 digital_ldo_top_VIA4 $T=99470 101460 0 0 $X=99220 $Y=101230
X6040 3 digital_ldo_top_VIA4 $T=99470 105540 0 0 $X=99220 $Y=105310
X6041 3 digital_ldo_top_VIA4 $T=99470 109620 0 0 $X=99220 $Y=109390
X6042 3 digital_ldo_top_VIA4 $T=99470 113700 0 0 $X=99220 $Y=113470
X6043 3 digital_ldo_top_VIA4 $T=99470 117780 0 0 $X=99220 $Y=117550
X6044 3 digital_ldo_top_VIA4 $T=99470 121860 0 0 $X=99220 $Y=121630
X6045 3 digital_ldo_top_VIA4 $T=99470 125940 0 0 $X=99220 $Y=125710
X6046 2 digital_ldo_top_VIA4 $T=100850 13060 0 0 $X=100600 $Y=12830
X6047 2 digital_ldo_top_VIA4 $T=100850 17140 0 0 $X=100600 $Y=16910
X6048 2 digital_ldo_top_VIA4 $T=100850 21220 0 0 $X=100600 $Y=20990
X6049 2 digital_ldo_top_VIA4 $T=100850 25300 0 0 $X=100600 $Y=25070
X6050 2 digital_ldo_top_VIA4 $T=100850 29380 0 0 $X=100600 $Y=29150
X6051 2 digital_ldo_top_VIA4 $T=100850 33460 0 0 $X=100600 $Y=33230
X6052 2 digital_ldo_top_VIA4 $T=100850 37540 0 0 $X=100600 $Y=37310
X6053 2 digital_ldo_top_VIA4 $T=100850 41620 0 0 $X=100600 $Y=41390
X6054 2 digital_ldo_top_VIA4 $T=100850 45700 0 0 $X=100600 $Y=45470
X6055 2 digital_ldo_top_VIA4 $T=100850 49780 0 0 $X=100600 $Y=49550
X6056 2 digital_ldo_top_VIA4 $T=100850 53860 0 0 $X=100600 $Y=53630
X6057 2 digital_ldo_top_VIA4 $T=100850 57940 0 0 $X=100600 $Y=57710
X6058 2 digital_ldo_top_VIA4 $T=100850 62020 0 0 $X=100600 $Y=61790
X6059 2 digital_ldo_top_VIA4 $T=100850 66100 0 0 $X=100600 $Y=65870
X6060 2 digital_ldo_top_VIA4 $T=100850 70180 0 0 $X=100600 $Y=69950
X6061 2 digital_ldo_top_VIA4 $T=100850 74260 0 0 $X=100600 $Y=74030
X6062 2 digital_ldo_top_VIA4 $T=100850 78340 0 0 $X=100600 $Y=78110
X6063 2 digital_ldo_top_VIA4 $T=100850 82420 0 0 $X=100600 $Y=82190
X6064 2 digital_ldo_top_VIA4 $T=100850 86500 0 0 $X=100600 $Y=86270
X6065 2 digital_ldo_top_VIA4 $T=100850 90580 0 0 $X=100600 $Y=90350
X6066 2 digital_ldo_top_VIA4 $T=100850 94660 0 0 $X=100600 $Y=94430
X6067 2 digital_ldo_top_VIA4 $T=100850 98740 0 0 $X=100600 $Y=98510
X6068 2 digital_ldo_top_VIA4 $T=100850 102820 0 0 $X=100600 $Y=102590
X6069 2 digital_ldo_top_VIA4 $T=100850 106900 0 0 $X=100600 $Y=106670
X6070 2 digital_ldo_top_VIA4 $T=100850 110980 0 0 $X=100600 $Y=110750
X6071 2 digital_ldo_top_VIA4 $T=100850 115060 0 0 $X=100600 $Y=114830
X6072 2 digital_ldo_top_VIA4 $T=100850 119140 0 0 $X=100600 $Y=118910
X6073 2 digital_ldo_top_VIA4 $T=100850 123220 0 0 $X=100600 $Y=122990
X6074 2 digital_ldo_top_VIA4 $T=100850 127300 0 0 $X=100600 $Y=127070
X6075 3 digital_ldo_top_VIA4 $T=103150 11700 0 0 $X=102900 $Y=11470
X6076 3 digital_ldo_top_VIA4 $T=103150 15780 0 0 $X=102900 $Y=15550
X6077 3 digital_ldo_top_VIA4 $T=103150 19860 0 0 $X=102900 $Y=19630
X6078 3 digital_ldo_top_VIA4 $T=103150 23940 0 0 $X=102900 $Y=23710
X6079 3 digital_ldo_top_VIA4 $T=103150 32100 0 0 $X=102900 $Y=31870
X6080 3 digital_ldo_top_VIA4 $T=103150 85140 0 0 $X=102900 $Y=84910
X6081 3 digital_ldo_top_VIA4 $T=103150 89220 0 0 $X=102900 $Y=88990
X6082 3 digital_ldo_top_VIA4 $T=103150 93300 0 0 $X=102900 $Y=93070
X6083 3 digital_ldo_top_VIA4 $T=103150 97380 0 0 $X=102900 $Y=97150
X6084 3 digital_ldo_top_VIA4 $T=103150 101460 0 0 $X=102900 $Y=101230
X6085 3 digital_ldo_top_VIA4 $T=103150 105540 0 0 $X=102900 $Y=105310
X6086 3 digital_ldo_top_VIA4 $T=103150 109620 0 0 $X=102900 $Y=109390
X6087 3 digital_ldo_top_VIA4 $T=103150 113700 0 0 $X=102900 $Y=113470
X6088 3 digital_ldo_top_VIA4 $T=103150 117780 0 0 $X=102900 $Y=117550
X6089 3 digital_ldo_top_VIA4 $T=103150 121860 0 0 $X=102900 $Y=121630
X6090 3 digital_ldo_top_VIA4 $T=103150 125940 0 0 $X=102900 $Y=125710
X6091 2 digital_ldo_top_VIA4 $T=104530 13060 0 0 $X=104280 $Y=12830
X6092 2 digital_ldo_top_VIA4 $T=104530 17140 0 0 $X=104280 $Y=16910
X6093 2 digital_ldo_top_VIA4 $T=104530 21220 0 0 $X=104280 $Y=20990
X6094 2 digital_ldo_top_VIA4 $T=104530 25300 0 0 $X=104280 $Y=25070
X6095 2 digital_ldo_top_VIA4 $T=104530 86500 0 0 $X=104280 $Y=86270
X6096 2 digital_ldo_top_VIA4 $T=104530 90580 0 0 $X=104280 $Y=90350
X6097 2 digital_ldo_top_VIA4 $T=104530 94660 0 0 $X=104280 $Y=94430
X6098 2 digital_ldo_top_VIA4 $T=104530 98740 0 0 $X=104280 $Y=98510
X6099 2 digital_ldo_top_VIA4 $T=104530 102820 0 0 $X=104280 $Y=102590
X6100 2 digital_ldo_top_VIA4 $T=104530 106900 0 0 $X=104280 $Y=106670
X6101 2 digital_ldo_top_VIA4 $T=104530 110980 0 0 $X=104280 $Y=110750
X6102 2 digital_ldo_top_VIA4 $T=104530 115060 0 0 $X=104280 $Y=114830
X6103 2 digital_ldo_top_VIA4 $T=104530 119140 0 0 $X=104280 $Y=118910
X6104 2 digital_ldo_top_VIA4 $T=104530 123220 0 0 $X=104280 $Y=122990
X6105 2 digital_ldo_top_VIA4 $T=104530 127300 0 0 $X=104280 $Y=127070
X6106 3 digital_ldo_top_VIA4 $T=106830 11700 0 0 $X=106580 $Y=11470
X6107 3 digital_ldo_top_VIA4 $T=106830 15780 0 0 $X=106580 $Y=15550
X6108 3 digital_ldo_top_VIA4 $T=106830 19860 0 0 $X=106580 $Y=19630
X6109 3 digital_ldo_top_VIA4 $T=106830 23940 0 0 $X=106580 $Y=23710
X6110 3 digital_ldo_top_VIA4 $T=106830 32100 0 0 $X=106580 $Y=31870
X6111 3 digital_ldo_top_VIA4 $T=106830 85140 0 0 $X=106580 $Y=84910
X6112 3 digital_ldo_top_VIA4 $T=106830 89220 0 0 $X=106580 $Y=88990
X6113 3 digital_ldo_top_VIA4 $T=106830 93300 0 0 $X=106580 $Y=93070
X6114 3 digital_ldo_top_VIA4 $T=106830 97380 0 0 $X=106580 $Y=97150
X6115 3 digital_ldo_top_VIA4 $T=106830 101460 0 0 $X=106580 $Y=101230
X6116 3 digital_ldo_top_VIA4 $T=106830 105540 0 0 $X=106580 $Y=105310
X6117 3 digital_ldo_top_VIA4 $T=106830 109620 0 0 $X=106580 $Y=109390
X6118 3 digital_ldo_top_VIA4 $T=106830 113700 0 0 $X=106580 $Y=113470
X6119 3 digital_ldo_top_VIA4 $T=106830 117780 0 0 $X=106580 $Y=117550
X6120 3 digital_ldo_top_VIA4 $T=106830 121860 0 0 $X=106580 $Y=121630
X6121 3 digital_ldo_top_VIA4 $T=106830 125940 0 0 $X=106580 $Y=125710
X6122 2 digital_ldo_top_VIA4 $T=108210 13060 0 0 $X=107960 $Y=12830
X6123 2 digital_ldo_top_VIA4 $T=108210 17140 0 0 $X=107960 $Y=16910
X6124 2 digital_ldo_top_VIA4 $T=108210 21220 0 0 $X=107960 $Y=20990
X6125 2 digital_ldo_top_VIA4 $T=108210 25300 0 0 $X=107960 $Y=25070
X6126 2 digital_ldo_top_VIA4 $T=108210 86500 0 0 $X=107960 $Y=86270
X6127 2 digital_ldo_top_VIA4 $T=108210 90580 0 0 $X=107960 $Y=90350
X6128 2 digital_ldo_top_VIA4 $T=108210 94660 0 0 $X=107960 $Y=94430
X6129 2 digital_ldo_top_VIA4 $T=108210 98740 0 0 $X=107960 $Y=98510
X6130 2 digital_ldo_top_VIA4 $T=108210 102820 0 0 $X=107960 $Y=102590
X6131 2 digital_ldo_top_VIA4 $T=108210 106900 0 0 $X=107960 $Y=106670
X6132 2 digital_ldo_top_VIA4 $T=108210 110980 0 0 $X=107960 $Y=110750
X6133 2 digital_ldo_top_VIA4 $T=108210 115060 0 0 $X=107960 $Y=114830
X6134 2 digital_ldo_top_VIA4 $T=108210 119140 0 0 $X=107960 $Y=118910
X6135 2 digital_ldo_top_VIA4 $T=108210 123220 0 0 $X=107960 $Y=122990
X6136 2 digital_ldo_top_VIA4 $T=108210 127300 0 0 $X=107960 $Y=127070
X6137 3 digital_ldo_top_VIA4 $T=110510 11700 0 0 $X=110260 $Y=11470
X6138 3 digital_ldo_top_VIA4 $T=110510 15780 0 0 $X=110260 $Y=15550
X6139 3 digital_ldo_top_VIA4 $T=110510 19860 0 0 $X=110260 $Y=19630
X6140 3 digital_ldo_top_VIA4 $T=110510 23940 0 0 $X=110260 $Y=23710
X6141 3 digital_ldo_top_VIA4 $T=110510 32100 0 0 $X=110260 $Y=31870
X6142 3 digital_ldo_top_VIA4 $T=110510 85140 0 0 $X=110260 $Y=84910
X6143 3 digital_ldo_top_VIA4 $T=110510 89220 0 0 $X=110260 $Y=88990
X6144 3 digital_ldo_top_VIA4 $T=110510 93300 0 0 $X=110260 $Y=93070
X6145 3 digital_ldo_top_VIA4 $T=110510 97380 0 0 $X=110260 $Y=97150
X6146 3 digital_ldo_top_VIA4 $T=110510 101460 0 0 $X=110260 $Y=101230
X6147 3 digital_ldo_top_VIA4 $T=110510 105540 0 0 $X=110260 $Y=105310
X6148 3 digital_ldo_top_VIA4 $T=110510 109620 0 0 $X=110260 $Y=109390
X6149 3 digital_ldo_top_VIA4 $T=110510 113700 0 0 $X=110260 $Y=113470
X6150 3 digital_ldo_top_VIA4 $T=110510 117780 0 0 $X=110260 $Y=117550
X6151 3 digital_ldo_top_VIA4 $T=110510 121860 0 0 $X=110260 $Y=121630
X6152 3 digital_ldo_top_VIA4 $T=110510 125940 0 0 $X=110260 $Y=125710
X6153 2 digital_ldo_top_VIA4 $T=111890 13060 0 0 $X=111640 $Y=12830
X6154 2 digital_ldo_top_VIA4 $T=111890 17140 0 0 $X=111640 $Y=16910
X6155 2 digital_ldo_top_VIA4 $T=111890 21220 0 0 $X=111640 $Y=20990
X6156 2 digital_ldo_top_VIA4 $T=111890 25300 0 0 $X=111640 $Y=25070
X6157 2 digital_ldo_top_VIA4 $T=111890 86500 0 0 $X=111640 $Y=86270
X6158 2 digital_ldo_top_VIA4 $T=111890 90580 0 0 $X=111640 $Y=90350
X6159 2 digital_ldo_top_VIA4 $T=111890 94660 0 0 $X=111640 $Y=94430
X6160 2 digital_ldo_top_VIA4 $T=111890 98740 0 0 $X=111640 $Y=98510
X6161 2 digital_ldo_top_VIA4 $T=111890 102820 0 0 $X=111640 $Y=102590
X6162 2 digital_ldo_top_VIA4 $T=111890 106900 0 0 $X=111640 $Y=106670
X6163 2 digital_ldo_top_VIA4 $T=111890 110980 0 0 $X=111640 $Y=110750
X6164 2 digital_ldo_top_VIA4 $T=111890 115060 0 0 $X=111640 $Y=114830
X6165 2 digital_ldo_top_VIA4 $T=111890 119140 0 0 $X=111640 $Y=118910
X6166 2 digital_ldo_top_VIA4 $T=111890 123220 0 0 $X=111640 $Y=122990
X6167 2 digital_ldo_top_VIA4 $T=111890 127300 0 0 $X=111640 $Y=127070
X6168 3 digital_ldo_top_VIA4 $T=114190 11700 0 0 $X=113940 $Y=11470
X6169 3 digital_ldo_top_VIA4 $T=114190 15780 0 0 $X=113940 $Y=15550
X6170 3 digital_ldo_top_VIA4 $T=114190 19860 0 0 $X=113940 $Y=19630
X6171 3 digital_ldo_top_VIA4 $T=114190 23940 0 0 $X=113940 $Y=23710
X6172 3 digital_ldo_top_VIA4 $T=114190 32100 0 0 $X=113940 $Y=31870
X6173 3 digital_ldo_top_VIA4 $T=114190 85140 0 0 $X=113940 $Y=84910
X6174 3 digital_ldo_top_VIA4 $T=114190 89220 0 0 $X=113940 $Y=88990
X6175 3 digital_ldo_top_VIA4 $T=114190 93300 0 0 $X=113940 $Y=93070
X6176 3 digital_ldo_top_VIA4 $T=114190 97380 0 0 $X=113940 $Y=97150
X6177 3 digital_ldo_top_VIA4 $T=114190 101460 0 0 $X=113940 $Y=101230
X6178 3 digital_ldo_top_VIA4 $T=114190 105540 0 0 $X=113940 $Y=105310
X6179 3 digital_ldo_top_VIA4 $T=114190 109620 0 0 $X=113940 $Y=109390
X6180 3 digital_ldo_top_VIA4 $T=114190 113700 0 0 $X=113940 $Y=113470
X6181 3 digital_ldo_top_VIA4 $T=114190 117780 0 0 $X=113940 $Y=117550
X6182 3 digital_ldo_top_VIA4 $T=114190 121860 0 0 $X=113940 $Y=121630
X6183 3 digital_ldo_top_VIA4 $T=114190 125940 0 0 $X=113940 $Y=125710
X6184 2 digital_ldo_top_VIA4 $T=115570 13060 0 0 $X=115320 $Y=12830
X6185 2 digital_ldo_top_VIA4 $T=115570 17140 0 0 $X=115320 $Y=16910
X6186 2 digital_ldo_top_VIA4 $T=115570 94660 0 0 $X=115320 $Y=94430
X6187 2 digital_ldo_top_VIA4 $T=115570 98740 0 0 $X=115320 $Y=98510
X6188 2 digital_ldo_top_VIA4 $T=115570 102820 0 0 $X=115320 $Y=102590
X6189 2 digital_ldo_top_VIA4 $T=115570 106900 0 0 $X=115320 $Y=106670
X6190 2 digital_ldo_top_VIA4 $T=115570 110980 0 0 $X=115320 $Y=110750
X6191 2 digital_ldo_top_VIA4 $T=115570 115060 0 0 $X=115320 $Y=114830
X6192 2 digital_ldo_top_VIA4 $T=115570 119140 0 0 $X=115320 $Y=118910
X6193 2 digital_ldo_top_VIA4 $T=115570 123220 0 0 $X=115320 $Y=122990
X6194 2 digital_ldo_top_VIA4 $T=115570 127300 0 0 $X=115320 $Y=127070
X6195 3 digital_ldo_top_VIA4 $T=117870 11700 0 0 $X=117620 $Y=11470
X6196 3 digital_ldo_top_VIA4 $T=117870 15780 0 0 $X=117620 $Y=15550
X6197 3 digital_ldo_top_VIA4 $T=117870 19860 0 0 $X=117620 $Y=19630
X6198 3 digital_ldo_top_VIA4 $T=117870 23940 0 0 $X=117620 $Y=23710
X6199 3 digital_ldo_top_VIA4 $T=117870 32100 0 0 $X=117620 $Y=31870
X6200 3 digital_ldo_top_VIA4 $T=117870 85140 0 0 $X=117620 $Y=84910
X6201 3 digital_ldo_top_VIA4 $T=117870 89220 0 0 $X=117620 $Y=88990
X6202 3 digital_ldo_top_VIA4 $T=117870 93300 0 0 $X=117620 $Y=93070
X6203 3 digital_ldo_top_VIA4 $T=117870 97380 0 0 $X=117620 $Y=97150
X6204 3 digital_ldo_top_VIA4 $T=117870 101460 0 0 $X=117620 $Y=101230
X6205 3 digital_ldo_top_VIA4 $T=117870 105540 0 0 $X=117620 $Y=105310
X6206 3 digital_ldo_top_VIA4 $T=117870 109620 0 0 $X=117620 $Y=109390
X6207 3 digital_ldo_top_VIA4 $T=117870 113700 0 0 $X=117620 $Y=113470
X6208 3 digital_ldo_top_VIA4 $T=117870 117780 0 0 $X=117620 $Y=117550
X6209 3 digital_ldo_top_VIA4 $T=117870 121860 0 0 $X=117620 $Y=121630
X6210 3 digital_ldo_top_VIA4 $T=117870 125940 0 0 $X=117620 $Y=125710
X6211 2 digital_ldo_top_VIA4 $T=119250 13060 0 0 $X=119000 $Y=12830
X6212 2 digital_ldo_top_VIA4 $T=119250 17140 0 0 $X=119000 $Y=16910
X6213 2 digital_ldo_top_VIA4 $T=119250 21220 0 0 $X=119000 $Y=20990
X6214 2 digital_ldo_top_VIA4 $T=119250 25300 0 0 $X=119000 $Y=25070
X6215 2 digital_ldo_top_VIA4 $T=119250 94660 0 0 $X=119000 $Y=94430
X6216 2 digital_ldo_top_VIA4 $T=119250 98740 0 0 $X=119000 $Y=98510
X6217 2 digital_ldo_top_VIA4 $T=119250 102820 0 0 $X=119000 $Y=102590
X6218 2 digital_ldo_top_VIA4 $T=119250 106900 0 0 $X=119000 $Y=106670
X6219 2 digital_ldo_top_VIA4 $T=119250 110980 0 0 $X=119000 $Y=110750
X6220 2 digital_ldo_top_VIA4 $T=119250 115060 0 0 $X=119000 $Y=114830
X6221 2 digital_ldo_top_VIA4 $T=119250 119140 0 0 $X=119000 $Y=118910
X6222 2 digital_ldo_top_VIA4 $T=119250 123220 0 0 $X=119000 $Y=122990
X6223 2 digital_ldo_top_VIA4 $T=119250 127300 0 0 $X=119000 $Y=127070
X6224 3 digital_ldo_top_VIA4 $T=121550 11700 0 0 $X=121300 $Y=11470
X6225 3 digital_ldo_top_VIA4 $T=121550 15780 0 0 $X=121300 $Y=15550
X6226 3 digital_ldo_top_VIA4 $T=121550 19860 0 0 $X=121300 $Y=19630
X6227 3 digital_ldo_top_VIA4 $T=121550 23940 0 0 $X=121300 $Y=23710
X6228 3 digital_ldo_top_VIA4 $T=121550 32100 0 0 $X=121300 $Y=31870
X6229 3 digital_ldo_top_VIA4 $T=121550 85140 0 0 $X=121300 $Y=84910
X6230 3 digital_ldo_top_VIA4 $T=121550 89220 0 0 $X=121300 $Y=88990
X6231 3 digital_ldo_top_VIA4 $T=121550 93300 0 0 $X=121300 $Y=93070
X6232 3 digital_ldo_top_VIA4 $T=121550 97380 0 0 $X=121300 $Y=97150
X6233 3 digital_ldo_top_VIA4 $T=121550 101460 0 0 $X=121300 $Y=101230
X6234 3 digital_ldo_top_VIA4 $T=121550 105540 0 0 $X=121300 $Y=105310
X6235 3 digital_ldo_top_VIA4 $T=121550 109620 0 0 $X=121300 $Y=109390
X6236 3 digital_ldo_top_VIA4 $T=121550 113700 0 0 $X=121300 $Y=113470
X6237 3 digital_ldo_top_VIA4 $T=121550 117780 0 0 $X=121300 $Y=117550
X6238 3 digital_ldo_top_VIA4 $T=121550 121860 0 0 $X=121300 $Y=121630
X6239 3 digital_ldo_top_VIA4 $T=121550 125940 0 0 $X=121300 $Y=125710
X6240 2 digital_ldo_top_VIA4 $T=122930 13060 0 0 $X=122680 $Y=12830
X6241 2 digital_ldo_top_VIA4 $T=122930 17140 0 0 $X=122680 $Y=16910
X6242 2 digital_ldo_top_VIA4 $T=122930 21220 0 0 $X=122680 $Y=20990
X6243 2 digital_ldo_top_VIA4 $T=122930 25300 0 0 $X=122680 $Y=25070
X6244 2 digital_ldo_top_VIA4 $T=122930 86500 0 0 $X=122680 $Y=86270
X6245 2 digital_ldo_top_VIA4 $T=122930 90580 0 0 $X=122680 $Y=90350
X6246 2 digital_ldo_top_VIA4 $T=122930 94660 0 0 $X=122680 $Y=94430
X6247 2 digital_ldo_top_VIA4 $T=122930 98740 0 0 $X=122680 $Y=98510
X6248 2 digital_ldo_top_VIA4 $T=122930 102820 0 0 $X=122680 $Y=102590
X6249 2 digital_ldo_top_VIA4 $T=122930 106900 0 0 $X=122680 $Y=106670
X6250 2 digital_ldo_top_VIA4 $T=122930 110980 0 0 $X=122680 $Y=110750
X6251 2 digital_ldo_top_VIA4 $T=122930 115060 0 0 $X=122680 $Y=114830
X6252 2 digital_ldo_top_VIA4 $T=122930 119140 0 0 $X=122680 $Y=118910
X6253 2 digital_ldo_top_VIA4 $T=122930 123220 0 0 $X=122680 $Y=122990
X6254 2 digital_ldo_top_VIA4 $T=122930 127300 0 0 $X=122680 $Y=127070
X6255 3 digital_ldo_top_VIA4 $T=125230 11700 0 0 $X=124980 $Y=11470
X6256 3 digital_ldo_top_VIA4 $T=125230 15780 0 0 $X=124980 $Y=15550
X6257 3 digital_ldo_top_VIA4 $T=125230 93300 0 0 $X=124980 $Y=93070
X6258 3 digital_ldo_top_VIA4 $T=125230 97380 0 0 $X=124980 $Y=97150
X6259 3 digital_ldo_top_VIA4 $T=125230 101460 0 0 $X=124980 $Y=101230
X6260 3 digital_ldo_top_VIA4 $T=125230 105540 0 0 $X=124980 $Y=105310
X6261 3 digital_ldo_top_VIA4 $T=125230 109620 0 0 $X=124980 $Y=109390
X6262 3 digital_ldo_top_VIA4 $T=125230 113700 0 0 $X=124980 $Y=113470
X6263 3 digital_ldo_top_VIA4 $T=125230 117780 0 0 $X=124980 $Y=117550
X6264 3 digital_ldo_top_VIA4 $T=125230 121860 0 0 $X=124980 $Y=121630
X6265 3 digital_ldo_top_VIA4 $T=125230 125940 0 0 $X=124980 $Y=125710
X6266 2 digital_ldo_top_VIA4 $T=126610 13060 0 0 $X=126360 $Y=12830
X6267 2 digital_ldo_top_VIA4 $T=126610 17140 0 0 $X=126360 $Y=16910
X6268 2 digital_ldo_top_VIA4 $T=126610 21220 0 0 $X=126360 $Y=20990
X6269 2 digital_ldo_top_VIA4 $T=126610 25300 0 0 $X=126360 $Y=25070
X6270 2 digital_ldo_top_VIA4 $T=126610 94660 0 0 $X=126360 $Y=94430
X6271 2 digital_ldo_top_VIA4 $T=126610 98740 0 0 $X=126360 $Y=98510
X6272 2 digital_ldo_top_VIA4 $T=126610 102820 0 0 $X=126360 $Y=102590
X6273 2 digital_ldo_top_VIA4 $T=126610 106900 0 0 $X=126360 $Y=106670
X6274 2 digital_ldo_top_VIA4 $T=126610 110980 0 0 $X=126360 $Y=110750
X6275 2 digital_ldo_top_VIA4 $T=126610 115060 0 0 $X=126360 $Y=114830
X6276 2 digital_ldo_top_VIA4 $T=126610 119140 0 0 $X=126360 $Y=118910
X6277 2 digital_ldo_top_VIA4 $T=126610 123220 0 0 $X=126360 $Y=122990
X6278 2 digital_ldo_top_VIA4 $T=126610 127300 0 0 $X=126360 $Y=127070
X6279 3 digital_ldo_top_VIA4 $T=128910 11700 0 0 $X=128660 $Y=11470
X6280 3 digital_ldo_top_VIA4 $T=128910 15780 0 0 $X=128660 $Y=15550
X6281 3 digital_ldo_top_VIA4 $T=128910 19860 0 0 $X=128660 $Y=19630
X6282 3 digital_ldo_top_VIA4 $T=128910 23940 0 0 $X=128660 $Y=23710
X6283 3 digital_ldo_top_VIA4 $T=128910 32100 0 0 $X=128660 $Y=31870
X6284 3 digital_ldo_top_VIA4 $T=128910 85140 0 0 $X=128660 $Y=84910
X6285 3 digital_ldo_top_VIA4 $T=128910 89220 0 0 $X=128660 $Y=88990
X6286 3 digital_ldo_top_VIA4 $T=128910 93300 0 0 $X=128660 $Y=93070
X6287 3 digital_ldo_top_VIA4 $T=128910 97380 0 0 $X=128660 $Y=97150
X6288 3 digital_ldo_top_VIA4 $T=128910 101460 0 0 $X=128660 $Y=101230
X6289 3 digital_ldo_top_VIA4 $T=128910 105540 0 0 $X=128660 $Y=105310
X6290 3 digital_ldo_top_VIA4 $T=128910 109620 0 0 $X=128660 $Y=109390
X6291 3 digital_ldo_top_VIA4 $T=128910 113700 0 0 $X=128660 $Y=113470
X6292 3 digital_ldo_top_VIA4 $T=128910 117780 0 0 $X=128660 $Y=117550
X6293 3 digital_ldo_top_VIA4 $T=128910 121860 0 0 $X=128660 $Y=121630
X6294 3 digital_ldo_top_VIA4 $T=128910 125940 0 0 $X=128660 $Y=125710
X6295 2 digital_ldo_top_VIA4 $T=130290 13060 0 0 $X=130040 $Y=12830
X6296 2 digital_ldo_top_VIA4 $T=130290 17140 0 0 $X=130040 $Y=16910
X6297 2 digital_ldo_top_VIA4 $T=130290 21220 0 0 $X=130040 $Y=20990
X6298 2 digital_ldo_top_VIA4 $T=130290 25300 0 0 $X=130040 $Y=25070
X6299 2 digital_ldo_top_VIA4 $T=130290 94660 0 0 $X=130040 $Y=94430
X6300 2 digital_ldo_top_VIA4 $T=130290 98740 0 0 $X=130040 $Y=98510
X6301 2 digital_ldo_top_VIA4 $T=130290 102820 0 0 $X=130040 $Y=102590
X6302 2 digital_ldo_top_VIA4 $T=130290 106900 0 0 $X=130040 $Y=106670
X6303 2 digital_ldo_top_VIA4 $T=130290 110980 0 0 $X=130040 $Y=110750
X6304 2 digital_ldo_top_VIA4 $T=130290 115060 0 0 $X=130040 $Y=114830
X6305 2 digital_ldo_top_VIA4 $T=130290 119140 0 0 $X=130040 $Y=118910
X6306 2 digital_ldo_top_VIA4 $T=130290 123220 0 0 $X=130040 $Y=122990
X6307 2 digital_ldo_top_VIA4 $T=130290 127300 0 0 $X=130040 $Y=127070
X6308 3 digital_ldo_top_VIA4 $T=132590 11700 0 0 $X=132340 $Y=11470
X6309 3 digital_ldo_top_VIA4 $T=132590 15780 0 0 $X=132340 $Y=15550
X6310 3 digital_ldo_top_VIA4 $T=132590 19860 0 0 $X=132340 $Y=19630
X6311 3 digital_ldo_top_VIA4 $T=132590 23940 0 0 $X=132340 $Y=23710
X6312 3 digital_ldo_top_VIA4 $T=132590 32100 0 0 $X=132340 $Y=31870
X6313 3 digital_ldo_top_VIA4 $T=132590 85140 0 0 $X=132340 $Y=84910
X6314 3 digital_ldo_top_VIA4 $T=132590 89220 0 0 $X=132340 $Y=88990
X6315 3 digital_ldo_top_VIA4 $T=132590 93300 0 0 $X=132340 $Y=93070
X6316 3 digital_ldo_top_VIA4 $T=132590 97380 0 0 $X=132340 $Y=97150
X6317 3 digital_ldo_top_VIA4 $T=132590 101460 0 0 $X=132340 $Y=101230
X6318 3 digital_ldo_top_VIA4 $T=132590 105540 0 0 $X=132340 $Y=105310
X6319 3 digital_ldo_top_VIA4 $T=132590 109620 0 0 $X=132340 $Y=109390
X6320 3 digital_ldo_top_VIA4 $T=132590 113700 0 0 $X=132340 $Y=113470
X6321 3 digital_ldo_top_VIA4 $T=132590 117780 0 0 $X=132340 $Y=117550
X6322 3 digital_ldo_top_VIA4 $T=132590 121860 0 0 $X=132340 $Y=121630
X6323 3 digital_ldo_top_VIA4 $T=132590 125940 0 0 $X=132340 $Y=125710
X6324 2 digital_ldo_top_VIA4 $T=133970 13060 0 0 $X=133720 $Y=12830
X6325 2 digital_ldo_top_VIA4 $T=133970 17140 0 0 $X=133720 $Y=16910
X6326 2 digital_ldo_top_VIA4 $T=133970 21220 0 0 $X=133720 $Y=20990
X6327 2 digital_ldo_top_VIA4 $T=133970 25300 0 0 $X=133720 $Y=25070
X6328 2 digital_ldo_top_VIA4 $T=133970 86500 0 0 $X=133720 $Y=86270
X6329 2 digital_ldo_top_VIA4 $T=133970 90580 0 0 $X=133720 $Y=90350
X6330 2 digital_ldo_top_VIA4 $T=133970 94660 0 0 $X=133720 $Y=94430
X6331 2 digital_ldo_top_VIA4 $T=133970 98740 0 0 $X=133720 $Y=98510
X6332 2 digital_ldo_top_VIA4 $T=133970 102820 0 0 $X=133720 $Y=102590
X6333 2 digital_ldo_top_VIA4 $T=133970 106900 0 0 $X=133720 $Y=106670
X6334 2 digital_ldo_top_VIA4 $T=133970 110980 0 0 $X=133720 $Y=110750
X6335 2 digital_ldo_top_VIA4 $T=133970 115060 0 0 $X=133720 $Y=114830
X6336 2 digital_ldo_top_VIA4 $T=133970 119140 0 0 $X=133720 $Y=118910
X6337 2 digital_ldo_top_VIA4 $T=133970 123220 0 0 $X=133720 $Y=122990
X6338 2 digital_ldo_top_VIA4 $T=133970 127300 0 0 $X=133720 $Y=127070
X6339 3 digital_ldo_top_VIA4 $T=136270 11700 0 0 $X=136020 $Y=11470
X6340 3 digital_ldo_top_VIA4 $T=136270 15780 0 0 $X=136020 $Y=15550
X6341 3 digital_ldo_top_VIA4 $T=136270 93300 0 0 $X=136020 $Y=93070
X6342 3 digital_ldo_top_VIA4 $T=136270 97380 0 0 $X=136020 $Y=97150
X6343 3 digital_ldo_top_VIA4 $T=136270 101460 0 0 $X=136020 $Y=101230
X6344 3 digital_ldo_top_VIA4 $T=136270 105540 0 0 $X=136020 $Y=105310
X6345 3 digital_ldo_top_VIA4 $T=136270 109620 0 0 $X=136020 $Y=109390
X6346 3 digital_ldo_top_VIA4 $T=136270 113700 0 0 $X=136020 $Y=113470
X6347 3 digital_ldo_top_VIA4 $T=136270 117780 0 0 $X=136020 $Y=117550
X6348 3 digital_ldo_top_VIA4 $T=136270 121860 0 0 $X=136020 $Y=121630
X6349 3 digital_ldo_top_VIA4 $T=136270 125940 0 0 $X=136020 $Y=125710
X6350 2 digital_ldo_top_VIA4 $T=137650 13060 0 0 $X=137400 $Y=12830
X6351 2 digital_ldo_top_VIA4 $T=137650 17140 0 0 $X=137400 $Y=16910
X6352 2 digital_ldo_top_VIA4 $T=137650 21220 0 0 $X=137400 $Y=20990
X6353 2 digital_ldo_top_VIA4 $T=137650 25300 0 0 $X=137400 $Y=25070
X6354 2 digital_ldo_top_VIA4 $T=137650 94660 0 0 $X=137400 $Y=94430
X6355 2 digital_ldo_top_VIA4 $T=137650 98740 0 0 $X=137400 $Y=98510
X6356 2 digital_ldo_top_VIA4 $T=137650 102820 0 0 $X=137400 $Y=102590
X6357 2 digital_ldo_top_VIA4 $T=137650 106900 0 0 $X=137400 $Y=106670
X6358 2 digital_ldo_top_VIA4 $T=137650 110980 0 0 $X=137400 $Y=110750
X6359 2 digital_ldo_top_VIA4 $T=137650 115060 0 0 $X=137400 $Y=114830
X6360 2 digital_ldo_top_VIA4 $T=137650 119140 0 0 $X=137400 $Y=118910
X6361 2 digital_ldo_top_VIA4 $T=137650 123220 0 0 $X=137400 $Y=122990
X6362 2 digital_ldo_top_VIA4 $T=137650 127300 0 0 $X=137400 $Y=127070
X6363 3 digital_ldo_top_VIA4 $T=139950 11700 0 0 $X=139700 $Y=11470
X6364 3 digital_ldo_top_VIA4 $T=139950 15780 0 0 $X=139700 $Y=15550
X6365 3 digital_ldo_top_VIA4 $T=139950 85140 0 0 $X=139700 $Y=84910
X6366 3 digital_ldo_top_VIA4 $T=139950 89220 0 0 $X=139700 $Y=88990
X6367 3 digital_ldo_top_VIA4 $T=139950 93300 0 0 $X=139700 $Y=93070
X6368 3 digital_ldo_top_VIA4 $T=139950 97380 0 0 $X=139700 $Y=97150
X6369 3 digital_ldo_top_VIA4 $T=139950 101460 0 0 $X=139700 $Y=101230
X6370 3 digital_ldo_top_VIA4 $T=139950 105540 0 0 $X=139700 $Y=105310
X6371 3 digital_ldo_top_VIA4 $T=139950 109620 0 0 $X=139700 $Y=109390
X6372 3 digital_ldo_top_VIA4 $T=139950 113700 0 0 $X=139700 $Y=113470
X6373 3 digital_ldo_top_VIA4 $T=139950 117780 0 0 $X=139700 $Y=117550
X6374 3 digital_ldo_top_VIA4 $T=139950 121860 0 0 $X=139700 $Y=121630
X6375 3 digital_ldo_top_VIA4 $T=139950 125940 0 0 $X=139700 $Y=125710
X6376 2 digital_ldo_top_VIA4 $T=141330 13060 0 0 $X=141080 $Y=12830
X6377 2 digital_ldo_top_VIA4 $T=141330 17140 0 0 $X=141080 $Y=16910
X6378 2 digital_ldo_top_VIA4 $T=141330 21220 0 0 $X=141080 $Y=20990
X6379 2 digital_ldo_top_VIA4 $T=141330 25300 0 0 $X=141080 $Y=25070
X6380 2 digital_ldo_top_VIA4 $T=141330 94660 0 0 $X=141080 $Y=94430
X6381 2 digital_ldo_top_VIA4 $T=141330 98740 0 0 $X=141080 $Y=98510
X6382 2 digital_ldo_top_VIA4 $T=141330 102820 0 0 $X=141080 $Y=102590
X6383 2 digital_ldo_top_VIA4 $T=141330 106900 0 0 $X=141080 $Y=106670
X6384 2 digital_ldo_top_VIA4 $T=141330 110980 0 0 $X=141080 $Y=110750
X6385 2 digital_ldo_top_VIA4 $T=141330 115060 0 0 $X=141080 $Y=114830
X6386 2 digital_ldo_top_VIA4 $T=141330 119140 0 0 $X=141080 $Y=118910
X6387 2 digital_ldo_top_VIA4 $T=141330 123220 0 0 $X=141080 $Y=122990
X6388 2 digital_ldo_top_VIA4 $T=141330 127300 0 0 $X=141080 $Y=127070
X6389 3 digital_ldo_top_VIA4 $T=143630 11700 0 0 $X=143380 $Y=11470
X6390 3 digital_ldo_top_VIA4 $T=143630 15780 0 0 $X=143380 $Y=15550
X6391 3 digital_ldo_top_VIA4 $T=143630 85140 0 0 $X=143380 $Y=84910
X6392 3 digital_ldo_top_VIA4 $T=143630 89220 0 0 $X=143380 $Y=88990
X6393 3 digital_ldo_top_VIA4 $T=143630 93300 0 0 $X=143380 $Y=93070
X6394 3 digital_ldo_top_VIA4 $T=143630 97380 0 0 $X=143380 $Y=97150
X6395 3 digital_ldo_top_VIA4 $T=143630 101460 0 0 $X=143380 $Y=101230
X6396 3 digital_ldo_top_VIA4 $T=143630 105540 0 0 $X=143380 $Y=105310
X6397 3 digital_ldo_top_VIA4 $T=143630 109620 0 0 $X=143380 $Y=109390
X6398 3 digital_ldo_top_VIA4 $T=143630 113700 0 0 $X=143380 $Y=113470
X6399 3 digital_ldo_top_VIA4 $T=143630 117780 0 0 $X=143380 $Y=117550
X6400 3 digital_ldo_top_VIA4 $T=143630 121860 0 0 $X=143380 $Y=121630
X6401 3 digital_ldo_top_VIA4 $T=143630 125940 0 0 $X=143380 $Y=125710
X6402 2 digital_ldo_top_VIA4 $T=145010 13060 0 0 $X=144760 $Y=12830
X6403 2 digital_ldo_top_VIA4 $T=145010 17140 0 0 $X=144760 $Y=16910
X6404 2 digital_ldo_top_VIA4 $T=145010 21220 0 0 $X=144760 $Y=20990
X6405 2 digital_ldo_top_VIA4 $T=145010 25300 0 0 $X=144760 $Y=25070
X6406 2 digital_ldo_top_VIA4 $T=145010 86500 0 0 $X=144760 $Y=86270
X6407 2 digital_ldo_top_VIA4 $T=145010 90580 0 0 $X=144760 $Y=90350
X6408 2 digital_ldo_top_VIA4 $T=145010 94660 0 0 $X=144760 $Y=94430
X6409 2 digital_ldo_top_VIA4 $T=145010 98740 0 0 $X=144760 $Y=98510
X6410 2 digital_ldo_top_VIA4 $T=145010 102820 0 0 $X=144760 $Y=102590
X6411 2 digital_ldo_top_VIA4 $T=145010 106900 0 0 $X=144760 $Y=106670
X6412 2 digital_ldo_top_VIA4 $T=145010 110980 0 0 $X=144760 $Y=110750
X6413 2 digital_ldo_top_VIA4 $T=145010 115060 0 0 $X=144760 $Y=114830
X6414 2 digital_ldo_top_VIA4 $T=145010 119140 0 0 $X=144760 $Y=118910
X6415 2 digital_ldo_top_VIA4 $T=145010 123220 0 0 $X=144760 $Y=122990
X6416 2 digital_ldo_top_VIA4 $T=145010 127300 0 0 $X=144760 $Y=127070
X6417 3 digital_ldo_top_VIA4 $T=147310 11700 0 0 $X=147060 $Y=11470
X6418 3 digital_ldo_top_VIA4 $T=147310 15780 0 0 $X=147060 $Y=15550
X6419 3 digital_ldo_top_VIA4 $T=147310 93300 0 0 $X=147060 $Y=93070
X6420 3 digital_ldo_top_VIA4 $T=147310 97380 0 0 $X=147060 $Y=97150
X6421 3 digital_ldo_top_VIA4 $T=147310 101460 0 0 $X=147060 $Y=101230
X6422 3 digital_ldo_top_VIA4 $T=147310 105540 0 0 $X=147060 $Y=105310
X6423 3 digital_ldo_top_VIA4 $T=147310 109620 0 0 $X=147060 $Y=109390
X6424 3 digital_ldo_top_VIA4 $T=147310 113700 0 0 $X=147060 $Y=113470
X6425 3 digital_ldo_top_VIA4 $T=147310 117780 0 0 $X=147060 $Y=117550
X6426 3 digital_ldo_top_VIA4 $T=147310 121860 0 0 $X=147060 $Y=121630
X6427 3 digital_ldo_top_VIA4 $T=147310 125940 0 0 $X=147060 $Y=125710
X6428 2 digital_ldo_top_VIA4 $T=148690 13060 0 0 $X=148440 $Y=12830
X6429 2 digital_ldo_top_VIA4 $T=148690 17140 0 0 $X=148440 $Y=16910
X6430 2 digital_ldo_top_VIA4 $T=148690 21220 0 0 $X=148440 $Y=20990
X6431 2 digital_ldo_top_VIA4 $T=148690 25300 0 0 $X=148440 $Y=25070
X6432 2 digital_ldo_top_VIA4 $T=148690 94660 0 0 $X=148440 $Y=94430
X6433 2 digital_ldo_top_VIA4 $T=148690 98740 0 0 $X=148440 $Y=98510
X6434 2 digital_ldo_top_VIA4 $T=148690 102820 0 0 $X=148440 $Y=102590
X6435 2 digital_ldo_top_VIA4 $T=148690 106900 0 0 $X=148440 $Y=106670
X6436 2 digital_ldo_top_VIA4 $T=148690 110980 0 0 $X=148440 $Y=110750
X6437 2 digital_ldo_top_VIA4 $T=148690 115060 0 0 $X=148440 $Y=114830
X6438 2 digital_ldo_top_VIA4 $T=148690 119140 0 0 $X=148440 $Y=118910
X6439 2 digital_ldo_top_VIA4 $T=148690 123220 0 0 $X=148440 $Y=122990
X6440 2 digital_ldo_top_VIA4 $T=148690 127300 0 0 $X=148440 $Y=127070
X6441 3 digital_ldo_top_VIA4 $T=150990 11700 0 0 $X=150740 $Y=11470
X6442 3 digital_ldo_top_VIA4 $T=150990 15780 0 0 $X=150740 $Y=15550
X6443 3 digital_ldo_top_VIA4 $T=150990 85140 0 0 $X=150740 $Y=84910
X6444 3 digital_ldo_top_VIA4 $T=150990 89220 0 0 $X=150740 $Y=88990
X6445 3 digital_ldo_top_VIA4 $T=150990 93300 0 0 $X=150740 $Y=93070
X6446 3 digital_ldo_top_VIA4 $T=150990 97380 0 0 $X=150740 $Y=97150
X6447 3 digital_ldo_top_VIA4 $T=150990 101460 0 0 $X=150740 $Y=101230
X6448 3 digital_ldo_top_VIA4 $T=150990 105540 0 0 $X=150740 $Y=105310
X6449 3 digital_ldo_top_VIA4 $T=150990 109620 0 0 $X=150740 $Y=109390
X6450 3 digital_ldo_top_VIA4 $T=150990 113700 0 0 $X=150740 $Y=113470
X6451 3 digital_ldo_top_VIA4 $T=150990 117780 0 0 $X=150740 $Y=117550
X6452 3 digital_ldo_top_VIA4 $T=150990 121860 0 0 $X=150740 $Y=121630
X6453 3 digital_ldo_top_VIA4 $T=150990 125940 0 0 $X=150740 $Y=125710
X6454 2 digital_ldo_top_VIA4 $T=152370 13060 0 0 $X=152120 $Y=12830
X6455 2 digital_ldo_top_VIA4 $T=152370 17140 0 0 $X=152120 $Y=16910
X6456 2 digital_ldo_top_VIA4 $T=152370 21220 0 0 $X=152120 $Y=20990
X6457 2 digital_ldo_top_VIA4 $T=152370 25300 0 0 $X=152120 $Y=25070
X6458 2 digital_ldo_top_VIA4 $T=152370 94660 0 0 $X=152120 $Y=94430
X6459 2 digital_ldo_top_VIA4 $T=152370 98740 0 0 $X=152120 $Y=98510
X6460 2 digital_ldo_top_VIA4 $T=152370 102820 0 0 $X=152120 $Y=102590
X6461 2 digital_ldo_top_VIA4 $T=152370 106900 0 0 $X=152120 $Y=106670
X6462 2 digital_ldo_top_VIA4 $T=152370 110980 0 0 $X=152120 $Y=110750
X6463 2 digital_ldo_top_VIA4 $T=152370 115060 0 0 $X=152120 $Y=114830
X6464 2 digital_ldo_top_VIA4 $T=152370 119140 0 0 $X=152120 $Y=118910
X6465 2 digital_ldo_top_VIA4 $T=152370 123220 0 0 $X=152120 $Y=122990
X6466 2 digital_ldo_top_VIA4 $T=152370 127300 0 0 $X=152120 $Y=127070
X6467 3 digital_ldo_top_VIA4 $T=154670 11700 0 0 $X=154420 $Y=11470
X6468 3 digital_ldo_top_VIA4 $T=154670 15780 0 0 $X=154420 $Y=15550
X6469 3 digital_ldo_top_VIA4 $T=154670 85140 0 0 $X=154420 $Y=84910
X6470 3 digital_ldo_top_VIA4 $T=154670 89220 0 0 $X=154420 $Y=88990
X6471 3 digital_ldo_top_VIA4 $T=154670 93300 0 0 $X=154420 $Y=93070
X6472 3 digital_ldo_top_VIA4 $T=154670 97380 0 0 $X=154420 $Y=97150
X6473 3 digital_ldo_top_VIA4 $T=154670 101460 0 0 $X=154420 $Y=101230
X6474 3 digital_ldo_top_VIA4 $T=154670 105540 0 0 $X=154420 $Y=105310
X6475 3 digital_ldo_top_VIA4 $T=154670 109620 0 0 $X=154420 $Y=109390
X6476 3 digital_ldo_top_VIA4 $T=154670 113700 0 0 $X=154420 $Y=113470
X6477 3 digital_ldo_top_VIA4 $T=154670 117780 0 0 $X=154420 $Y=117550
X6478 3 digital_ldo_top_VIA4 $T=154670 121860 0 0 $X=154420 $Y=121630
X6479 3 digital_ldo_top_VIA4 $T=154670 125940 0 0 $X=154420 $Y=125710
X6480 2 digital_ldo_top_VIA4 $T=156050 13060 0 0 $X=155800 $Y=12830
X6481 2 digital_ldo_top_VIA4 $T=156050 17140 0 0 $X=155800 $Y=16910
X6482 2 digital_ldo_top_VIA4 $T=156050 21220 0 0 $X=155800 $Y=20990
X6483 2 digital_ldo_top_VIA4 $T=156050 25300 0 0 $X=155800 $Y=25070
X6484 2 digital_ldo_top_VIA4 $T=156050 86500 0 0 $X=155800 $Y=86270
X6485 2 digital_ldo_top_VIA4 $T=156050 90580 0 0 $X=155800 $Y=90350
X6486 2 digital_ldo_top_VIA4 $T=156050 94660 0 0 $X=155800 $Y=94430
X6487 2 digital_ldo_top_VIA4 $T=156050 98740 0 0 $X=155800 $Y=98510
X6488 2 digital_ldo_top_VIA4 $T=156050 102820 0 0 $X=155800 $Y=102590
X6489 2 digital_ldo_top_VIA4 $T=156050 106900 0 0 $X=155800 $Y=106670
X6490 2 digital_ldo_top_VIA4 $T=156050 110980 0 0 $X=155800 $Y=110750
X6491 2 digital_ldo_top_VIA4 $T=156050 115060 0 0 $X=155800 $Y=114830
X6492 2 digital_ldo_top_VIA4 $T=156050 119140 0 0 $X=155800 $Y=118910
X6493 2 digital_ldo_top_VIA4 $T=156050 123220 0 0 $X=155800 $Y=122990
X6494 2 digital_ldo_top_VIA4 $T=156050 127300 0 0 $X=155800 $Y=127070
X6495 3 digital_ldo_top_VIA4 $T=158350 11700 0 0 $X=158100 $Y=11470
X6496 3 digital_ldo_top_VIA4 $T=158350 15780 0 0 $X=158100 $Y=15550
X6497 3 digital_ldo_top_VIA4 $T=158350 93300 0 0 $X=158100 $Y=93070
X6498 3 digital_ldo_top_VIA4 $T=158350 97380 0 0 $X=158100 $Y=97150
X6499 3 digital_ldo_top_VIA4 $T=158350 101460 0 0 $X=158100 $Y=101230
X6500 3 digital_ldo_top_VIA4 $T=158350 105540 0 0 $X=158100 $Y=105310
X6501 3 digital_ldo_top_VIA4 $T=158350 109620 0 0 $X=158100 $Y=109390
X6502 3 digital_ldo_top_VIA4 $T=158350 113700 0 0 $X=158100 $Y=113470
X6503 3 digital_ldo_top_VIA4 $T=158350 117780 0 0 $X=158100 $Y=117550
X6504 3 digital_ldo_top_VIA4 $T=158350 121860 0 0 $X=158100 $Y=121630
X6505 3 digital_ldo_top_VIA4 $T=158350 125940 0 0 $X=158100 $Y=125710
X6506 2 digital_ldo_top_VIA4 $T=159730 13060 0 0 $X=159480 $Y=12830
X6507 2 digital_ldo_top_VIA4 $T=159730 17140 0 0 $X=159480 $Y=16910
X6508 2 digital_ldo_top_VIA4 $T=159730 21220 0 0 $X=159480 $Y=20990
X6509 2 digital_ldo_top_VIA4 $T=159730 25300 0 0 $X=159480 $Y=25070
X6510 2 digital_ldo_top_VIA4 $T=159730 94660 0 0 $X=159480 $Y=94430
X6511 2 digital_ldo_top_VIA4 $T=159730 98740 0 0 $X=159480 $Y=98510
X6512 2 digital_ldo_top_VIA4 $T=159730 102820 0 0 $X=159480 $Y=102590
X6513 2 digital_ldo_top_VIA4 $T=159730 106900 0 0 $X=159480 $Y=106670
X6514 2 digital_ldo_top_VIA4 $T=159730 110980 0 0 $X=159480 $Y=110750
X6515 2 digital_ldo_top_VIA4 $T=159730 115060 0 0 $X=159480 $Y=114830
X6516 2 digital_ldo_top_VIA4 $T=159730 119140 0 0 $X=159480 $Y=118910
X6517 2 digital_ldo_top_VIA4 $T=159730 123220 0 0 $X=159480 $Y=122990
X6518 2 digital_ldo_top_VIA4 $T=159730 127300 0 0 $X=159480 $Y=127070
X6519 3 digital_ldo_top_VIA4 $T=162030 11700 0 0 $X=161780 $Y=11470
X6520 3 digital_ldo_top_VIA4 $T=162030 15780 0 0 $X=161780 $Y=15550
X6521 3 digital_ldo_top_VIA4 $T=162030 85140 0 0 $X=161780 $Y=84910
X6522 3 digital_ldo_top_VIA4 $T=162030 89220 0 0 $X=161780 $Y=88990
X6523 3 digital_ldo_top_VIA4 $T=162030 93300 0 0 $X=161780 $Y=93070
X6524 3 digital_ldo_top_VIA4 $T=162030 97380 0 0 $X=161780 $Y=97150
X6525 3 digital_ldo_top_VIA4 $T=162030 101460 0 0 $X=161780 $Y=101230
X6526 3 digital_ldo_top_VIA4 $T=162030 105540 0 0 $X=161780 $Y=105310
X6527 3 digital_ldo_top_VIA4 $T=162030 109620 0 0 $X=161780 $Y=109390
X6528 3 digital_ldo_top_VIA4 $T=162030 113700 0 0 $X=161780 $Y=113470
X6529 3 digital_ldo_top_VIA4 $T=162030 117780 0 0 $X=161780 $Y=117550
X6530 3 digital_ldo_top_VIA4 $T=162030 121860 0 0 $X=161780 $Y=121630
X6531 3 digital_ldo_top_VIA4 $T=162030 125940 0 0 $X=161780 $Y=125710
X6532 2 digital_ldo_top_VIA4 $T=163410 13060 0 0 $X=163160 $Y=12830
X6533 2 digital_ldo_top_VIA4 $T=163410 17140 0 0 $X=163160 $Y=16910
X6534 2 digital_ldo_top_VIA4 $T=163410 21220 0 0 $X=163160 $Y=20990
X6535 2 digital_ldo_top_VIA4 $T=163410 25300 0 0 $X=163160 $Y=25070
X6536 2 digital_ldo_top_VIA4 $T=163410 94660 0 0 $X=163160 $Y=94430
X6537 2 digital_ldo_top_VIA4 $T=163410 98740 0 0 $X=163160 $Y=98510
X6538 2 digital_ldo_top_VIA4 $T=163410 102820 0 0 $X=163160 $Y=102590
X6539 2 digital_ldo_top_VIA4 $T=163410 106900 0 0 $X=163160 $Y=106670
X6540 2 digital_ldo_top_VIA4 $T=163410 110980 0 0 $X=163160 $Y=110750
X6541 2 digital_ldo_top_VIA4 $T=163410 115060 0 0 $X=163160 $Y=114830
X6542 2 digital_ldo_top_VIA4 $T=163410 119140 0 0 $X=163160 $Y=118910
X6543 2 digital_ldo_top_VIA4 $T=163410 123220 0 0 $X=163160 $Y=122990
X6544 2 digital_ldo_top_VIA4 $T=163410 127300 0 0 $X=163160 $Y=127070
X6545 3 digital_ldo_top_VIA4 $T=165710 11700 0 0 $X=165460 $Y=11470
X6546 3 digital_ldo_top_VIA4 $T=165710 15780 0 0 $X=165460 $Y=15550
X6547 3 digital_ldo_top_VIA4 $T=165710 19860 0 0 $X=165460 $Y=19630
X6548 3 digital_ldo_top_VIA4 $T=165710 23940 0 0 $X=165460 $Y=23710
X6549 3 digital_ldo_top_VIA4 $T=165710 32100 0 0 $X=165460 $Y=31870
X6550 3 digital_ldo_top_VIA4 $T=165710 85140 0 0 $X=165460 $Y=84910
X6551 3 digital_ldo_top_VIA4 $T=165710 89220 0 0 $X=165460 $Y=88990
X6552 3 digital_ldo_top_VIA4 $T=165710 93300 0 0 $X=165460 $Y=93070
X6553 3 digital_ldo_top_VIA4 $T=165710 97380 0 0 $X=165460 $Y=97150
X6554 3 digital_ldo_top_VIA4 $T=165710 101460 0 0 $X=165460 $Y=101230
X6555 3 digital_ldo_top_VIA4 $T=165710 105540 0 0 $X=165460 $Y=105310
X6556 3 digital_ldo_top_VIA4 $T=165710 109620 0 0 $X=165460 $Y=109390
X6557 3 digital_ldo_top_VIA4 $T=165710 113700 0 0 $X=165460 $Y=113470
X6558 3 digital_ldo_top_VIA4 $T=165710 117780 0 0 $X=165460 $Y=117550
X6559 3 digital_ldo_top_VIA4 $T=165710 121860 0 0 $X=165460 $Y=121630
X6560 3 digital_ldo_top_VIA4 $T=165710 125940 0 0 $X=165460 $Y=125710
X6561 2 digital_ldo_top_VIA4 $T=167090 13060 0 0 $X=166840 $Y=12830
X6562 2 digital_ldo_top_VIA4 $T=167090 17140 0 0 $X=166840 $Y=16910
X6563 2 digital_ldo_top_VIA4 $T=167090 21220 0 0 $X=166840 $Y=20990
X6564 2 digital_ldo_top_VIA4 $T=167090 25300 0 0 $X=166840 $Y=25070
X6565 2 digital_ldo_top_VIA4 $T=167090 86500 0 0 $X=166840 $Y=86270
X6566 2 digital_ldo_top_VIA4 $T=167090 90580 0 0 $X=166840 $Y=90350
X6567 2 digital_ldo_top_VIA4 $T=167090 94660 0 0 $X=166840 $Y=94430
X6568 2 digital_ldo_top_VIA4 $T=167090 98740 0 0 $X=166840 $Y=98510
X6569 2 digital_ldo_top_VIA4 $T=167090 102820 0 0 $X=166840 $Y=102590
X6570 2 digital_ldo_top_VIA4 $T=167090 106900 0 0 $X=166840 $Y=106670
X6571 2 digital_ldo_top_VIA4 $T=167090 110980 0 0 $X=166840 $Y=110750
X6572 2 digital_ldo_top_VIA4 $T=167090 115060 0 0 $X=166840 $Y=114830
X6573 2 digital_ldo_top_VIA4 $T=167090 119140 0 0 $X=166840 $Y=118910
X6574 2 digital_ldo_top_VIA4 $T=167090 123220 0 0 $X=166840 $Y=122990
X6575 2 digital_ldo_top_VIA4 $T=167090 127300 0 0 $X=166840 $Y=127070
X6576 3 digital_ldo_top_VIA4 $T=169390 11700 0 0 $X=169140 $Y=11470
X6577 3 digital_ldo_top_VIA4 $T=169390 15780 0 0 $X=169140 $Y=15550
X6578 3 digital_ldo_top_VIA4 $T=169390 93300 0 0 $X=169140 $Y=93070
X6579 3 digital_ldo_top_VIA4 $T=169390 97380 0 0 $X=169140 $Y=97150
X6580 3 digital_ldo_top_VIA4 $T=169390 101460 0 0 $X=169140 $Y=101230
X6581 3 digital_ldo_top_VIA4 $T=169390 105540 0 0 $X=169140 $Y=105310
X6582 3 digital_ldo_top_VIA4 $T=169390 109620 0 0 $X=169140 $Y=109390
X6583 3 digital_ldo_top_VIA4 $T=169390 113700 0 0 $X=169140 $Y=113470
X6584 3 digital_ldo_top_VIA4 $T=169390 117780 0 0 $X=169140 $Y=117550
X6585 3 digital_ldo_top_VIA4 $T=169390 121860 0 0 $X=169140 $Y=121630
X6586 3 digital_ldo_top_VIA4 $T=169390 125940 0 0 $X=169140 $Y=125710
X6587 2 digital_ldo_top_VIA4 $T=170770 13060 0 0 $X=170520 $Y=12830
X6588 2 digital_ldo_top_VIA4 $T=170770 17140 0 0 $X=170520 $Y=16910
X6589 2 digital_ldo_top_VIA4 $T=170770 94660 0 0 $X=170520 $Y=94430
X6590 2 digital_ldo_top_VIA4 $T=170770 98740 0 0 $X=170520 $Y=98510
X6591 2 digital_ldo_top_VIA4 $T=170770 102820 0 0 $X=170520 $Y=102590
X6592 2 digital_ldo_top_VIA4 $T=170770 106900 0 0 $X=170520 $Y=106670
X6593 2 digital_ldo_top_VIA4 $T=170770 110980 0 0 $X=170520 $Y=110750
X6594 2 digital_ldo_top_VIA4 $T=170770 115060 0 0 $X=170520 $Y=114830
X6595 2 digital_ldo_top_VIA4 $T=170770 119140 0 0 $X=170520 $Y=118910
X6596 2 digital_ldo_top_VIA4 $T=170770 123220 0 0 $X=170520 $Y=122990
X6597 2 digital_ldo_top_VIA4 $T=170770 127300 0 0 $X=170520 $Y=127070
X6598 3 digital_ldo_top_VIA4 $T=173070 11700 0 0 $X=172820 $Y=11470
X6599 3 digital_ldo_top_VIA4 $T=173070 15780 0 0 $X=172820 $Y=15550
X6600 3 digital_ldo_top_VIA4 $T=173070 85140 0 0 $X=172820 $Y=84910
X6601 3 digital_ldo_top_VIA4 $T=173070 89220 0 0 $X=172820 $Y=88990
X6602 3 digital_ldo_top_VIA4 $T=173070 93300 0 0 $X=172820 $Y=93070
X6603 3 digital_ldo_top_VIA4 $T=173070 97380 0 0 $X=172820 $Y=97150
X6604 3 digital_ldo_top_VIA4 $T=173070 101460 0 0 $X=172820 $Y=101230
X6605 3 digital_ldo_top_VIA4 $T=173070 105540 0 0 $X=172820 $Y=105310
X6606 3 digital_ldo_top_VIA4 $T=173070 109620 0 0 $X=172820 $Y=109390
X6607 3 digital_ldo_top_VIA4 $T=173070 113700 0 0 $X=172820 $Y=113470
X6608 3 digital_ldo_top_VIA4 $T=173070 117780 0 0 $X=172820 $Y=117550
X6609 3 digital_ldo_top_VIA4 $T=173070 121860 0 0 $X=172820 $Y=121630
X6610 3 digital_ldo_top_VIA4 $T=173070 125940 0 0 $X=172820 $Y=125710
X6611 2 digital_ldo_top_VIA4 $T=174450 13060 0 0 $X=174200 $Y=12830
X6612 2 digital_ldo_top_VIA4 $T=174450 17140 0 0 $X=174200 $Y=16910
X6613 2 digital_ldo_top_VIA4 $T=174450 21220 0 0 $X=174200 $Y=20990
X6614 2 digital_ldo_top_VIA4 $T=174450 25300 0 0 $X=174200 $Y=25070
X6615 2 digital_ldo_top_VIA4 $T=174450 94660 0 0 $X=174200 $Y=94430
X6616 2 digital_ldo_top_VIA4 $T=174450 98740 0 0 $X=174200 $Y=98510
X6617 2 digital_ldo_top_VIA4 $T=174450 102820 0 0 $X=174200 $Y=102590
X6618 2 digital_ldo_top_VIA4 $T=174450 106900 0 0 $X=174200 $Y=106670
X6619 2 digital_ldo_top_VIA4 $T=174450 110980 0 0 $X=174200 $Y=110750
X6620 2 digital_ldo_top_VIA4 $T=174450 115060 0 0 $X=174200 $Y=114830
X6621 2 digital_ldo_top_VIA4 $T=174450 119140 0 0 $X=174200 $Y=118910
X6622 2 digital_ldo_top_VIA4 $T=174450 123220 0 0 $X=174200 $Y=122990
X6623 2 digital_ldo_top_VIA4 $T=174450 127300 0 0 $X=174200 $Y=127070
X6624 3 digital_ldo_top_VIA4 $T=176750 11700 0 0 $X=176500 $Y=11470
X6625 3 digital_ldo_top_VIA4 $T=176750 15780 0 0 $X=176500 $Y=15550
X6626 3 digital_ldo_top_VIA4 $T=176750 19860 0 0 $X=176500 $Y=19630
X6627 3 digital_ldo_top_VIA4 $T=176750 23940 0 0 $X=176500 $Y=23710
X6628 3 digital_ldo_top_VIA4 $T=176750 32100 0 0 $X=176500 $Y=31870
X6629 3 digital_ldo_top_VIA4 $T=176750 85140 0 0 $X=176500 $Y=84910
X6630 3 digital_ldo_top_VIA4 $T=176750 89220 0 0 $X=176500 $Y=88990
X6631 3 digital_ldo_top_VIA4 $T=176750 93300 0 0 $X=176500 $Y=93070
X6632 3 digital_ldo_top_VIA4 $T=176750 97380 0 0 $X=176500 $Y=97150
X6633 3 digital_ldo_top_VIA4 $T=176750 101460 0 0 $X=176500 $Y=101230
X6634 3 digital_ldo_top_VIA4 $T=176750 105540 0 0 $X=176500 $Y=105310
X6635 3 digital_ldo_top_VIA4 $T=176750 109620 0 0 $X=176500 $Y=109390
X6636 3 digital_ldo_top_VIA4 $T=176750 113700 0 0 $X=176500 $Y=113470
X6637 3 digital_ldo_top_VIA4 $T=176750 117780 0 0 $X=176500 $Y=117550
X6638 3 digital_ldo_top_VIA4 $T=176750 121860 0 0 $X=176500 $Y=121630
X6639 3 digital_ldo_top_VIA4 $T=176750 125940 0 0 $X=176500 $Y=125710
X6640 2 digital_ldo_top_VIA4 $T=178130 13060 0 0 $X=177880 $Y=12830
X6641 2 digital_ldo_top_VIA4 $T=178130 17140 0 0 $X=177880 $Y=16910
X6642 2 digital_ldo_top_VIA4 $T=178130 21220 0 0 $X=177880 $Y=20990
X6643 2 digital_ldo_top_VIA4 $T=178130 25300 0 0 $X=177880 $Y=25070
X6644 2 digital_ldo_top_VIA4 $T=178130 86500 0 0 $X=177880 $Y=86270
X6645 2 digital_ldo_top_VIA4 $T=178130 90580 0 0 $X=177880 $Y=90350
X6646 2 digital_ldo_top_VIA4 $T=178130 94660 0 0 $X=177880 $Y=94430
X6647 2 digital_ldo_top_VIA4 $T=178130 98740 0 0 $X=177880 $Y=98510
X6648 2 digital_ldo_top_VIA4 $T=178130 102820 0 0 $X=177880 $Y=102590
X6649 2 digital_ldo_top_VIA4 $T=178130 106900 0 0 $X=177880 $Y=106670
X6650 2 digital_ldo_top_VIA4 $T=178130 110980 0 0 $X=177880 $Y=110750
X6651 2 digital_ldo_top_VIA4 $T=178130 115060 0 0 $X=177880 $Y=114830
X6652 2 digital_ldo_top_VIA4 $T=178130 119140 0 0 $X=177880 $Y=118910
X6653 2 digital_ldo_top_VIA4 $T=178130 123220 0 0 $X=177880 $Y=122990
X6654 2 digital_ldo_top_VIA4 $T=178130 127300 0 0 $X=177880 $Y=127070
X6655 3 digital_ldo_top_VIA4 $T=180430 11700 0 0 $X=180180 $Y=11470
X6656 3 digital_ldo_top_VIA4 $T=180430 15780 0 0 $X=180180 $Y=15550
X6657 3 digital_ldo_top_VIA4 $T=180430 93300 0 0 $X=180180 $Y=93070
X6658 3 digital_ldo_top_VIA4 $T=180430 97380 0 0 $X=180180 $Y=97150
X6659 3 digital_ldo_top_VIA4 $T=180430 101460 0 0 $X=180180 $Y=101230
X6660 3 digital_ldo_top_VIA4 $T=180430 105540 0 0 $X=180180 $Y=105310
X6661 3 digital_ldo_top_VIA4 $T=180430 109620 0 0 $X=180180 $Y=109390
X6662 3 digital_ldo_top_VIA4 $T=180430 113700 0 0 $X=180180 $Y=113470
X6663 3 digital_ldo_top_VIA4 $T=180430 117780 0 0 $X=180180 $Y=117550
X6664 3 digital_ldo_top_VIA4 $T=180430 121860 0 0 $X=180180 $Y=121630
X6665 3 digital_ldo_top_VIA4 $T=180430 125940 0 0 $X=180180 $Y=125710
X6666 2 digital_ldo_top_VIA4 $T=181810 13060 0 0 $X=181560 $Y=12830
X6667 2 digital_ldo_top_VIA4 $T=181810 17140 0 0 $X=181560 $Y=16910
X6668 2 digital_ldo_top_VIA4 $T=181810 94660 0 0 $X=181560 $Y=94430
X6669 2 digital_ldo_top_VIA4 $T=181810 98740 0 0 $X=181560 $Y=98510
X6670 2 digital_ldo_top_VIA4 $T=181810 102820 0 0 $X=181560 $Y=102590
X6671 2 digital_ldo_top_VIA4 $T=181810 106900 0 0 $X=181560 $Y=106670
X6672 2 digital_ldo_top_VIA4 $T=181810 110980 0 0 $X=181560 $Y=110750
X6673 2 digital_ldo_top_VIA4 $T=181810 115060 0 0 $X=181560 $Y=114830
X6674 2 digital_ldo_top_VIA4 $T=181810 119140 0 0 $X=181560 $Y=118910
X6675 2 digital_ldo_top_VIA4 $T=181810 123220 0 0 $X=181560 $Y=122990
X6676 2 digital_ldo_top_VIA4 $T=181810 127300 0 0 $X=181560 $Y=127070
X6677 3 digital_ldo_top_VIA4 $T=184110 11700 0 0 $X=183860 $Y=11470
X6678 3 digital_ldo_top_VIA4 $T=184110 15780 0 0 $X=183860 $Y=15550
X6679 3 digital_ldo_top_VIA4 $T=184110 85140 0 0 $X=183860 $Y=84910
X6680 3 digital_ldo_top_VIA4 $T=184110 89220 0 0 $X=183860 $Y=88990
X6681 3 digital_ldo_top_VIA4 $T=184110 93300 0 0 $X=183860 $Y=93070
X6682 3 digital_ldo_top_VIA4 $T=184110 97380 0 0 $X=183860 $Y=97150
X6683 3 digital_ldo_top_VIA4 $T=184110 101460 0 0 $X=183860 $Y=101230
X6684 3 digital_ldo_top_VIA4 $T=184110 105540 0 0 $X=183860 $Y=105310
X6685 3 digital_ldo_top_VIA4 $T=184110 109620 0 0 $X=183860 $Y=109390
X6686 3 digital_ldo_top_VIA4 $T=184110 113700 0 0 $X=183860 $Y=113470
X6687 3 digital_ldo_top_VIA4 $T=184110 117780 0 0 $X=183860 $Y=117550
X6688 3 digital_ldo_top_VIA4 $T=184110 121860 0 0 $X=183860 $Y=121630
X6689 3 digital_ldo_top_VIA4 $T=184110 125940 0 0 $X=183860 $Y=125710
X6690 2 digital_ldo_top_VIA4 $T=185490 13060 0 0 $X=185240 $Y=12830
X6691 2 digital_ldo_top_VIA4 $T=185490 17140 0 0 $X=185240 $Y=16910
X6692 2 digital_ldo_top_VIA4 $T=185490 21220 0 0 $X=185240 $Y=20990
X6693 2 digital_ldo_top_VIA4 $T=185490 25300 0 0 $X=185240 $Y=25070
X6694 2 digital_ldo_top_VIA4 $T=185490 94660 0 0 $X=185240 $Y=94430
X6695 2 digital_ldo_top_VIA4 $T=185490 98740 0 0 $X=185240 $Y=98510
X6696 2 digital_ldo_top_VIA4 $T=185490 102820 0 0 $X=185240 $Y=102590
X6697 2 digital_ldo_top_VIA4 $T=185490 106900 0 0 $X=185240 $Y=106670
X6698 2 digital_ldo_top_VIA4 $T=185490 110980 0 0 $X=185240 $Y=110750
X6699 2 digital_ldo_top_VIA4 $T=185490 115060 0 0 $X=185240 $Y=114830
X6700 2 digital_ldo_top_VIA4 $T=185490 119140 0 0 $X=185240 $Y=118910
X6701 2 digital_ldo_top_VIA4 $T=185490 123220 0 0 $X=185240 $Y=122990
X6702 2 digital_ldo_top_VIA4 $T=185490 127300 0 0 $X=185240 $Y=127070
X6703 3 digital_ldo_top_VIA4 $T=187790 11700 0 0 $X=187540 $Y=11470
X6704 3 digital_ldo_top_VIA4 $T=187790 15780 0 0 $X=187540 $Y=15550
X6705 3 digital_ldo_top_VIA4 $T=187790 19860 0 0 $X=187540 $Y=19630
X6706 3 digital_ldo_top_VIA4 $T=187790 23940 0 0 $X=187540 $Y=23710
X6707 3 digital_ldo_top_VIA4 $T=187790 32100 0 0 $X=187540 $Y=31870
X6708 3 digital_ldo_top_VIA4 $T=187790 85140 0 0 $X=187540 $Y=84910
X6709 3 digital_ldo_top_VIA4 $T=187790 89220 0 0 $X=187540 $Y=88990
X6710 3 digital_ldo_top_VIA4 $T=187790 93300 0 0 $X=187540 $Y=93070
X6711 3 digital_ldo_top_VIA4 $T=187790 97380 0 0 $X=187540 $Y=97150
X6712 3 digital_ldo_top_VIA4 $T=187790 101460 0 0 $X=187540 $Y=101230
X6713 3 digital_ldo_top_VIA4 $T=187790 105540 0 0 $X=187540 $Y=105310
X6714 3 digital_ldo_top_VIA4 $T=187790 109620 0 0 $X=187540 $Y=109390
X6715 3 digital_ldo_top_VIA4 $T=187790 113700 0 0 $X=187540 $Y=113470
X6716 3 digital_ldo_top_VIA4 $T=187790 117780 0 0 $X=187540 $Y=117550
X6717 3 digital_ldo_top_VIA4 $T=187790 121860 0 0 $X=187540 $Y=121630
X6718 3 digital_ldo_top_VIA4 $T=187790 125940 0 0 $X=187540 $Y=125710
X6719 2 digital_ldo_top_VIA4 $T=189170 13060 0 0 $X=188920 $Y=12830
X6720 2 digital_ldo_top_VIA4 $T=189170 17140 0 0 $X=188920 $Y=16910
X6721 2 digital_ldo_top_VIA4 $T=189170 21220 0 0 $X=188920 $Y=20990
X6722 2 digital_ldo_top_VIA4 $T=189170 25300 0 0 $X=188920 $Y=25070
X6723 2 digital_ldo_top_VIA4 $T=189170 86500 0 0 $X=188920 $Y=86270
X6724 2 digital_ldo_top_VIA4 $T=189170 90580 0 0 $X=188920 $Y=90350
X6725 2 digital_ldo_top_VIA4 $T=189170 94660 0 0 $X=188920 $Y=94430
X6726 2 digital_ldo_top_VIA4 $T=189170 98740 0 0 $X=188920 $Y=98510
X6727 2 digital_ldo_top_VIA4 $T=189170 102820 0 0 $X=188920 $Y=102590
X6728 2 digital_ldo_top_VIA4 $T=189170 106900 0 0 $X=188920 $Y=106670
X6729 2 digital_ldo_top_VIA4 $T=189170 110980 0 0 $X=188920 $Y=110750
X6730 2 digital_ldo_top_VIA4 $T=189170 115060 0 0 $X=188920 $Y=114830
X6731 2 digital_ldo_top_VIA4 $T=189170 119140 0 0 $X=188920 $Y=118910
X6732 2 digital_ldo_top_VIA4 $T=189170 123220 0 0 $X=188920 $Y=122990
X6733 2 digital_ldo_top_VIA4 $T=189170 127300 0 0 $X=188920 $Y=127070
X6734 3 digital_ldo_top_VIA4 $T=191470 11700 0 0 $X=191220 $Y=11470
X6735 3 digital_ldo_top_VIA4 $T=191470 15780 0 0 $X=191220 $Y=15550
X6736 3 digital_ldo_top_VIA4 $T=191470 93300 0 0 $X=191220 $Y=93070
X6737 3 digital_ldo_top_VIA4 $T=191470 97380 0 0 $X=191220 $Y=97150
X6738 3 digital_ldo_top_VIA4 $T=191470 101460 0 0 $X=191220 $Y=101230
X6739 3 digital_ldo_top_VIA4 $T=191470 105540 0 0 $X=191220 $Y=105310
X6740 3 digital_ldo_top_VIA4 $T=191470 109620 0 0 $X=191220 $Y=109390
X6741 3 digital_ldo_top_VIA4 $T=191470 113700 0 0 $X=191220 $Y=113470
X6742 3 digital_ldo_top_VIA4 $T=191470 117780 0 0 $X=191220 $Y=117550
X6743 3 digital_ldo_top_VIA4 $T=191470 121860 0 0 $X=191220 $Y=121630
X6744 3 digital_ldo_top_VIA4 $T=191470 125940 0 0 $X=191220 $Y=125710
X6745 2 digital_ldo_top_VIA4 $T=192850 13060 0 0 $X=192600 $Y=12830
X6746 2 digital_ldo_top_VIA4 $T=192850 17140 0 0 $X=192600 $Y=16910
X6747 2 digital_ldo_top_VIA4 $T=192850 21220 0 0 $X=192600 $Y=20990
X6748 2 digital_ldo_top_VIA4 $T=192850 25300 0 0 $X=192600 $Y=25070
X6749 2 digital_ldo_top_VIA4 $T=192850 94660 0 0 $X=192600 $Y=94430
X6750 2 digital_ldo_top_VIA4 $T=192850 98740 0 0 $X=192600 $Y=98510
X6751 2 digital_ldo_top_VIA4 $T=192850 102820 0 0 $X=192600 $Y=102590
X6752 2 digital_ldo_top_VIA4 $T=192850 106900 0 0 $X=192600 $Y=106670
X6753 2 digital_ldo_top_VIA4 $T=192850 110980 0 0 $X=192600 $Y=110750
X6754 2 digital_ldo_top_VIA4 $T=192850 115060 0 0 $X=192600 $Y=114830
X6755 2 digital_ldo_top_VIA4 $T=192850 119140 0 0 $X=192600 $Y=118910
X6756 2 digital_ldo_top_VIA4 $T=192850 123220 0 0 $X=192600 $Y=122990
X6757 2 digital_ldo_top_VIA4 $T=192850 127300 0 0 $X=192600 $Y=127070
X6758 3 digital_ldo_top_VIA4 $T=195150 11700 0 0 $X=194900 $Y=11470
X6759 3 digital_ldo_top_VIA4 $T=195150 15780 0 0 $X=194900 $Y=15550
X6760 3 digital_ldo_top_VIA4 $T=195150 85140 0 0 $X=194900 $Y=84910
X6761 3 digital_ldo_top_VIA4 $T=195150 89220 0 0 $X=194900 $Y=88990
X6762 3 digital_ldo_top_VIA4 $T=195150 93300 0 0 $X=194900 $Y=93070
X6763 3 digital_ldo_top_VIA4 $T=195150 97380 0 0 $X=194900 $Y=97150
X6764 3 digital_ldo_top_VIA4 $T=195150 101460 0 0 $X=194900 $Y=101230
X6765 3 digital_ldo_top_VIA4 $T=195150 105540 0 0 $X=194900 $Y=105310
X6766 3 digital_ldo_top_VIA4 $T=195150 109620 0 0 $X=194900 $Y=109390
X6767 3 digital_ldo_top_VIA4 $T=195150 113700 0 0 $X=194900 $Y=113470
X6768 3 digital_ldo_top_VIA4 $T=195150 117780 0 0 $X=194900 $Y=117550
X6769 3 digital_ldo_top_VIA4 $T=195150 121860 0 0 $X=194900 $Y=121630
X6770 3 digital_ldo_top_VIA4 $T=195150 125940 0 0 $X=194900 $Y=125710
X6771 2 digital_ldo_top_VIA4 $T=196530 13060 0 0 $X=196280 $Y=12830
X6772 2 digital_ldo_top_VIA4 $T=196530 17140 0 0 $X=196280 $Y=16910
X6773 2 digital_ldo_top_VIA4 $T=196530 21220 0 0 $X=196280 $Y=20990
X6774 2 digital_ldo_top_VIA4 $T=196530 25300 0 0 $X=196280 $Y=25070
X6775 2 digital_ldo_top_VIA4 $T=196530 94660 0 0 $X=196280 $Y=94430
X6776 2 digital_ldo_top_VIA4 $T=196530 98740 0 0 $X=196280 $Y=98510
X6777 2 digital_ldo_top_VIA4 $T=196530 102820 0 0 $X=196280 $Y=102590
X6778 2 digital_ldo_top_VIA4 $T=196530 106900 0 0 $X=196280 $Y=106670
X6779 2 digital_ldo_top_VIA4 $T=196530 110980 0 0 $X=196280 $Y=110750
X6780 2 digital_ldo_top_VIA4 $T=196530 115060 0 0 $X=196280 $Y=114830
X6781 2 digital_ldo_top_VIA4 $T=196530 119140 0 0 $X=196280 $Y=118910
X6782 2 digital_ldo_top_VIA4 $T=196530 123220 0 0 $X=196280 $Y=122990
X6783 2 digital_ldo_top_VIA4 $T=196530 127300 0 0 $X=196280 $Y=127070
X6784 3 digital_ldo_top_VIA4 $T=198830 11700 0 0 $X=198580 $Y=11470
X6785 3 digital_ldo_top_VIA4 $T=198830 15780 0 0 $X=198580 $Y=15550
X6786 3 digital_ldo_top_VIA4 $T=198830 19860 0 0 $X=198580 $Y=19630
X6787 3 digital_ldo_top_VIA4 $T=198830 23940 0 0 $X=198580 $Y=23710
X6788 3 digital_ldo_top_VIA4 $T=198830 32100 0 0 $X=198580 $Y=31870
X6789 3 digital_ldo_top_VIA4 $T=198830 85140 0 0 $X=198580 $Y=84910
X6790 3 digital_ldo_top_VIA4 $T=198830 89220 0 0 $X=198580 $Y=88990
X6791 3 digital_ldo_top_VIA4 $T=198830 93300 0 0 $X=198580 $Y=93070
X6792 3 digital_ldo_top_VIA4 $T=198830 97380 0 0 $X=198580 $Y=97150
X6793 3 digital_ldo_top_VIA4 $T=198830 101460 0 0 $X=198580 $Y=101230
X6794 3 digital_ldo_top_VIA4 $T=198830 105540 0 0 $X=198580 $Y=105310
X6795 3 digital_ldo_top_VIA4 $T=198830 109620 0 0 $X=198580 $Y=109390
X6796 3 digital_ldo_top_VIA4 $T=198830 113700 0 0 $X=198580 $Y=113470
X6797 3 digital_ldo_top_VIA4 $T=198830 117780 0 0 $X=198580 $Y=117550
X6798 3 digital_ldo_top_VIA4 $T=198830 121860 0 0 $X=198580 $Y=121630
X6799 3 digital_ldo_top_VIA4 $T=198830 125940 0 0 $X=198580 $Y=125710
X6800 2 digital_ldo_top_VIA4 $T=200210 13060 0 0 $X=199960 $Y=12830
X6801 2 digital_ldo_top_VIA4 $T=200210 17140 0 0 $X=199960 $Y=16910
X6802 2 digital_ldo_top_VIA4 $T=200210 86500 0 0 $X=199960 $Y=86270
X6803 2 digital_ldo_top_VIA4 $T=200210 90580 0 0 $X=199960 $Y=90350
X6804 2 digital_ldo_top_VIA4 $T=200210 94660 0 0 $X=199960 $Y=94430
X6805 2 digital_ldo_top_VIA4 $T=200210 98740 0 0 $X=199960 $Y=98510
X6806 2 digital_ldo_top_VIA4 $T=200210 102820 0 0 $X=199960 $Y=102590
X6807 2 digital_ldo_top_VIA4 $T=200210 106900 0 0 $X=199960 $Y=106670
X6808 2 digital_ldo_top_VIA4 $T=200210 110980 0 0 $X=199960 $Y=110750
X6809 2 digital_ldo_top_VIA4 $T=200210 115060 0 0 $X=199960 $Y=114830
X6810 2 digital_ldo_top_VIA4 $T=200210 119140 0 0 $X=199960 $Y=118910
X6811 2 digital_ldo_top_VIA4 $T=200210 123220 0 0 $X=199960 $Y=122990
X6812 2 digital_ldo_top_VIA4 $T=200210 127300 0 0 $X=199960 $Y=127070
X6813 3 digital_ldo_top_VIA4 $T=202510 11700 0 0 $X=202260 $Y=11470
X6814 3 digital_ldo_top_VIA4 $T=202510 15780 0 0 $X=202260 $Y=15550
X6815 3 digital_ldo_top_VIA4 $T=202510 93300 0 0 $X=202260 $Y=93070
X6816 3 digital_ldo_top_VIA4 $T=202510 97380 0 0 $X=202260 $Y=97150
X6817 3 digital_ldo_top_VIA4 $T=202510 101460 0 0 $X=202260 $Y=101230
X6818 3 digital_ldo_top_VIA4 $T=202510 105540 0 0 $X=202260 $Y=105310
X6819 3 digital_ldo_top_VIA4 $T=202510 109620 0 0 $X=202260 $Y=109390
X6820 3 digital_ldo_top_VIA4 $T=202510 113700 0 0 $X=202260 $Y=113470
X6821 3 digital_ldo_top_VIA4 $T=202510 117780 0 0 $X=202260 $Y=117550
X6822 3 digital_ldo_top_VIA4 $T=202510 121860 0 0 $X=202260 $Y=121630
X6823 3 digital_ldo_top_VIA4 $T=202510 125940 0 0 $X=202260 $Y=125710
X6824 2 digital_ldo_top_VIA4 $T=203890 13060 0 0 $X=203640 $Y=12830
X6825 2 digital_ldo_top_VIA4 $T=203890 17140 0 0 $X=203640 $Y=16910
X6826 2 digital_ldo_top_VIA4 $T=203890 21220 0 0 $X=203640 $Y=20990
X6827 2 digital_ldo_top_VIA4 $T=203890 25300 0 0 $X=203640 $Y=25070
X6828 2 digital_ldo_top_VIA4 $T=203890 94660 0 0 $X=203640 $Y=94430
X6829 2 digital_ldo_top_VIA4 $T=203890 98740 0 0 $X=203640 $Y=98510
X6830 2 digital_ldo_top_VIA4 $T=203890 102820 0 0 $X=203640 $Y=102590
X6831 2 digital_ldo_top_VIA4 $T=203890 106900 0 0 $X=203640 $Y=106670
X6832 2 digital_ldo_top_VIA4 $T=203890 110980 0 0 $X=203640 $Y=110750
X6833 2 digital_ldo_top_VIA4 $T=203890 115060 0 0 $X=203640 $Y=114830
X6834 2 digital_ldo_top_VIA4 $T=203890 119140 0 0 $X=203640 $Y=118910
X6835 2 digital_ldo_top_VIA4 $T=203890 123220 0 0 $X=203640 $Y=122990
X6836 2 digital_ldo_top_VIA4 $T=203890 127300 0 0 $X=203640 $Y=127070
X6837 3 digital_ldo_top_VIA4 $T=206190 11700 0 0 $X=205940 $Y=11470
X6838 3 digital_ldo_top_VIA4 $T=206190 15780 0 0 $X=205940 $Y=15550
X6839 3 digital_ldo_top_VIA4 $T=206190 85140 0 0 $X=205940 $Y=84910
X6840 3 digital_ldo_top_VIA4 $T=206190 89220 0 0 $X=205940 $Y=88990
X6841 3 digital_ldo_top_VIA4 $T=206190 93300 0 0 $X=205940 $Y=93070
X6842 3 digital_ldo_top_VIA4 $T=206190 97380 0 0 $X=205940 $Y=97150
X6843 3 digital_ldo_top_VIA4 $T=206190 101460 0 0 $X=205940 $Y=101230
X6844 3 digital_ldo_top_VIA4 $T=206190 105540 0 0 $X=205940 $Y=105310
X6845 3 digital_ldo_top_VIA4 $T=206190 109620 0 0 $X=205940 $Y=109390
X6846 3 digital_ldo_top_VIA4 $T=206190 113700 0 0 $X=205940 $Y=113470
X6847 3 digital_ldo_top_VIA4 $T=206190 117780 0 0 $X=205940 $Y=117550
X6848 3 digital_ldo_top_VIA4 $T=206190 121860 0 0 $X=205940 $Y=121630
X6849 3 digital_ldo_top_VIA4 $T=206190 125940 0 0 $X=205940 $Y=125710
X6850 2 digital_ldo_top_VIA4 $T=207570 13060 0 0 $X=207320 $Y=12830
X6851 2 digital_ldo_top_VIA4 $T=207570 17140 0 0 $X=207320 $Y=16910
X6852 2 digital_ldo_top_VIA4 $T=207570 21220 0 0 $X=207320 $Y=20990
X6853 2 digital_ldo_top_VIA4 $T=207570 25300 0 0 $X=207320 $Y=25070
X6854 2 digital_ldo_top_VIA4 $T=207570 94660 0 0 $X=207320 $Y=94430
X6855 2 digital_ldo_top_VIA4 $T=207570 98740 0 0 $X=207320 $Y=98510
X6856 2 digital_ldo_top_VIA4 $T=207570 102820 0 0 $X=207320 $Y=102590
X6857 2 digital_ldo_top_VIA4 $T=207570 106900 0 0 $X=207320 $Y=106670
X6858 2 digital_ldo_top_VIA4 $T=207570 110980 0 0 $X=207320 $Y=110750
X6859 2 digital_ldo_top_VIA4 $T=207570 115060 0 0 $X=207320 $Y=114830
X6860 2 digital_ldo_top_VIA4 $T=207570 119140 0 0 $X=207320 $Y=118910
X6861 2 digital_ldo_top_VIA4 $T=207570 123220 0 0 $X=207320 $Y=122990
X6862 2 digital_ldo_top_VIA4 $T=207570 127300 0 0 $X=207320 $Y=127070
X6863 3 digital_ldo_top_VIA4 $T=209870 11700 0 0 $X=209620 $Y=11470
X6864 3 digital_ldo_top_VIA4 $T=209870 15780 0 0 $X=209620 $Y=15550
X6865 3 digital_ldo_top_VIA4 $T=209870 32100 0 0 $X=209620 $Y=31870
X6866 3 digital_ldo_top_VIA4 $T=209870 85140 0 0 $X=209620 $Y=84910
X6867 3 digital_ldo_top_VIA4 $T=209870 89220 0 0 $X=209620 $Y=88990
X6868 3 digital_ldo_top_VIA4 $T=209870 93300 0 0 $X=209620 $Y=93070
X6869 3 digital_ldo_top_VIA4 $T=209870 97380 0 0 $X=209620 $Y=97150
X6870 3 digital_ldo_top_VIA4 $T=209870 101460 0 0 $X=209620 $Y=101230
X6871 3 digital_ldo_top_VIA4 $T=209870 105540 0 0 $X=209620 $Y=105310
X6872 3 digital_ldo_top_VIA4 $T=209870 109620 0 0 $X=209620 $Y=109390
X6873 3 digital_ldo_top_VIA4 $T=209870 113700 0 0 $X=209620 $Y=113470
X6874 3 digital_ldo_top_VIA4 $T=209870 117780 0 0 $X=209620 $Y=117550
X6875 3 digital_ldo_top_VIA4 $T=209870 121860 0 0 $X=209620 $Y=121630
X6876 3 digital_ldo_top_VIA4 $T=209870 125940 0 0 $X=209620 $Y=125710
X6877 2 digital_ldo_top_VIA4 $T=211250 13060 0 0 $X=211000 $Y=12830
X6878 2 digital_ldo_top_VIA4 $T=211250 17140 0 0 $X=211000 $Y=16910
X6879 2 digital_ldo_top_VIA4 $T=211250 21220 0 0 $X=211000 $Y=20990
X6880 2 digital_ldo_top_VIA4 $T=211250 25300 0 0 $X=211000 $Y=25070
X6881 2 digital_ldo_top_VIA4 $T=211250 86500 0 0 $X=211000 $Y=86270
X6882 2 digital_ldo_top_VIA4 $T=211250 90580 0 0 $X=211000 $Y=90350
X6883 2 digital_ldo_top_VIA4 $T=211250 94660 0 0 $X=211000 $Y=94430
X6884 2 digital_ldo_top_VIA4 $T=211250 98740 0 0 $X=211000 $Y=98510
X6885 2 digital_ldo_top_VIA4 $T=211250 102820 0 0 $X=211000 $Y=102590
X6886 2 digital_ldo_top_VIA4 $T=211250 106900 0 0 $X=211000 $Y=106670
X6887 2 digital_ldo_top_VIA4 $T=211250 110980 0 0 $X=211000 $Y=110750
X6888 2 digital_ldo_top_VIA4 $T=211250 115060 0 0 $X=211000 $Y=114830
X6889 2 digital_ldo_top_VIA4 $T=211250 119140 0 0 $X=211000 $Y=118910
X6890 2 digital_ldo_top_VIA4 $T=211250 123220 0 0 $X=211000 $Y=122990
X6891 2 digital_ldo_top_VIA4 $T=211250 127300 0 0 $X=211000 $Y=127070
X6892 3 digital_ldo_top_VIA4 $T=213550 11700 0 0 $X=213300 $Y=11470
X6893 3 digital_ldo_top_VIA4 $T=213550 15780 0 0 $X=213300 $Y=15550
X6894 3 digital_ldo_top_VIA4 $T=213550 93300 0 0 $X=213300 $Y=93070
X6895 3 digital_ldo_top_VIA4 $T=213550 97380 0 0 $X=213300 $Y=97150
X6896 3 digital_ldo_top_VIA4 $T=213550 101460 0 0 $X=213300 $Y=101230
X6897 3 digital_ldo_top_VIA4 $T=213550 105540 0 0 $X=213300 $Y=105310
X6898 3 digital_ldo_top_VIA4 $T=213550 109620 0 0 $X=213300 $Y=109390
X6899 3 digital_ldo_top_VIA4 $T=213550 113700 0 0 $X=213300 $Y=113470
X6900 3 digital_ldo_top_VIA4 $T=213550 117780 0 0 $X=213300 $Y=117550
X6901 3 digital_ldo_top_VIA4 $T=213550 121860 0 0 $X=213300 $Y=121630
X6902 3 digital_ldo_top_VIA4 $T=213550 125940 0 0 $X=213300 $Y=125710
X6903 2 digital_ldo_top_VIA4 $T=214930 13060 0 0 $X=214680 $Y=12830
X6904 2 digital_ldo_top_VIA4 $T=214930 17140 0 0 $X=214680 $Y=16910
X6905 2 digital_ldo_top_VIA4 $T=214930 21220 0 0 $X=214680 $Y=20990
X6906 2 digital_ldo_top_VIA4 $T=214930 25300 0 0 $X=214680 $Y=25070
X6907 2 digital_ldo_top_VIA4 $T=214930 94660 0 0 $X=214680 $Y=94430
X6908 2 digital_ldo_top_VIA4 $T=214930 98740 0 0 $X=214680 $Y=98510
X6909 2 digital_ldo_top_VIA4 $T=214930 102820 0 0 $X=214680 $Y=102590
X6910 2 digital_ldo_top_VIA4 $T=214930 106900 0 0 $X=214680 $Y=106670
X6911 2 digital_ldo_top_VIA4 $T=214930 110980 0 0 $X=214680 $Y=110750
X6912 2 digital_ldo_top_VIA4 $T=214930 115060 0 0 $X=214680 $Y=114830
X6913 2 digital_ldo_top_VIA4 $T=214930 119140 0 0 $X=214680 $Y=118910
X6914 2 digital_ldo_top_VIA4 $T=214930 123220 0 0 $X=214680 $Y=122990
X6915 2 digital_ldo_top_VIA4 $T=214930 127300 0 0 $X=214680 $Y=127070
X6916 3 digital_ldo_top_VIA4 $T=217230 11700 0 0 $X=216980 $Y=11470
X6917 3 digital_ldo_top_VIA4 $T=217230 15780 0 0 $X=216980 $Y=15550
X6918 3 digital_ldo_top_VIA4 $T=217230 19860 0 0 $X=216980 $Y=19630
X6919 3 digital_ldo_top_VIA4 $T=217230 23940 0 0 $X=216980 $Y=23710
X6920 3 digital_ldo_top_VIA4 $T=217230 32100 0 0 $X=216980 $Y=31870
X6921 3 digital_ldo_top_VIA4 $T=217230 85140 0 0 $X=216980 $Y=84910
X6922 3 digital_ldo_top_VIA4 $T=217230 89220 0 0 $X=216980 $Y=88990
X6923 3 digital_ldo_top_VIA4 $T=217230 93300 0 0 $X=216980 $Y=93070
X6924 3 digital_ldo_top_VIA4 $T=217230 97380 0 0 $X=216980 $Y=97150
X6925 3 digital_ldo_top_VIA4 $T=217230 101460 0 0 $X=216980 $Y=101230
X6926 3 digital_ldo_top_VIA4 $T=217230 105540 0 0 $X=216980 $Y=105310
X6927 3 digital_ldo_top_VIA4 $T=217230 109620 0 0 $X=216980 $Y=109390
X6928 3 digital_ldo_top_VIA4 $T=217230 113700 0 0 $X=216980 $Y=113470
X6929 3 digital_ldo_top_VIA4 $T=217230 117780 0 0 $X=216980 $Y=117550
X6930 3 digital_ldo_top_VIA4 $T=217230 121860 0 0 $X=216980 $Y=121630
X6931 3 digital_ldo_top_VIA4 $T=217230 125940 0 0 $X=216980 $Y=125710
X6932 2 digital_ldo_top_VIA4 $T=218610 13060 0 0 $X=218360 $Y=12830
X6933 2 digital_ldo_top_VIA4 $T=218610 17140 0 0 $X=218360 $Y=16910
X6934 2 digital_ldo_top_VIA4 $T=218610 21220 0 0 $X=218360 $Y=20990
X6935 2 digital_ldo_top_VIA4 $T=218610 25300 0 0 $X=218360 $Y=25070
X6936 2 digital_ldo_top_VIA4 $T=218610 94660 0 0 $X=218360 $Y=94430
X6937 2 digital_ldo_top_VIA4 $T=218610 98740 0 0 $X=218360 $Y=98510
X6938 2 digital_ldo_top_VIA4 $T=218610 102820 0 0 $X=218360 $Y=102590
X6939 2 digital_ldo_top_VIA4 $T=218610 106900 0 0 $X=218360 $Y=106670
X6940 2 digital_ldo_top_VIA4 $T=218610 110980 0 0 $X=218360 $Y=110750
X6941 2 digital_ldo_top_VIA4 $T=218610 115060 0 0 $X=218360 $Y=114830
X6942 2 digital_ldo_top_VIA4 $T=218610 119140 0 0 $X=218360 $Y=118910
X6943 2 digital_ldo_top_VIA4 $T=218610 123220 0 0 $X=218360 $Y=122990
X6944 2 digital_ldo_top_VIA4 $T=218610 127300 0 0 $X=218360 $Y=127070
X6945 3 digital_ldo_top_VIA4 $T=220910 11700 0 0 $X=220660 $Y=11470
X6946 3 digital_ldo_top_VIA4 $T=220910 15780 0 0 $X=220660 $Y=15550
X6947 3 digital_ldo_top_VIA4 $T=220910 19860 0 0 $X=220660 $Y=19630
X6948 3 digital_ldo_top_VIA4 $T=220910 23940 0 0 $X=220660 $Y=23710
X6949 3 digital_ldo_top_VIA4 $T=220910 32100 0 0 $X=220660 $Y=31870
X6950 3 digital_ldo_top_VIA4 $T=220910 85140 0 0 $X=220660 $Y=84910
X6951 3 digital_ldo_top_VIA4 $T=220910 89220 0 0 $X=220660 $Y=88990
X6952 3 digital_ldo_top_VIA4 $T=220910 93300 0 0 $X=220660 $Y=93070
X6953 3 digital_ldo_top_VIA4 $T=220910 97380 0 0 $X=220660 $Y=97150
X6954 3 digital_ldo_top_VIA4 $T=220910 101460 0 0 $X=220660 $Y=101230
X6955 3 digital_ldo_top_VIA4 $T=220910 105540 0 0 $X=220660 $Y=105310
X6956 3 digital_ldo_top_VIA4 $T=220910 109620 0 0 $X=220660 $Y=109390
X6957 3 digital_ldo_top_VIA4 $T=220910 113700 0 0 $X=220660 $Y=113470
X6958 3 digital_ldo_top_VIA4 $T=220910 117780 0 0 $X=220660 $Y=117550
X6959 3 digital_ldo_top_VIA4 $T=220910 121860 0 0 $X=220660 $Y=121630
X6960 3 digital_ldo_top_VIA4 $T=220910 125940 0 0 $X=220660 $Y=125710
X6961 2 digital_ldo_top_VIA4 $T=222290 13060 0 0 $X=222040 $Y=12830
X6962 2 digital_ldo_top_VIA4 $T=222290 17140 0 0 $X=222040 $Y=16910
X6963 2 digital_ldo_top_VIA4 $T=222290 21220 0 0 $X=222040 $Y=20990
X6964 2 digital_ldo_top_VIA4 $T=222290 25300 0 0 $X=222040 $Y=25070
X6965 2 digital_ldo_top_VIA4 $T=222290 86500 0 0 $X=222040 $Y=86270
X6966 2 digital_ldo_top_VIA4 $T=222290 90580 0 0 $X=222040 $Y=90350
X6967 2 digital_ldo_top_VIA4 $T=222290 94660 0 0 $X=222040 $Y=94430
X6968 2 digital_ldo_top_VIA4 $T=222290 98740 0 0 $X=222040 $Y=98510
X6969 2 digital_ldo_top_VIA4 $T=222290 102820 0 0 $X=222040 $Y=102590
X6970 2 digital_ldo_top_VIA4 $T=222290 106900 0 0 $X=222040 $Y=106670
X6971 2 digital_ldo_top_VIA4 $T=222290 110980 0 0 $X=222040 $Y=110750
X6972 2 digital_ldo_top_VIA4 $T=222290 115060 0 0 $X=222040 $Y=114830
X6973 2 digital_ldo_top_VIA4 $T=222290 119140 0 0 $X=222040 $Y=118910
X6974 2 digital_ldo_top_VIA4 $T=222290 123220 0 0 $X=222040 $Y=122990
X6975 2 digital_ldo_top_VIA4 $T=222290 127300 0 0 $X=222040 $Y=127070
X6976 3 digital_ldo_top_VIA4 $T=224590 11700 0 0 $X=224340 $Y=11470
X6977 3 digital_ldo_top_VIA4 $T=224590 15780 0 0 $X=224340 $Y=15550
X6978 3 digital_ldo_top_VIA4 $T=224590 93300 0 0 $X=224340 $Y=93070
X6979 3 digital_ldo_top_VIA4 $T=224590 97380 0 0 $X=224340 $Y=97150
X6980 3 digital_ldo_top_VIA4 $T=224590 101460 0 0 $X=224340 $Y=101230
X6981 3 digital_ldo_top_VIA4 $T=224590 105540 0 0 $X=224340 $Y=105310
X6982 3 digital_ldo_top_VIA4 $T=224590 109620 0 0 $X=224340 $Y=109390
X6983 3 digital_ldo_top_VIA4 $T=224590 113700 0 0 $X=224340 $Y=113470
X6984 3 digital_ldo_top_VIA4 $T=224590 117780 0 0 $X=224340 $Y=117550
X6985 3 digital_ldo_top_VIA4 $T=224590 121860 0 0 $X=224340 $Y=121630
X6986 3 digital_ldo_top_VIA4 $T=224590 125940 0 0 $X=224340 $Y=125710
X6987 2 digital_ldo_top_VIA4 $T=225970 13060 0 0 $X=225720 $Y=12830
X6988 2 digital_ldo_top_VIA4 $T=225970 17140 0 0 $X=225720 $Y=16910
X6989 2 digital_ldo_top_VIA4 $T=225970 21220 0 0 $X=225720 $Y=20990
X6990 2 digital_ldo_top_VIA4 $T=225970 25300 0 0 $X=225720 $Y=25070
X6991 2 digital_ldo_top_VIA4 $T=225970 94660 0 0 $X=225720 $Y=94430
X6992 2 digital_ldo_top_VIA4 $T=225970 98740 0 0 $X=225720 $Y=98510
X6993 2 digital_ldo_top_VIA4 $T=225970 102820 0 0 $X=225720 $Y=102590
X6994 2 digital_ldo_top_VIA4 $T=225970 106900 0 0 $X=225720 $Y=106670
X6995 2 digital_ldo_top_VIA4 $T=225970 110980 0 0 $X=225720 $Y=110750
X6996 2 digital_ldo_top_VIA4 $T=225970 115060 0 0 $X=225720 $Y=114830
X6997 2 digital_ldo_top_VIA4 $T=225970 119140 0 0 $X=225720 $Y=118910
X6998 2 digital_ldo_top_VIA4 $T=225970 123220 0 0 $X=225720 $Y=122990
X6999 2 digital_ldo_top_VIA4 $T=225970 127300 0 0 $X=225720 $Y=127070
X7000 3 digital_ldo_top_VIA4 $T=228270 11700 0 0 $X=228020 $Y=11470
X7001 3 digital_ldo_top_VIA4 $T=228270 15780 0 0 $X=228020 $Y=15550
X7002 3 digital_ldo_top_VIA4 $T=228270 85140 0 0 $X=228020 $Y=84910
X7003 3 digital_ldo_top_VIA4 $T=228270 89220 0 0 $X=228020 $Y=88990
X7004 3 digital_ldo_top_VIA4 $T=228270 93300 0 0 $X=228020 $Y=93070
X7005 3 digital_ldo_top_VIA4 $T=228270 97380 0 0 $X=228020 $Y=97150
X7006 3 digital_ldo_top_VIA4 $T=228270 101460 0 0 $X=228020 $Y=101230
X7007 3 digital_ldo_top_VIA4 $T=228270 105540 0 0 $X=228020 $Y=105310
X7008 3 digital_ldo_top_VIA4 $T=228270 109620 0 0 $X=228020 $Y=109390
X7009 3 digital_ldo_top_VIA4 $T=228270 113700 0 0 $X=228020 $Y=113470
X7010 3 digital_ldo_top_VIA4 $T=228270 117780 0 0 $X=228020 $Y=117550
X7011 3 digital_ldo_top_VIA4 $T=228270 121860 0 0 $X=228020 $Y=121630
X7012 3 digital_ldo_top_VIA4 $T=228270 125940 0 0 $X=228020 $Y=125710
X7013 2 digital_ldo_top_VIA4 $T=229650 13060 0 0 $X=229400 $Y=12830
X7014 2 digital_ldo_top_VIA4 $T=229650 17140 0 0 $X=229400 $Y=16910
X7015 2 digital_ldo_top_VIA4 $T=229650 21220 0 0 $X=229400 $Y=20990
X7016 2 digital_ldo_top_VIA4 $T=229650 25300 0 0 $X=229400 $Y=25070
X7017 2 digital_ldo_top_VIA4 $T=229650 94660 0 0 $X=229400 $Y=94430
X7018 2 digital_ldo_top_VIA4 $T=229650 98740 0 0 $X=229400 $Y=98510
X7019 2 digital_ldo_top_VIA4 $T=229650 102820 0 0 $X=229400 $Y=102590
X7020 2 digital_ldo_top_VIA4 $T=229650 106900 0 0 $X=229400 $Y=106670
X7021 2 digital_ldo_top_VIA4 $T=229650 110980 0 0 $X=229400 $Y=110750
X7022 2 digital_ldo_top_VIA4 $T=229650 115060 0 0 $X=229400 $Y=114830
X7023 2 digital_ldo_top_VIA4 $T=229650 119140 0 0 $X=229400 $Y=118910
X7024 2 digital_ldo_top_VIA4 $T=229650 123220 0 0 $X=229400 $Y=122990
X7025 2 digital_ldo_top_VIA4 $T=229650 127300 0 0 $X=229400 $Y=127070
X7026 3 digital_ldo_top_VIA4 $T=231950 11700 0 0 $X=231700 $Y=11470
X7027 3 digital_ldo_top_VIA4 $T=231950 15780 0 0 $X=231700 $Y=15550
X7028 3 digital_ldo_top_VIA4 $T=231950 19860 0 0 $X=231700 $Y=19630
X7029 3 digital_ldo_top_VIA4 $T=231950 23940 0 0 $X=231700 $Y=23710
X7030 3 digital_ldo_top_VIA4 $T=231950 32100 0 0 $X=231700 $Y=31870
X7031 3 digital_ldo_top_VIA4 $T=231950 85140 0 0 $X=231700 $Y=84910
X7032 3 digital_ldo_top_VIA4 $T=231950 89220 0 0 $X=231700 $Y=88990
X7033 3 digital_ldo_top_VIA4 $T=231950 93300 0 0 $X=231700 $Y=93070
X7034 3 digital_ldo_top_VIA4 $T=231950 97380 0 0 $X=231700 $Y=97150
X7035 3 digital_ldo_top_VIA4 $T=231950 101460 0 0 $X=231700 $Y=101230
X7036 3 digital_ldo_top_VIA4 $T=231950 105540 0 0 $X=231700 $Y=105310
X7037 3 digital_ldo_top_VIA4 $T=231950 109620 0 0 $X=231700 $Y=109390
X7038 3 digital_ldo_top_VIA4 $T=231950 113700 0 0 $X=231700 $Y=113470
X7039 3 digital_ldo_top_VIA4 $T=231950 117780 0 0 $X=231700 $Y=117550
X7040 3 digital_ldo_top_VIA4 $T=231950 121860 0 0 $X=231700 $Y=121630
X7041 3 digital_ldo_top_VIA4 $T=231950 125940 0 0 $X=231700 $Y=125710
X7042 2 digital_ldo_top_VIA4 $T=233330 13060 0 0 $X=233080 $Y=12830
X7043 2 digital_ldo_top_VIA4 $T=233330 17140 0 0 $X=233080 $Y=16910
X7044 2 digital_ldo_top_VIA4 $T=233330 21220 0 0 $X=233080 $Y=20990
X7045 2 digital_ldo_top_VIA4 $T=233330 25300 0 0 $X=233080 $Y=25070
X7046 2 digital_ldo_top_VIA4 $T=233330 86500 0 0 $X=233080 $Y=86270
X7047 2 digital_ldo_top_VIA4 $T=233330 90580 0 0 $X=233080 $Y=90350
X7048 2 digital_ldo_top_VIA4 $T=233330 94660 0 0 $X=233080 $Y=94430
X7049 2 digital_ldo_top_VIA4 $T=233330 98740 0 0 $X=233080 $Y=98510
X7050 2 digital_ldo_top_VIA4 $T=233330 102820 0 0 $X=233080 $Y=102590
X7051 2 digital_ldo_top_VIA4 $T=233330 106900 0 0 $X=233080 $Y=106670
X7052 2 digital_ldo_top_VIA4 $T=233330 110980 0 0 $X=233080 $Y=110750
X7053 2 digital_ldo_top_VIA4 $T=233330 115060 0 0 $X=233080 $Y=114830
X7054 2 digital_ldo_top_VIA4 $T=233330 119140 0 0 $X=233080 $Y=118910
X7055 2 digital_ldo_top_VIA4 $T=233330 123220 0 0 $X=233080 $Y=122990
X7056 2 digital_ldo_top_VIA4 $T=233330 127300 0 0 $X=233080 $Y=127070
X7057 3 digital_ldo_top_VIA4 $T=235630 11700 0 0 $X=235380 $Y=11470
X7058 3 digital_ldo_top_VIA4 $T=235630 15780 0 0 $X=235380 $Y=15550
X7059 3 digital_ldo_top_VIA4 $T=235630 93300 0 0 $X=235380 $Y=93070
X7060 3 digital_ldo_top_VIA4 $T=235630 97380 0 0 $X=235380 $Y=97150
X7061 3 digital_ldo_top_VIA4 $T=235630 101460 0 0 $X=235380 $Y=101230
X7062 3 digital_ldo_top_VIA4 $T=235630 105540 0 0 $X=235380 $Y=105310
X7063 3 digital_ldo_top_VIA4 $T=235630 109620 0 0 $X=235380 $Y=109390
X7064 3 digital_ldo_top_VIA4 $T=235630 113700 0 0 $X=235380 $Y=113470
X7065 3 digital_ldo_top_VIA4 $T=235630 117780 0 0 $X=235380 $Y=117550
X7066 3 digital_ldo_top_VIA4 $T=235630 121860 0 0 $X=235380 $Y=121630
X7067 3 digital_ldo_top_VIA4 $T=235630 125940 0 0 $X=235380 $Y=125710
X7068 2 digital_ldo_top_VIA4 $T=237010 13060 0 0 $X=236760 $Y=12830
X7069 2 digital_ldo_top_VIA4 $T=237010 17140 0 0 $X=236760 $Y=16910
X7070 2 digital_ldo_top_VIA4 $T=237010 21220 0 0 $X=236760 $Y=20990
X7071 2 digital_ldo_top_VIA4 $T=237010 25300 0 0 $X=236760 $Y=25070
X7072 2 digital_ldo_top_VIA4 $T=237010 94660 0 0 $X=236760 $Y=94430
X7073 2 digital_ldo_top_VIA4 $T=237010 98740 0 0 $X=236760 $Y=98510
X7074 2 digital_ldo_top_VIA4 $T=237010 102820 0 0 $X=236760 $Y=102590
X7075 2 digital_ldo_top_VIA4 $T=237010 106900 0 0 $X=236760 $Y=106670
X7076 2 digital_ldo_top_VIA4 $T=237010 110980 0 0 $X=236760 $Y=110750
X7077 2 digital_ldo_top_VIA4 $T=237010 115060 0 0 $X=236760 $Y=114830
X7078 2 digital_ldo_top_VIA4 $T=237010 119140 0 0 $X=236760 $Y=118910
X7079 2 digital_ldo_top_VIA4 $T=237010 123220 0 0 $X=236760 $Y=122990
X7080 2 digital_ldo_top_VIA4 $T=237010 127300 0 0 $X=236760 $Y=127070
X7081 3 digital_ldo_top_VIA4 $T=239310 11700 0 0 $X=239060 $Y=11470
X7082 3 digital_ldo_top_VIA4 $T=239310 15780 0 0 $X=239060 $Y=15550
X7083 3 digital_ldo_top_VIA4 $T=239310 85140 0 0 $X=239060 $Y=84910
X7084 3 digital_ldo_top_VIA4 $T=239310 89220 0 0 $X=239060 $Y=88990
X7085 3 digital_ldo_top_VIA4 $T=239310 93300 0 0 $X=239060 $Y=93070
X7086 3 digital_ldo_top_VIA4 $T=239310 97380 0 0 $X=239060 $Y=97150
X7087 3 digital_ldo_top_VIA4 $T=239310 101460 0 0 $X=239060 $Y=101230
X7088 3 digital_ldo_top_VIA4 $T=239310 105540 0 0 $X=239060 $Y=105310
X7089 3 digital_ldo_top_VIA4 $T=239310 109620 0 0 $X=239060 $Y=109390
X7090 3 digital_ldo_top_VIA4 $T=239310 113700 0 0 $X=239060 $Y=113470
X7091 3 digital_ldo_top_VIA4 $T=239310 117780 0 0 $X=239060 $Y=117550
X7092 3 digital_ldo_top_VIA4 $T=239310 121860 0 0 $X=239060 $Y=121630
X7093 3 digital_ldo_top_VIA4 $T=239310 125940 0 0 $X=239060 $Y=125710
X7094 2 digital_ldo_top_VIA4 $T=240690 13060 0 0 $X=240440 $Y=12830
X7095 2 digital_ldo_top_VIA4 $T=240690 17140 0 0 $X=240440 $Y=16910
X7096 2 digital_ldo_top_VIA4 $T=240690 21220 0 0 $X=240440 $Y=20990
X7097 2 digital_ldo_top_VIA4 $T=240690 25300 0 0 $X=240440 $Y=25070
X7098 2 digital_ldo_top_VIA4 $T=240690 94660 0 0 $X=240440 $Y=94430
X7099 2 digital_ldo_top_VIA4 $T=240690 98740 0 0 $X=240440 $Y=98510
X7100 2 digital_ldo_top_VIA4 $T=240690 102820 0 0 $X=240440 $Y=102590
X7101 2 digital_ldo_top_VIA4 $T=240690 106900 0 0 $X=240440 $Y=106670
X7102 2 digital_ldo_top_VIA4 $T=240690 110980 0 0 $X=240440 $Y=110750
X7103 2 digital_ldo_top_VIA4 $T=240690 115060 0 0 $X=240440 $Y=114830
X7104 2 digital_ldo_top_VIA4 $T=240690 119140 0 0 $X=240440 $Y=118910
X7105 2 digital_ldo_top_VIA4 $T=240690 123220 0 0 $X=240440 $Y=122990
X7106 2 digital_ldo_top_VIA4 $T=240690 127300 0 0 $X=240440 $Y=127070
X7107 3 digital_ldo_top_VIA4 $T=242990 11700 0 0 $X=242740 $Y=11470
X7108 3 digital_ldo_top_VIA4 $T=242990 15780 0 0 $X=242740 $Y=15550
X7109 3 digital_ldo_top_VIA4 $T=242990 19860 0 0 $X=242740 $Y=19630
X7110 3 digital_ldo_top_VIA4 $T=242990 23940 0 0 $X=242740 $Y=23710
X7111 3 digital_ldo_top_VIA4 $T=242990 32100 0 0 $X=242740 $Y=31870
X7112 3 digital_ldo_top_VIA4 $T=242990 85140 0 0 $X=242740 $Y=84910
X7113 3 digital_ldo_top_VIA4 $T=242990 89220 0 0 $X=242740 $Y=88990
X7114 3 digital_ldo_top_VIA4 $T=242990 93300 0 0 $X=242740 $Y=93070
X7115 3 digital_ldo_top_VIA4 $T=242990 97380 0 0 $X=242740 $Y=97150
X7116 3 digital_ldo_top_VIA4 $T=242990 101460 0 0 $X=242740 $Y=101230
X7117 3 digital_ldo_top_VIA4 $T=242990 105540 0 0 $X=242740 $Y=105310
X7118 3 digital_ldo_top_VIA4 $T=242990 109620 0 0 $X=242740 $Y=109390
X7119 3 digital_ldo_top_VIA4 $T=242990 113700 0 0 $X=242740 $Y=113470
X7120 3 digital_ldo_top_VIA4 $T=242990 117780 0 0 $X=242740 $Y=117550
X7121 3 digital_ldo_top_VIA4 $T=242990 121860 0 0 $X=242740 $Y=121630
X7122 3 digital_ldo_top_VIA4 $T=242990 125940 0 0 $X=242740 $Y=125710
X7123 2 digital_ldo_top_VIA4 $T=244370 13060 0 0 $X=244120 $Y=12830
X7124 2 digital_ldo_top_VIA4 $T=244370 17140 0 0 $X=244120 $Y=16910
X7125 2 digital_ldo_top_VIA4 $T=244370 21220 0 0 $X=244120 $Y=20990
X7126 2 digital_ldo_top_VIA4 $T=244370 25300 0 0 $X=244120 $Y=25070
X7127 2 digital_ldo_top_VIA4 $T=244370 86500 0 0 $X=244120 $Y=86270
X7128 2 digital_ldo_top_VIA4 $T=244370 90580 0 0 $X=244120 $Y=90350
X7129 2 digital_ldo_top_VIA4 $T=244370 94660 0 0 $X=244120 $Y=94430
X7130 2 digital_ldo_top_VIA4 $T=244370 98740 0 0 $X=244120 $Y=98510
X7131 2 digital_ldo_top_VIA4 $T=244370 102820 0 0 $X=244120 $Y=102590
X7132 2 digital_ldo_top_VIA4 $T=244370 106900 0 0 $X=244120 $Y=106670
X7133 2 digital_ldo_top_VIA4 $T=244370 110980 0 0 $X=244120 $Y=110750
X7134 2 digital_ldo_top_VIA4 $T=244370 115060 0 0 $X=244120 $Y=114830
X7135 2 digital_ldo_top_VIA4 $T=244370 119140 0 0 $X=244120 $Y=118910
X7136 2 digital_ldo_top_VIA4 $T=244370 123220 0 0 $X=244120 $Y=122990
X7137 2 digital_ldo_top_VIA4 $T=244370 127300 0 0 $X=244120 $Y=127070
X7138 3 digital_ldo_top_VIA4 $T=246670 11700 0 0 $X=246420 $Y=11470
X7139 3 digital_ldo_top_VIA4 $T=246670 15780 0 0 $X=246420 $Y=15550
X7140 3 digital_ldo_top_VIA4 $T=246670 93300 0 0 $X=246420 $Y=93070
X7141 3 digital_ldo_top_VIA4 $T=246670 97380 0 0 $X=246420 $Y=97150
X7142 3 digital_ldo_top_VIA4 $T=246670 101460 0 0 $X=246420 $Y=101230
X7143 3 digital_ldo_top_VIA4 $T=246670 105540 0 0 $X=246420 $Y=105310
X7144 3 digital_ldo_top_VIA4 $T=246670 109620 0 0 $X=246420 $Y=109390
X7145 3 digital_ldo_top_VIA4 $T=246670 113700 0 0 $X=246420 $Y=113470
X7146 3 digital_ldo_top_VIA4 $T=246670 117780 0 0 $X=246420 $Y=117550
X7147 3 digital_ldo_top_VIA4 $T=246670 121860 0 0 $X=246420 $Y=121630
X7148 3 digital_ldo_top_VIA4 $T=246670 125940 0 0 $X=246420 $Y=125710
X7149 2 digital_ldo_top_VIA4 $T=248050 13060 0 0 $X=247800 $Y=12830
X7150 2 digital_ldo_top_VIA4 $T=248050 17140 0 0 $X=247800 $Y=16910
X7151 2 digital_ldo_top_VIA4 $T=248050 94660 0 0 $X=247800 $Y=94430
X7152 2 digital_ldo_top_VIA4 $T=248050 98740 0 0 $X=247800 $Y=98510
X7153 2 digital_ldo_top_VIA4 $T=248050 102820 0 0 $X=247800 $Y=102590
X7154 2 digital_ldo_top_VIA4 $T=248050 106900 0 0 $X=247800 $Y=106670
X7155 2 digital_ldo_top_VIA4 $T=248050 110980 0 0 $X=247800 $Y=110750
X7156 2 digital_ldo_top_VIA4 $T=248050 115060 0 0 $X=247800 $Y=114830
X7157 2 digital_ldo_top_VIA4 $T=248050 119140 0 0 $X=247800 $Y=118910
X7158 2 digital_ldo_top_VIA4 $T=248050 123220 0 0 $X=247800 $Y=122990
X7159 2 digital_ldo_top_VIA4 $T=248050 127300 0 0 $X=247800 $Y=127070
X7160 3 digital_ldo_top_VIA4 $T=250350 11700 0 0 $X=250100 $Y=11470
X7161 3 digital_ldo_top_VIA4 $T=250350 15780 0 0 $X=250100 $Y=15550
X7162 3 digital_ldo_top_VIA4 $T=250350 19860 0 0 $X=250100 $Y=19630
X7163 3 digital_ldo_top_VIA4 $T=250350 23940 0 0 $X=250100 $Y=23710
X7164 3 digital_ldo_top_VIA4 $T=250350 32100 0 0 $X=250100 $Y=31870
X7165 3 digital_ldo_top_VIA4 $T=250350 85140 0 0 $X=250100 $Y=84910
X7166 3 digital_ldo_top_VIA4 $T=250350 89220 0 0 $X=250100 $Y=88990
X7167 3 digital_ldo_top_VIA4 $T=250350 93300 0 0 $X=250100 $Y=93070
X7168 3 digital_ldo_top_VIA4 $T=250350 97380 0 0 $X=250100 $Y=97150
X7169 3 digital_ldo_top_VIA4 $T=250350 101460 0 0 $X=250100 $Y=101230
X7170 3 digital_ldo_top_VIA4 $T=250350 105540 0 0 $X=250100 $Y=105310
X7171 3 digital_ldo_top_VIA4 $T=250350 109620 0 0 $X=250100 $Y=109390
X7172 3 digital_ldo_top_VIA4 $T=250350 113700 0 0 $X=250100 $Y=113470
X7173 3 digital_ldo_top_VIA4 $T=250350 117780 0 0 $X=250100 $Y=117550
X7174 3 digital_ldo_top_VIA4 $T=250350 121860 0 0 $X=250100 $Y=121630
X7175 3 digital_ldo_top_VIA4 $T=250350 125940 0 0 $X=250100 $Y=125710
X7176 2 digital_ldo_top_VIA4 $T=251730 13060 0 0 $X=251480 $Y=12830
X7177 2 digital_ldo_top_VIA4 $T=251730 17140 0 0 $X=251480 $Y=16910
X7178 2 digital_ldo_top_VIA4 $T=251730 21220 0 0 $X=251480 $Y=20990
X7179 2 digital_ldo_top_VIA4 $T=251730 25300 0 0 $X=251480 $Y=25070
X7180 2 digital_ldo_top_VIA4 $T=251730 94660 0 0 $X=251480 $Y=94430
X7181 2 digital_ldo_top_VIA4 $T=251730 98740 0 0 $X=251480 $Y=98510
X7182 2 digital_ldo_top_VIA4 $T=251730 102820 0 0 $X=251480 $Y=102590
X7183 2 digital_ldo_top_VIA4 $T=251730 106900 0 0 $X=251480 $Y=106670
X7184 2 digital_ldo_top_VIA4 $T=251730 110980 0 0 $X=251480 $Y=110750
X7185 2 digital_ldo_top_VIA4 $T=251730 115060 0 0 $X=251480 $Y=114830
X7186 2 digital_ldo_top_VIA4 $T=251730 119140 0 0 $X=251480 $Y=118910
X7187 2 digital_ldo_top_VIA4 $T=251730 123220 0 0 $X=251480 $Y=122990
X7188 2 digital_ldo_top_VIA4 $T=251730 127300 0 0 $X=251480 $Y=127070
X7189 3 digital_ldo_top_VIA4 $T=254030 11700 0 0 $X=253780 $Y=11470
X7190 3 digital_ldo_top_VIA4 $T=254030 15780 0 0 $X=253780 $Y=15550
X7191 3 digital_ldo_top_VIA4 $T=254030 19860 0 0 $X=253780 $Y=19630
X7192 3 digital_ldo_top_VIA4 $T=254030 23940 0 0 $X=253780 $Y=23710
X7193 3 digital_ldo_top_VIA4 $T=254030 32100 0 0 $X=253780 $Y=31870
X7194 3 digital_ldo_top_VIA4 $T=254030 85140 0 0 $X=253780 $Y=84910
X7195 3 digital_ldo_top_VIA4 $T=254030 89220 0 0 $X=253780 $Y=88990
X7196 3 digital_ldo_top_VIA4 $T=254030 93300 0 0 $X=253780 $Y=93070
X7197 3 digital_ldo_top_VIA4 $T=254030 97380 0 0 $X=253780 $Y=97150
X7198 3 digital_ldo_top_VIA4 $T=254030 101460 0 0 $X=253780 $Y=101230
X7199 3 digital_ldo_top_VIA4 $T=254030 105540 0 0 $X=253780 $Y=105310
X7200 3 digital_ldo_top_VIA4 $T=254030 109620 0 0 $X=253780 $Y=109390
X7201 3 digital_ldo_top_VIA4 $T=254030 113700 0 0 $X=253780 $Y=113470
X7202 3 digital_ldo_top_VIA4 $T=254030 117780 0 0 $X=253780 $Y=117550
X7203 3 digital_ldo_top_VIA4 $T=254030 121860 0 0 $X=253780 $Y=121630
X7204 3 digital_ldo_top_VIA4 $T=254030 125940 0 0 $X=253780 $Y=125710
X7205 2 digital_ldo_top_VIA4 $T=255410 13060 0 0 $X=255160 $Y=12830
X7206 2 digital_ldo_top_VIA4 $T=255410 17140 0 0 $X=255160 $Y=16910
X7207 2 digital_ldo_top_VIA4 $T=255410 86500 0 0 $X=255160 $Y=86270
X7208 2 digital_ldo_top_VIA4 $T=255410 90580 0 0 $X=255160 $Y=90350
X7209 2 digital_ldo_top_VIA4 $T=255410 94660 0 0 $X=255160 $Y=94430
X7210 2 digital_ldo_top_VIA4 $T=255410 98740 0 0 $X=255160 $Y=98510
X7211 2 digital_ldo_top_VIA4 $T=255410 102820 0 0 $X=255160 $Y=102590
X7212 2 digital_ldo_top_VIA4 $T=255410 106900 0 0 $X=255160 $Y=106670
X7213 2 digital_ldo_top_VIA4 $T=255410 110980 0 0 $X=255160 $Y=110750
X7214 2 digital_ldo_top_VIA4 $T=255410 115060 0 0 $X=255160 $Y=114830
X7215 2 digital_ldo_top_VIA4 $T=255410 119140 0 0 $X=255160 $Y=118910
X7216 2 digital_ldo_top_VIA4 $T=255410 123220 0 0 $X=255160 $Y=122990
X7217 2 digital_ldo_top_VIA4 $T=255410 127300 0 0 $X=255160 $Y=127070
X7218 3 digital_ldo_top_VIA4 $T=257710 11700 0 0 $X=257460 $Y=11470
X7219 3 digital_ldo_top_VIA4 $T=257710 15780 0 0 $X=257460 $Y=15550
X7220 3 digital_ldo_top_VIA4 $T=257710 93300 0 0 $X=257460 $Y=93070
X7221 3 digital_ldo_top_VIA4 $T=257710 97380 0 0 $X=257460 $Y=97150
X7222 3 digital_ldo_top_VIA4 $T=257710 101460 0 0 $X=257460 $Y=101230
X7223 3 digital_ldo_top_VIA4 $T=257710 105540 0 0 $X=257460 $Y=105310
X7224 3 digital_ldo_top_VIA4 $T=257710 109620 0 0 $X=257460 $Y=109390
X7225 3 digital_ldo_top_VIA4 $T=257710 113700 0 0 $X=257460 $Y=113470
X7226 3 digital_ldo_top_VIA4 $T=257710 117780 0 0 $X=257460 $Y=117550
X7227 3 digital_ldo_top_VIA4 $T=257710 121860 0 0 $X=257460 $Y=121630
X7228 3 digital_ldo_top_VIA4 $T=257710 125940 0 0 $X=257460 $Y=125710
X7229 2 digital_ldo_top_VIA4 $T=259090 13060 0 0 $X=258840 $Y=12830
X7230 2 digital_ldo_top_VIA4 $T=259090 17140 0 0 $X=258840 $Y=16910
X7231 2 digital_ldo_top_VIA4 $T=259090 94660 0 0 $X=258840 $Y=94430
X7232 2 digital_ldo_top_VIA4 $T=259090 98740 0 0 $X=258840 $Y=98510
X7233 2 digital_ldo_top_VIA4 $T=259090 102820 0 0 $X=258840 $Y=102590
X7234 2 digital_ldo_top_VIA4 $T=259090 106900 0 0 $X=258840 $Y=106670
X7235 2 digital_ldo_top_VIA4 $T=259090 110980 0 0 $X=258840 $Y=110750
X7236 2 digital_ldo_top_VIA4 $T=259090 115060 0 0 $X=258840 $Y=114830
X7237 2 digital_ldo_top_VIA4 $T=259090 119140 0 0 $X=258840 $Y=118910
X7238 2 digital_ldo_top_VIA4 $T=259090 123220 0 0 $X=258840 $Y=122990
X7239 2 digital_ldo_top_VIA4 $T=259090 127300 0 0 $X=258840 $Y=127070
X7240 3 digital_ldo_top_VIA4 $T=261390 11700 0 0 $X=261140 $Y=11470
X7241 3 digital_ldo_top_VIA4 $T=261390 15780 0 0 $X=261140 $Y=15550
X7242 3 digital_ldo_top_VIA4 $T=261390 19860 0 0 $X=261140 $Y=19630
X7243 3 digital_ldo_top_VIA4 $T=261390 23940 0 0 $X=261140 $Y=23710
X7244 3 digital_ldo_top_VIA4 $T=261390 32100 0 0 $X=261140 $Y=31870
X7245 3 digital_ldo_top_VIA4 $T=261390 85140 0 0 $X=261140 $Y=84910
X7246 3 digital_ldo_top_VIA4 $T=261390 89220 0 0 $X=261140 $Y=88990
X7247 3 digital_ldo_top_VIA4 $T=261390 93300 0 0 $X=261140 $Y=93070
X7248 3 digital_ldo_top_VIA4 $T=261390 97380 0 0 $X=261140 $Y=97150
X7249 3 digital_ldo_top_VIA4 $T=261390 101460 0 0 $X=261140 $Y=101230
X7250 3 digital_ldo_top_VIA4 $T=261390 105540 0 0 $X=261140 $Y=105310
X7251 3 digital_ldo_top_VIA4 $T=261390 109620 0 0 $X=261140 $Y=109390
X7252 3 digital_ldo_top_VIA4 $T=261390 113700 0 0 $X=261140 $Y=113470
X7253 3 digital_ldo_top_VIA4 $T=261390 117780 0 0 $X=261140 $Y=117550
X7254 3 digital_ldo_top_VIA4 $T=261390 121860 0 0 $X=261140 $Y=121630
X7255 3 digital_ldo_top_VIA4 $T=261390 125940 0 0 $X=261140 $Y=125710
X7256 2 digital_ldo_top_VIA4 $T=262770 13060 0 0 $X=262520 $Y=12830
X7257 2 digital_ldo_top_VIA4 $T=262770 17140 0 0 $X=262520 $Y=16910
X7258 2 digital_ldo_top_VIA4 $T=262770 21220 0 0 $X=262520 $Y=20990
X7259 2 digital_ldo_top_VIA4 $T=262770 25300 0 0 $X=262520 $Y=25070
X7260 2 digital_ldo_top_VIA4 $T=262770 94660 0 0 $X=262520 $Y=94430
X7261 2 digital_ldo_top_VIA4 $T=262770 98740 0 0 $X=262520 $Y=98510
X7262 2 digital_ldo_top_VIA4 $T=262770 102820 0 0 $X=262520 $Y=102590
X7263 2 digital_ldo_top_VIA4 $T=262770 106900 0 0 $X=262520 $Y=106670
X7264 2 digital_ldo_top_VIA4 $T=262770 110980 0 0 $X=262520 $Y=110750
X7265 2 digital_ldo_top_VIA4 $T=262770 115060 0 0 $X=262520 $Y=114830
X7266 2 digital_ldo_top_VIA4 $T=262770 119140 0 0 $X=262520 $Y=118910
X7267 2 digital_ldo_top_VIA4 $T=262770 123220 0 0 $X=262520 $Y=122990
X7268 2 digital_ldo_top_VIA4 $T=262770 127300 0 0 $X=262520 $Y=127070
X7269 3 digital_ldo_top_VIA4 $T=265070 11700 0 0 $X=264820 $Y=11470
X7270 3 digital_ldo_top_VIA4 $T=265070 15780 0 0 $X=264820 $Y=15550
X7271 3 digital_ldo_top_VIA4 $T=265070 19860 0 0 $X=264820 $Y=19630
X7272 3 digital_ldo_top_VIA4 $T=265070 23940 0 0 $X=264820 $Y=23710
X7273 3 digital_ldo_top_VIA4 $T=265070 32100 0 0 $X=264820 $Y=31870
X7274 3 digital_ldo_top_VIA4 $T=265070 85140 0 0 $X=264820 $Y=84910
X7275 3 digital_ldo_top_VIA4 $T=265070 89220 0 0 $X=264820 $Y=88990
X7276 3 digital_ldo_top_VIA4 $T=265070 93300 0 0 $X=264820 $Y=93070
X7277 3 digital_ldo_top_VIA4 $T=265070 97380 0 0 $X=264820 $Y=97150
X7278 3 digital_ldo_top_VIA4 $T=265070 101460 0 0 $X=264820 $Y=101230
X7279 3 digital_ldo_top_VIA4 $T=265070 105540 0 0 $X=264820 $Y=105310
X7280 3 digital_ldo_top_VIA4 $T=265070 109620 0 0 $X=264820 $Y=109390
X7281 3 digital_ldo_top_VIA4 $T=265070 113700 0 0 $X=264820 $Y=113470
X7282 3 digital_ldo_top_VIA4 $T=265070 117780 0 0 $X=264820 $Y=117550
X7283 3 digital_ldo_top_VIA4 $T=265070 121860 0 0 $X=264820 $Y=121630
X7284 3 digital_ldo_top_VIA4 $T=265070 125940 0 0 $X=264820 $Y=125710
X7285 2 digital_ldo_top_VIA4 $T=266450 13060 0 0 $X=266200 $Y=12830
X7286 2 digital_ldo_top_VIA4 $T=266450 17140 0 0 $X=266200 $Y=16910
X7287 2 digital_ldo_top_VIA4 $T=266450 86500 0 0 $X=266200 $Y=86270
X7288 2 digital_ldo_top_VIA4 $T=266450 90580 0 0 $X=266200 $Y=90350
X7289 2 digital_ldo_top_VIA4 $T=266450 94660 0 0 $X=266200 $Y=94430
X7290 2 digital_ldo_top_VIA4 $T=266450 98740 0 0 $X=266200 $Y=98510
X7291 2 digital_ldo_top_VIA4 $T=266450 102820 0 0 $X=266200 $Y=102590
X7292 2 digital_ldo_top_VIA4 $T=266450 106900 0 0 $X=266200 $Y=106670
X7293 2 digital_ldo_top_VIA4 $T=266450 110980 0 0 $X=266200 $Y=110750
X7294 2 digital_ldo_top_VIA4 $T=266450 115060 0 0 $X=266200 $Y=114830
X7295 2 digital_ldo_top_VIA4 $T=266450 119140 0 0 $X=266200 $Y=118910
X7296 2 digital_ldo_top_VIA4 $T=266450 123220 0 0 $X=266200 $Y=122990
X7297 2 digital_ldo_top_VIA4 $T=266450 127300 0 0 $X=266200 $Y=127070
X7298 3 digital_ldo_top_VIA4 $T=268750 11700 0 0 $X=268500 $Y=11470
X7299 3 digital_ldo_top_VIA4 $T=268750 15780 0 0 $X=268500 $Y=15550
X7300 3 digital_ldo_top_VIA4 $T=268750 93300 0 0 $X=268500 $Y=93070
X7301 3 digital_ldo_top_VIA4 $T=268750 97380 0 0 $X=268500 $Y=97150
X7302 3 digital_ldo_top_VIA4 $T=268750 101460 0 0 $X=268500 $Y=101230
X7303 3 digital_ldo_top_VIA4 $T=268750 105540 0 0 $X=268500 $Y=105310
X7304 3 digital_ldo_top_VIA4 $T=268750 109620 0 0 $X=268500 $Y=109390
X7305 3 digital_ldo_top_VIA4 $T=268750 113700 0 0 $X=268500 $Y=113470
X7306 3 digital_ldo_top_VIA4 $T=268750 117780 0 0 $X=268500 $Y=117550
X7307 3 digital_ldo_top_VIA4 $T=268750 121860 0 0 $X=268500 $Y=121630
X7308 3 digital_ldo_top_VIA4 $T=268750 125940 0 0 $X=268500 $Y=125710
X7309 2 digital_ldo_top_VIA4 $T=270130 13060 0 0 $X=269880 $Y=12830
X7310 2 digital_ldo_top_VIA4 $T=270130 17140 0 0 $X=269880 $Y=16910
X7311 2 digital_ldo_top_VIA4 $T=270130 94660 0 0 $X=269880 $Y=94430
X7312 2 digital_ldo_top_VIA4 $T=270130 98740 0 0 $X=269880 $Y=98510
X7313 2 digital_ldo_top_VIA4 $T=270130 102820 0 0 $X=269880 $Y=102590
X7314 2 digital_ldo_top_VIA4 $T=270130 106900 0 0 $X=269880 $Y=106670
X7315 2 digital_ldo_top_VIA4 $T=270130 110980 0 0 $X=269880 $Y=110750
X7316 2 digital_ldo_top_VIA4 $T=270130 115060 0 0 $X=269880 $Y=114830
X7317 2 digital_ldo_top_VIA4 $T=270130 119140 0 0 $X=269880 $Y=118910
X7318 2 digital_ldo_top_VIA4 $T=270130 123220 0 0 $X=269880 $Y=122990
X7319 2 digital_ldo_top_VIA4 $T=270130 127300 0 0 $X=269880 $Y=127070
X7320 3 digital_ldo_top_VIA4 $T=272430 11700 0 0 $X=272180 $Y=11470
X7321 3 digital_ldo_top_VIA4 $T=272430 15780 0 0 $X=272180 $Y=15550
X7322 3 digital_ldo_top_VIA4 $T=272430 85140 0 0 $X=272180 $Y=84910
X7323 3 digital_ldo_top_VIA4 $T=272430 89220 0 0 $X=272180 $Y=88990
X7324 3 digital_ldo_top_VIA4 $T=272430 93300 0 0 $X=272180 $Y=93070
X7325 3 digital_ldo_top_VIA4 $T=272430 97380 0 0 $X=272180 $Y=97150
X7326 3 digital_ldo_top_VIA4 $T=272430 101460 0 0 $X=272180 $Y=101230
X7327 3 digital_ldo_top_VIA4 $T=272430 105540 0 0 $X=272180 $Y=105310
X7328 3 digital_ldo_top_VIA4 $T=272430 109620 0 0 $X=272180 $Y=109390
X7329 3 digital_ldo_top_VIA4 $T=272430 113700 0 0 $X=272180 $Y=113470
X7330 3 digital_ldo_top_VIA4 $T=272430 117780 0 0 $X=272180 $Y=117550
X7331 3 digital_ldo_top_VIA4 $T=272430 121860 0 0 $X=272180 $Y=121630
X7332 3 digital_ldo_top_VIA4 $T=272430 125940 0 0 $X=272180 $Y=125710
X7333 2 digital_ldo_top_VIA4 $T=273810 13060 0 0 $X=273560 $Y=12830
X7334 2 digital_ldo_top_VIA4 $T=273810 17140 0 0 $X=273560 $Y=16910
X7335 2 digital_ldo_top_VIA4 $T=273810 21220 0 0 $X=273560 $Y=20990
X7336 2 digital_ldo_top_VIA4 $T=273810 25300 0 0 $X=273560 $Y=25070
X7337 2 digital_ldo_top_VIA4 $T=273810 94660 0 0 $X=273560 $Y=94430
X7338 2 digital_ldo_top_VIA4 $T=273810 98740 0 0 $X=273560 $Y=98510
X7339 2 digital_ldo_top_VIA4 $T=273810 102820 0 0 $X=273560 $Y=102590
X7340 2 digital_ldo_top_VIA4 $T=273810 106900 0 0 $X=273560 $Y=106670
X7341 2 digital_ldo_top_VIA4 $T=273810 110980 0 0 $X=273560 $Y=110750
X7342 2 digital_ldo_top_VIA4 $T=273810 115060 0 0 $X=273560 $Y=114830
X7343 2 digital_ldo_top_VIA4 $T=273810 119140 0 0 $X=273560 $Y=118910
X7344 2 digital_ldo_top_VIA4 $T=273810 123220 0 0 $X=273560 $Y=122990
X7345 2 digital_ldo_top_VIA4 $T=273810 127300 0 0 $X=273560 $Y=127070
X7346 3 digital_ldo_top_VIA4 $T=276110 11700 0 0 $X=275860 $Y=11470
X7347 3 digital_ldo_top_VIA4 $T=276110 15780 0 0 $X=275860 $Y=15550
X7348 3 digital_ldo_top_VIA4 $T=276110 85140 0 0 $X=275860 $Y=84910
X7349 3 digital_ldo_top_VIA4 $T=276110 89220 0 0 $X=275860 $Y=88990
X7350 3 digital_ldo_top_VIA4 $T=276110 93300 0 0 $X=275860 $Y=93070
X7351 3 digital_ldo_top_VIA4 $T=276110 97380 0 0 $X=275860 $Y=97150
X7352 3 digital_ldo_top_VIA4 $T=276110 101460 0 0 $X=275860 $Y=101230
X7353 3 digital_ldo_top_VIA4 $T=276110 105540 0 0 $X=275860 $Y=105310
X7354 3 digital_ldo_top_VIA4 $T=276110 109620 0 0 $X=275860 $Y=109390
X7355 3 digital_ldo_top_VIA4 $T=276110 113700 0 0 $X=275860 $Y=113470
X7356 3 digital_ldo_top_VIA4 $T=276110 117780 0 0 $X=275860 $Y=117550
X7357 3 digital_ldo_top_VIA4 $T=276110 121860 0 0 $X=275860 $Y=121630
X7358 3 digital_ldo_top_VIA4 $T=276110 125940 0 0 $X=275860 $Y=125710
X7359 2 digital_ldo_top_VIA4 $T=277490 13060 0 0 $X=277240 $Y=12830
X7360 2 digital_ldo_top_VIA4 $T=277490 17140 0 0 $X=277240 $Y=16910
X7361 2 digital_ldo_top_VIA4 $T=277490 21220 0 0 $X=277240 $Y=20990
X7362 2 digital_ldo_top_VIA4 $T=277490 25300 0 0 $X=277240 $Y=25070
X7363 2 digital_ldo_top_VIA4 $T=277490 86500 0 0 $X=277240 $Y=86270
X7364 2 digital_ldo_top_VIA4 $T=277490 90580 0 0 $X=277240 $Y=90350
X7365 2 digital_ldo_top_VIA4 $T=277490 94660 0 0 $X=277240 $Y=94430
X7366 2 digital_ldo_top_VIA4 $T=277490 98740 0 0 $X=277240 $Y=98510
X7367 2 digital_ldo_top_VIA4 $T=277490 102820 0 0 $X=277240 $Y=102590
X7368 2 digital_ldo_top_VIA4 $T=277490 106900 0 0 $X=277240 $Y=106670
X7369 2 digital_ldo_top_VIA4 $T=277490 110980 0 0 $X=277240 $Y=110750
X7370 2 digital_ldo_top_VIA4 $T=277490 115060 0 0 $X=277240 $Y=114830
X7371 2 digital_ldo_top_VIA4 $T=277490 119140 0 0 $X=277240 $Y=118910
X7372 2 digital_ldo_top_VIA4 $T=277490 123220 0 0 $X=277240 $Y=122990
X7373 2 digital_ldo_top_VIA4 $T=277490 127300 0 0 $X=277240 $Y=127070
X7374 3 digital_ldo_top_VIA4 $T=279790 11700 0 0 $X=279540 $Y=11470
X7375 3 digital_ldo_top_VIA4 $T=279790 15780 0 0 $X=279540 $Y=15550
X7376 3 digital_ldo_top_VIA4 $T=279790 93300 0 0 $X=279540 $Y=93070
X7377 3 digital_ldo_top_VIA4 $T=279790 97380 0 0 $X=279540 $Y=97150
X7378 3 digital_ldo_top_VIA4 $T=279790 101460 0 0 $X=279540 $Y=101230
X7379 3 digital_ldo_top_VIA4 $T=279790 105540 0 0 $X=279540 $Y=105310
X7380 3 digital_ldo_top_VIA4 $T=279790 109620 0 0 $X=279540 $Y=109390
X7381 3 digital_ldo_top_VIA4 $T=279790 113700 0 0 $X=279540 $Y=113470
X7382 3 digital_ldo_top_VIA4 $T=279790 117780 0 0 $X=279540 $Y=117550
X7383 3 digital_ldo_top_VIA4 $T=279790 121860 0 0 $X=279540 $Y=121630
X7384 3 digital_ldo_top_VIA4 $T=279790 125940 0 0 $X=279540 $Y=125710
X7385 2 digital_ldo_top_VIA4 $T=281170 13060 0 0 $X=280920 $Y=12830
X7386 2 digital_ldo_top_VIA4 $T=281170 17140 0 0 $X=280920 $Y=16910
X7387 2 digital_ldo_top_VIA4 $T=281170 21220 0 0 $X=280920 $Y=20990
X7388 2 digital_ldo_top_VIA4 $T=281170 25300 0 0 $X=280920 $Y=25070
X7389 2 digital_ldo_top_VIA4 $T=281170 94660 0 0 $X=280920 $Y=94430
X7390 2 digital_ldo_top_VIA4 $T=281170 98740 0 0 $X=280920 $Y=98510
X7391 2 digital_ldo_top_VIA4 $T=281170 102820 0 0 $X=280920 $Y=102590
X7392 2 digital_ldo_top_VIA4 $T=281170 106900 0 0 $X=280920 $Y=106670
X7393 2 digital_ldo_top_VIA4 $T=281170 110980 0 0 $X=280920 $Y=110750
X7394 2 digital_ldo_top_VIA4 $T=281170 115060 0 0 $X=280920 $Y=114830
X7395 2 digital_ldo_top_VIA4 $T=281170 119140 0 0 $X=280920 $Y=118910
X7396 2 digital_ldo_top_VIA4 $T=281170 123220 0 0 $X=280920 $Y=122990
X7397 2 digital_ldo_top_VIA4 $T=281170 127300 0 0 $X=280920 $Y=127070
X7398 3 digital_ldo_top_VIA4 $T=283470 11700 0 0 $X=283220 $Y=11470
X7399 3 digital_ldo_top_VIA4 $T=283470 15780 0 0 $X=283220 $Y=15550
X7400 3 digital_ldo_top_VIA4 $T=283470 85140 0 0 $X=283220 $Y=84910
X7401 3 digital_ldo_top_VIA4 $T=283470 89220 0 0 $X=283220 $Y=88990
X7402 3 digital_ldo_top_VIA4 $T=283470 93300 0 0 $X=283220 $Y=93070
X7403 3 digital_ldo_top_VIA4 $T=283470 97380 0 0 $X=283220 $Y=97150
X7404 3 digital_ldo_top_VIA4 $T=283470 101460 0 0 $X=283220 $Y=101230
X7405 3 digital_ldo_top_VIA4 $T=283470 105540 0 0 $X=283220 $Y=105310
X7406 3 digital_ldo_top_VIA4 $T=283470 109620 0 0 $X=283220 $Y=109390
X7407 3 digital_ldo_top_VIA4 $T=283470 113700 0 0 $X=283220 $Y=113470
X7408 3 digital_ldo_top_VIA4 $T=283470 117780 0 0 $X=283220 $Y=117550
X7409 3 digital_ldo_top_VIA4 $T=283470 121860 0 0 $X=283220 $Y=121630
X7410 3 digital_ldo_top_VIA4 $T=283470 125940 0 0 $X=283220 $Y=125710
X7411 2 digital_ldo_top_VIA4 $T=284850 13060 0 0 $X=284600 $Y=12830
X7412 2 digital_ldo_top_VIA4 $T=284850 17140 0 0 $X=284600 $Y=16910
X7413 2 digital_ldo_top_VIA4 $T=284850 21220 0 0 $X=284600 $Y=20990
X7414 2 digital_ldo_top_VIA4 $T=284850 25300 0 0 $X=284600 $Y=25070
X7415 2 digital_ldo_top_VIA4 $T=284850 94660 0 0 $X=284600 $Y=94430
X7416 2 digital_ldo_top_VIA4 $T=284850 98740 0 0 $X=284600 $Y=98510
X7417 2 digital_ldo_top_VIA4 $T=284850 102820 0 0 $X=284600 $Y=102590
X7418 2 digital_ldo_top_VIA4 $T=284850 106900 0 0 $X=284600 $Y=106670
X7419 2 digital_ldo_top_VIA4 $T=284850 110980 0 0 $X=284600 $Y=110750
X7420 2 digital_ldo_top_VIA4 $T=284850 115060 0 0 $X=284600 $Y=114830
X7421 2 digital_ldo_top_VIA4 $T=284850 119140 0 0 $X=284600 $Y=118910
X7422 2 digital_ldo_top_VIA4 $T=284850 123220 0 0 $X=284600 $Y=122990
X7423 2 digital_ldo_top_VIA4 $T=284850 127300 0 0 $X=284600 $Y=127070
X7424 3 digital_ldo_top_VIA4 $T=287150 11700 0 0 $X=286900 $Y=11470
X7425 3 digital_ldo_top_VIA4 $T=287150 15780 0 0 $X=286900 $Y=15550
X7426 3 digital_ldo_top_VIA4 $T=287150 19860 0 0 $X=286900 $Y=19630
X7427 3 digital_ldo_top_VIA4 $T=287150 23940 0 0 $X=286900 $Y=23710
X7428 3 digital_ldo_top_VIA4 $T=287150 32100 0 0 $X=286900 $Y=31870
X7429 3 digital_ldo_top_VIA4 $T=287150 85140 0 0 $X=286900 $Y=84910
X7430 3 digital_ldo_top_VIA4 $T=287150 89220 0 0 $X=286900 $Y=88990
X7431 3 digital_ldo_top_VIA4 $T=287150 93300 0 0 $X=286900 $Y=93070
X7432 3 digital_ldo_top_VIA4 $T=287150 97380 0 0 $X=286900 $Y=97150
X7433 3 digital_ldo_top_VIA4 $T=287150 101460 0 0 $X=286900 $Y=101230
X7434 3 digital_ldo_top_VIA4 $T=287150 105540 0 0 $X=286900 $Y=105310
X7435 3 digital_ldo_top_VIA4 $T=287150 109620 0 0 $X=286900 $Y=109390
X7436 3 digital_ldo_top_VIA4 $T=287150 113700 0 0 $X=286900 $Y=113470
X7437 3 digital_ldo_top_VIA4 $T=287150 117780 0 0 $X=286900 $Y=117550
X7438 3 digital_ldo_top_VIA4 $T=287150 121860 0 0 $X=286900 $Y=121630
X7439 3 digital_ldo_top_VIA4 $T=287150 125940 0 0 $X=286900 $Y=125710
X7440 2 digital_ldo_top_VIA4 $T=288530 13060 0 0 $X=288280 $Y=12830
X7441 2 digital_ldo_top_VIA4 $T=288530 17140 0 0 $X=288280 $Y=16910
X7442 2 digital_ldo_top_VIA4 $T=288530 21220 0 0 $X=288280 $Y=20990
X7443 2 digital_ldo_top_VIA4 $T=288530 25300 0 0 $X=288280 $Y=25070
X7444 2 digital_ldo_top_VIA4 $T=288530 86500 0 0 $X=288280 $Y=86270
X7445 2 digital_ldo_top_VIA4 $T=288530 90580 0 0 $X=288280 $Y=90350
X7446 2 digital_ldo_top_VIA4 $T=288530 94660 0 0 $X=288280 $Y=94430
X7447 2 digital_ldo_top_VIA4 $T=288530 98740 0 0 $X=288280 $Y=98510
X7448 2 digital_ldo_top_VIA4 $T=288530 102820 0 0 $X=288280 $Y=102590
X7449 2 digital_ldo_top_VIA4 $T=288530 106900 0 0 $X=288280 $Y=106670
X7450 2 digital_ldo_top_VIA4 $T=288530 110980 0 0 $X=288280 $Y=110750
X7451 2 digital_ldo_top_VIA4 $T=288530 115060 0 0 $X=288280 $Y=114830
X7452 2 digital_ldo_top_VIA4 $T=288530 119140 0 0 $X=288280 $Y=118910
X7453 2 digital_ldo_top_VIA4 $T=288530 123220 0 0 $X=288280 $Y=122990
X7454 2 digital_ldo_top_VIA4 $T=288530 127300 0 0 $X=288280 $Y=127070
X7455 3 digital_ldo_top_VIA4 $T=290830 11700 0 0 $X=290580 $Y=11470
X7456 3 digital_ldo_top_VIA4 $T=290830 15780 0 0 $X=290580 $Y=15550
X7457 3 digital_ldo_top_VIA4 $T=290830 93300 0 0 $X=290580 $Y=93070
X7458 3 digital_ldo_top_VIA4 $T=290830 97380 0 0 $X=290580 $Y=97150
X7459 3 digital_ldo_top_VIA4 $T=290830 101460 0 0 $X=290580 $Y=101230
X7460 3 digital_ldo_top_VIA4 $T=290830 105540 0 0 $X=290580 $Y=105310
X7461 3 digital_ldo_top_VIA4 $T=290830 109620 0 0 $X=290580 $Y=109390
X7462 3 digital_ldo_top_VIA4 $T=290830 113700 0 0 $X=290580 $Y=113470
X7463 3 digital_ldo_top_VIA4 $T=290830 117780 0 0 $X=290580 $Y=117550
X7464 3 digital_ldo_top_VIA4 $T=290830 121860 0 0 $X=290580 $Y=121630
X7465 3 digital_ldo_top_VIA4 $T=290830 125940 0 0 $X=290580 $Y=125710
X7466 2 digital_ldo_top_VIA4 $T=292210 13060 0 0 $X=291960 $Y=12830
X7467 2 digital_ldo_top_VIA4 $T=292210 17140 0 0 $X=291960 $Y=16910
X7468 2 digital_ldo_top_VIA4 $T=292210 94660 0 0 $X=291960 $Y=94430
X7469 2 digital_ldo_top_VIA4 $T=292210 98740 0 0 $X=291960 $Y=98510
X7470 2 digital_ldo_top_VIA4 $T=292210 102820 0 0 $X=291960 $Y=102590
X7471 2 digital_ldo_top_VIA4 $T=292210 106900 0 0 $X=291960 $Y=106670
X7472 2 digital_ldo_top_VIA4 $T=292210 110980 0 0 $X=291960 $Y=110750
X7473 2 digital_ldo_top_VIA4 $T=292210 115060 0 0 $X=291960 $Y=114830
X7474 2 digital_ldo_top_VIA4 $T=292210 119140 0 0 $X=291960 $Y=118910
X7475 2 digital_ldo_top_VIA4 $T=292210 123220 0 0 $X=291960 $Y=122990
X7476 2 digital_ldo_top_VIA4 $T=292210 127300 0 0 $X=291960 $Y=127070
X7477 3 digital_ldo_top_VIA4 $T=294510 11700 0 0 $X=294260 $Y=11470
X7478 3 digital_ldo_top_VIA4 $T=294510 15780 0 0 $X=294260 $Y=15550
X7479 3 digital_ldo_top_VIA4 $T=294510 32100 0 0 $X=294260 $Y=31870
X7480 3 digital_ldo_top_VIA4 $T=294510 85140 0 0 $X=294260 $Y=84910
X7481 3 digital_ldo_top_VIA4 $T=294510 89220 0 0 $X=294260 $Y=88990
X7482 3 digital_ldo_top_VIA4 $T=294510 93300 0 0 $X=294260 $Y=93070
X7483 3 digital_ldo_top_VIA4 $T=294510 97380 0 0 $X=294260 $Y=97150
X7484 3 digital_ldo_top_VIA4 $T=294510 101460 0 0 $X=294260 $Y=101230
X7485 3 digital_ldo_top_VIA4 $T=294510 105540 0 0 $X=294260 $Y=105310
X7486 3 digital_ldo_top_VIA4 $T=294510 109620 0 0 $X=294260 $Y=109390
X7487 3 digital_ldo_top_VIA4 $T=294510 113700 0 0 $X=294260 $Y=113470
X7488 3 digital_ldo_top_VIA4 $T=294510 117780 0 0 $X=294260 $Y=117550
X7489 3 digital_ldo_top_VIA4 $T=294510 121860 0 0 $X=294260 $Y=121630
X7490 3 digital_ldo_top_VIA4 $T=294510 125940 0 0 $X=294260 $Y=125710
X7491 2 digital_ldo_top_VIA4 $T=295890 13060 0 0 $X=295640 $Y=12830
X7492 2 digital_ldo_top_VIA4 $T=295890 17140 0 0 $X=295640 $Y=16910
X7493 2 digital_ldo_top_VIA4 $T=295890 21220 0 0 $X=295640 $Y=20990
X7494 2 digital_ldo_top_VIA4 $T=295890 25300 0 0 $X=295640 $Y=25070
X7495 2 digital_ldo_top_VIA4 $T=295890 86500 0 0 $X=295640 $Y=86270
X7496 2 digital_ldo_top_VIA4 $T=295890 90580 0 0 $X=295640 $Y=90350
X7497 2 digital_ldo_top_VIA4 $T=295890 94660 0 0 $X=295640 $Y=94430
X7498 2 digital_ldo_top_VIA4 $T=295890 98740 0 0 $X=295640 $Y=98510
X7499 2 digital_ldo_top_VIA4 $T=295890 102820 0 0 $X=295640 $Y=102590
X7500 2 digital_ldo_top_VIA4 $T=295890 106900 0 0 $X=295640 $Y=106670
X7501 2 digital_ldo_top_VIA4 $T=295890 110980 0 0 $X=295640 $Y=110750
X7502 2 digital_ldo_top_VIA4 $T=295890 115060 0 0 $X=295640 $Y=114830
X7503 2 digital_ldo_top_VIA4 $T=295890 119140 0 0 $X=295640 $Y=118910
X7504 2 digital_ldo_top_VIA4 $T=295890 123220 0 0 $X=295640 $Y=122990
X7505 2 digital_ldo_top_VIA4 $T=295890 127300 0 0 $X=295640 $Y=127070
X7506 3 digital_ldo_top_VIA4 $T=298190 11700 0 0 $X=297940 $Y=11470
X7507 3 digital_ldo_top_VIA4 $T=298190 15780 0 0 $X=297940 $Y=15550
X7508 3 digital_ldo_top_VIA4 $T=298190 19860 0 0 $X=297940 $Y=19630
X7509 3 digital_ldo_top_VIA4 $T=298190 23940 0 0 $X=297940 $Y=23710
X7510 3 digital_ldo_top_VIA4 $T=298190 32100 0 0 $X=297940 $Y=31870
X7511 3 digital_ldo_top_VIA4 $T=298190 85140 0 0 $X=297940 $Y=84910
X7512 3 digital_ldo_top_VIA4 $T=298190 89220 0 0 $X=297940 $Y=88990
X7513 3 digital_ldo_top_VIA4 $T=298190 93300 0 0 $X=297940 $Y=93070
X7514 3 digital_ldo_top_VIA4 $T=298190 97380 0 0 $X=297940 $Y=97150
X7515 3 digital_ldo_top_VIA4 $T=298190 101460 0 0 $X=297940 $Y=101230
X7516 3 digital_ldo_top_VIA4 $T=298190 105540 0 0 $X=297940 $Y=105310
X7517 3 digital_ldo_top_VIA4 $T=298190 109620 0 0 $X=297940 $Y=109390
X7518 3 digital_ldo_top_VIA4 $T=298190 113700 0 0 $X=297940 $Y=113470
X7519 3 digital_ldo_top_VIA4 $T=298190 117780 0 0 $X=297940 $Y=117550
X7520 3 digital_ldo_top_VIA4 $T=298190 121860 0 0 $X=297940 $Y=121630
X7521 3 digital_ldo_top_VIA4 $T=298190 125940 0 0 $X=297940 $Y=125710
X7522 2 digital_ldo_top_VIA4 $T=299570 13060 0 0 $X=299320 $Y=12830
X7523 2 digital_ldo_top_VIA4 $T=299570 17140 0 0 $X=299320 $Y=16910
X7524 2 digital_ldo_top_VIA4 $T=299570 21220 0 0 $X=299320 $Y=20990
X7525 2 digital_ldo_top_VIA4 $T=299570 25300 0 0 $X=299320 $Y=25070
X7526 2 digital_ldo_top_VIA4 $T=299570 86500 0 0 $X=299320 $Y=86270
X7527 2 digital_ldo_top_VIA4 $T=299570 90580 0 0 $X=299320 $Y=90350
X7528 2 digital_ldo_top_VIA4 $T=299570 94660 0 0 $X=299320 $Y=94430
X7529 2 digital_ldo_top_VIA4 $T=299570 98740 0 0 $X=299320 $Y=98510
X7530 2 digital_ldo_top_VIA4 $T=299570 102820 0 0 $X=299320 $Y=102590
X7531 2 digital_ldo_top_VIA4 $T=299570 106900 0 0 $X=299320 $Y=106670
X7532 2 digital_ldo_top_VIA4 $T=299570 110980 0 0 $X=299320 $Y=110750
X7533 2 digital_ldo_top_VIA4 $T=299570 115060 0 0 $X=299320 $Y=114830
X7534 2 digital_ldo_top_VIA4 $T=299570 119140 0 0 $X=299320 $Y=118910
X7535 2 digital_ldo_top_VIA4 $T=299570 123220 0 0 $X=299320 $Y=122990
X7536 2 digital_ldo_top_VIA4 $T=299570 127300 0 0 $X=299320 $Y=127070
X7537 3 digital_ldo_top_VIA4 $T=301870 11700 0 0 $X=301620 $Y=11470
X7538 3 digital_ldo_top_VIA4 $T=301870 15780 0 0 $X=301620 $Y=15550
X7539 3 digital_ldo_top_VIA4 $T=301870 19860 0 0 $X=301620 $Y=19630
X7540 3 digital_ldo_top_VIA4 $T=301870 23940 0 0 $X=301620 $Y=23710
X7541 3 digital_ldo_top_VIA4 $T=301870 32100 0 0 $X=301620 $Y=31870
X7542 3 digital_ldo_top_VIA4 $T=301870 85140 0 0 $X=301620 $Y=84910
X7543 3 digital_ldo_top_VIA4 $T=301870 89220 0 0 $X=301620 $Y=88990
X7544 3 digital_ldo_top_VIA4 $T=301870 93300 0 0 $X=301620 $Y=93070
X7545 3 digital_ldo_top_VIA4 $T=301870 97380 0 0 $X=301620 $Y=97150
X7546 3 digital_ldo_top_VIA4 $T=301870 101460 0 0 $X=301620 $Y=101230
X7547 3 digital_ldo_top_VIA4 $T=301870 105540 0 0 $X=301620 $Y=105310
X7548 3 digital_ldo_top_VIA4 $T=301870 109620 0 0 $X=301620 $Y=109390
X7549 3 digital_ldo_top_VIA4 $T=301870 113700 0 0 $X=301620 $Y=113470
X7550 3 digital_ldo_top_VIA4 $T=301870 117780 0 0 $X=301620 $Y=117550
X7551 3 digital_ldo_top_VIA4 $T=301870 121860 0 0 $X=301620 $Y=121630
X7552 3 digital_ldo_top_VIA4 $T=301870 125940 0 0 $X=301620 $Y=125710
X7553 2 digital_ldo_top_VIA4 $T=303250 13060 0 0 $X=303000 $Y=12830
X7554 2 digital_ldo_top_VIA4 $T=303250 17140 0 0 $X=303000 $Y=16910
X7555 2 digital_ldo_top_VIA4 $T=303250 21220 0 0 $X=303000 $Y=20990
X7556 2 digital_ldo_top_VIA4 $T=303250 25300 0 0 $X=303000 $Y=25070
X7557 2 digital_ldo_top_VIA4 $T=303250 86500 0 0 $X=303000 $Y=86270
X7558 2 digital_ldo_top_VIA4 $T=303250 90580 0 0 $X=303000 $Y=90350
X7559 2 digital_ldo_top_VIA4 $T=303250 94660 0 0 $X=303000 $Y=94430
X7560 2 digital_ldo_top_VIA4 $T=303250 98740 0 0 $X=303000 $Y=98510
X7561 2 digital_ldo_top_VIA4 $T=303250 102820 0 0 $X=303000 $Y=102590
X7562 2 digital_ldo_top_VIA4 $T=303250 106900 0 0 $X=303000 $Y=106670
X7563 2 digital_ldo_top_VIA4 $T=303250 110980 0 0 $X=303000 $Y=110750
X7564 2 digital_ldo_top_VIA4 $T=303250 115060 0 0 $X=303000 $Y=114830
X7565 2 digital_ldo_top_VIA4 $T=303250 119140 0 0 $X=303000 $Y=118910
X7566 2 digital_ldo_top_VIA4 $T=303250 123220 0 0 $X=303000 $Y=122990
X7567 2 digital_ldo_top_VIA4 $T=303250 127300 0 0 $X=303000 $Y=127070
X7568 3 digital_ldo_top_VIA4 $T=305550 11700 0 0 $X=305300 $Y=11470
X7569 3 digital_ldo_top_VIA4 $T=305550 15780 0 0 $X=305300 $Y=15550
X7570 3 digital_ldo_top_VIA4 $T=305550 19860 0 0 $X=305300 $Y=19630
X7571 3 digital_ldo_top_VIA4 $T=305550 23940 0 0 $X=305300 $Y=23710
X7572 3 digital_ldo_top_VIA4 $T=305550 32100 0 0 $X=305300 $Y=31870
X7573 3 digital_ldo_top_VIA4 $T=305550 85140 0 0 $X=305300 $Y=84910
X7574 3 digital_ldo_top_VIA4 $T=305550 89220 0 0 $X=305300 $Y=88990
X7575 3 digital_ldo_top_VIA4 $T=305550 93300 0 0 $X=305300 $Y=93070
X7576 3 digital_ldo_top_VIA4 $T=305550 97380 0 0 $X=305300 $Y=97150
X7577 3 digital_ldo_top_VIA4 $T=305550 101460 0 0 $X=305300 $Y=101230
X7578 3 digital_ldo_top_VIA4 $T=305550 105540 0 0 $X=305300 $Y=105310
X7579 3 digital_ldo_top_VIA4 $T=305550 109620 0 0 $X=305300 $Y=109390
X7580 3 digital_ldo_top_VIA4 $T=305550 113700 0 0 $X=305300 $Y=113470
X7581 3 digital_ldo_top_VIA4 $T=305550 117780 0 0 $X=305300 $Y=117550
X7582 3 digital_ldo_top_VIA4 $T=305550 121860 0 0 $X=305300 $Y=121630
X7583 3 digital_ldo_top_VIA4 $T=305550 125940 0 0 $X=305300 $Y=125710
X7584 2 digital_ldo_top_VIA4 $T=306930 13060 0 0 $X=306680 $Y=12830
X7585 2 digital_ldo_top_VIA4 $T=306930 17140 0 0 $X=306680 $Y=16910
X7586 2 digital_ldo_top_VIA4 $T=306930 21220 0 0 $X=306680 $Y=20990
X7587 2 digital_ldo_top_VIA4 $T=306930 25300 0 0 $X=306680 $Y=25070
X7588 2 digital_ldo_top_VIA4 $T=306930 86500 0 0 $X=306680 $Y=86270
X7589 2 digital_ldo_top_VIA4 $T=306930 90580 0 0 $X=306680 $Y=90350
X7590 2 digital_ldo_top_VIA4 $T=306930 94660 0 0 $X=306680 $Y=94430
X7591 2 digital_ldo_top_VIA4 $T=306930 98740 0 0 $X=306680 $Y=98510
X7592 2 digital_ldo_top_VIA4 $T=306930 102820 0 0 $X=306680 $Y=102590
X7593 2 digital_ldo_top_VIA4 $T=306930 106900 0 0 $X=306680 $Y=106670
X7594 2 digital_ldo_top_VIA4 $T=306930 110980 0 0 $X=306680 $Y=110750
X7595 2 digital_ldo_top_VIA4 $T=306930 115060 0 0 $X=306680 $Y=114830
X7596 2 digital_ldo_top_VIA4 $T=306930 119140 0 0 $X=306680 $Y=118910
X7597 2 digital_ldo_top_VIA4 $T=306930 123220 0 0 $X=306680 $Y=122990
X7598 2 digital_ldo_top_VIA4 $T=306930 127300 0 0 $X=306680 $Y=127070
X7599 3 digital_ldo_top_VIA4 $T=309230 11700 0 0 $X=308980 $Y=11470
X7600 3 digital_ldo_top_VIA4 $T=309230 15780 0 0 $X=308980 $Y=15550
X7601 3 digital_ldo_top_VIA4 $T=309230 19860 0 0 $X=308980 $Y=19630
X7602 3 digital_ldo_top_VIA4 $T=309230 23940 0 0 $X=308980 $Y=23710
X7603 3 digital_ldo_top_VIA4 $T=309230 28020 0 0 $X=308980 $Y=27790
X7604 3 digital_ldo_top_VIA4 $T=309230 32100 0 0 $X=308980 $Y=31870
X7605 3 digital_ldo_top_VIA4 $T=309230 36180 0 0 $X=308980 $Y=35950
X7606 3 digital_ldo_top_VIA4 $T=309230 40260 0 0 $X=308980 $Y=40030
X7607 3 digital_ldo_top_VIA4 $T=309230 44340 0 0 $X=308980 $Y=44110
X7608 3 digital_ldo_top_VIA4 $T=309230 48420 0 0 $X=308980 $Y=48190
X7609 3 digital_ldo_top_VIA4 $T=309230 52500 0 0 $X=308980 $Y=52270
X7610 3 digital_ldo_top_VIA4 $T=309230 56580 0 0 $X=308980 $Y=56350
X7611 3 digital_ldo_top_VIA4 $T=309230 60660 0 0 $X=308980 $Y=60430
X7612 3 digital_ldo_top_VIA4 $T=309230 64740 0 0 $X=308980 $Y=64510
X7613 3 digital_ldo_top_VIA4 $T=309230 68820 0 0 $X=308980 $Y=68590
X7614 3 digital_ldo_top_VIA4 $T=309230 72900 0 0 $X=308980 $Y=72670
X7615 3 digital_ldo_top_VIA4 $T=309230 76980 0 0 $X=308980 $Y=76750
X7616 3 digital_ldo_top_VIA4 $T=309230 81060 0 0 $X=308980 $Y=80830
X7617 3 digital_ldo_top_VIA4 $T=309230 85140 0 0 $X=308980 $Y=84910
X7618 3 digital_ldo_top_VIA4 $T=309230 89220 0 0 $X=308980 $Y=88990
X7619 3 digital_ldo_top_VIA4 $T=309230 93300 0 0 $X=308980 $Y=93070
X7620 3 digital_ldo_top_VIA4 $T=309230 97380 0 0 $X=308980 $Y=97150
X7621 3 digital_ldo_top_VIA4 $T=309230 101460 0 0 $X=308980 $Y=101230
X7622 3 digital_ldo_top_VIA4 $T=309230 105540 0 0 $X=308980 $Y=105310
X7623 3 digital_ldo_top_VIA4 $T=309230 109620 0 0 $X=308980 $Y=109390
X7624 3 digital_ldo_top_VIA4 $T=309230 113700 0 0 $X=308980 $Y=113470
X7625 3 digital_ldo_top_VIA4 $T=309230 117780 0 0 $X=308980 $Y=117550
X7626 3 digital_ldo_top_VIA4 $T=309230 121860 0 0 $X=308980 $Y=121630
X7627 3 digital_ldo_top_VIA4 $T=309230 125940 0 0 $X=308980 $Y=125710
X7628 2 digital_ldo_top_VIA4 $T=310610 13060 0 0 $X=310360 $Y=12830
X7629 2 digital_ldo_top_VIA4 $T=310610 17140 0 0 $X=310360 $Y=16910
X7630 2 digital_ldo_top_VIA4 $T=310610 21220 0 0 $X=310360 $Y=20990
X7631 2 digital_ldo_top_VIA4 $T=310610 25300 0 0 $X=310360 $Y=25070
X7632 2 digital_ldo_top_VIA4 $T=310610 29380 0 0 $X=310360 $Y=29150
X7633 2 digital_ldo_top_VIA4 $T=310610 33460 0 0 $X=310360 $Y=33230
X7634 2 digital_ldo_top_VIA4 $T=310610 37540 0 0 $X=310360 $Y=37310
X7635 2 digital_ldo_top_VIA4 $T=310610 41620 0 0 $X=310360 $Y=41390
X7636 2 digital_ldo_top_VIA4 $T=310610 45700 0 0 $X=310360 $Y=45470
X7637 2 digital_ldo_top_VIA4 $T=310610 49780 0 0 $X=310360 $Y=49550
X7638 2 digital_ldo_top_VIA4 $T=310610 53860 0 0 $X=310360 $Y=53630
X7639 2 digital_ldo_top_VIA4 $T=310610 57940 0 0 $X=310360 $Y=57710
X7640 2 digital_ldo_top_VIA4 $T=310610 62020 0 0 $X=310360 $Y=61790
X7641 2 digital_ldo_top_VIA4 $T=310610 66100 0 0 $X=310360 $Y=65870
X7642 2 digital_ldo_top_VIA4 $T=310610 70180 0 0 $X=310360 $Y=69950
X7643 2 digital_ldo_top_VIA4 $T=310610 74260 0 0 $X=310360 $Y=74030
X7644 2 digital_ldo_top_VIA4 $T=310610 78340 0 0 $X=310360 $Y=78110
X7645 2 digital_ldo_top_VIA4 $T=310610 82420 0 0 $X=310360 $Y=82190
X7646 2 digital_ldo_top_VIA4 $T=310610 86500 0 0 $X=310360 $Y=86270
X7647 2 digital_ldo_top_VIA4 $T=310610 90580 0 0 $X=310360 $Y=90350
X7648 2 digital_ldo_top_VIA4 $T=310610 94660 0 0 $X=310360 $Y=94430
X7649 2 digital_ldo_top_VIA4 $T=310610 98740 0 0 $X=310360 $Y=98510
X7650 2 digital_ldo_top_VIA4 $T=310610 102820 0 0 $X=310360 $Y=102590
X7651 2 digital_ldo_top_VIA4 $T=310610 106900 0 0 $X=310360 $Y=106670
X7652 2 digital_ldo_top_VIA4 $T=310610 110980 0 0 $X=310360 $Y=110750
X7653 2 digital_ldo_top_VIA4 $T=310610 115060 0 0 $X=310360 $Y=114830
X7654 2 digital_ldo_top_VIA4 $T=310610 119140 0 0 $X=310360 $Y=118910
X7655 2 digital_ldo_top_VIA4 $T=310610 123220 0 0 $X=310360 $Y=122990
X7656 2 digital_ldo_top_VIA4 $T=310610 127300 0 0 $X=310360 $Y=127070
X7657 3 digital_ldo_top_VIA4 $T=312910 11700 0 0 $X=312660 $Y=11470
X7658 3 digital_ldo_top_VIA4 $T=312910 15780 0 0 $X=312660 $Y=15550
X7659 3 digital_ldo_top_VIA4 $T=312910 19860 0 0 $X=312660 $Y=19630
X7660 3 digital_ldo_top_VIA4 $T=312910 23940 0 0 $X=312660 $Y=23710
X7661 3 digital_ldo_top_VIA4 $T=312910 28020 0 0 $X=312660 $Y=27790
X7662 3 digital_ldo_top_VIA4 $T=312910 32100 0 0 $X=312660 $Y=31870
X7663 3 digital_ldo_top_VIA4 $T=312910 36180 0 0 $X=312660 $Y=35950
X7664 3 digital_ldo_top_VIA4 $T=312910 40260 0 0 $X=312660 $Y=40030
X7665 3 digital_ldo_top_VIA4 $T=312910 44340 0 0 $X=312660 $Y=44110
X7666 3 digital_ldo_top_VIA4 $T=312910 48420 0 0 $X=312660 $Y=48190
X7667 3 digital_ldo_top_VIA4 $T=312910 52500 0 0 $X=312660 $Y=52270
X7668 3 digital_ldo_top_VIA4 $T=312910 56580 0 0 $X=312660 $Y=56350
X7669 3 digital_ldo_top_VIA4 $T=312910 60660 0 0 $X=312660 $Y=60430
X7670 3 digital_ldo_top_VIA4 $T=312910 64740 0 0 $X=312660 $Y=64510
X7671 3 digital_ldo_top_VIA4 $T=312910 68820 0 0 $X=312660 $Y=68590
X7672 3 digital_ldo_top_VIA4 $T=312910 72900 0 0 $X=312660 $Y=72670
X7673 3 digital_ldo_top_VIA4 $T=312910 76980 0 0 $X=312660 $Y=76750
X7674 3 digital_ldo_top_VIA4 $T=312910 81060 0 0 $X=312660 $Y=80830
X7675 3 digital_ldo_top_VIA4 $T=312910 85140 0 0 $X=312660 $Y=84910
X7676 3 digital_ldo_top_VIA4 $T=312910 89220 0 0 $X=312660 $Y=88990
X7677 3 digital_ldo_top_VIA4 $T=312910 93300 0 0 $X=312660 $Y=93070
X7678 3 digital_ldo_top_VIA4 $T=312910 97380 0 0 $X=312660 $Y=97150
X7679 3 digital_ldo_top_VIA4 $T=312910 101460 0 0 $X=312660 $Y=101230
X7680 3 digital_ldo_top_VIA4 $T=312910 105540 0 0 $X=312660 $Y=105310
X7681 3 digital_ldo_top_VIA4 $T=312910 109620 0 0 $X=312660 $Y=109390
X7682 3 digital_ldo_top_VIA4 $T=312910 113700 0 0 $X=312660 $Y=113470
X7683 3 digital_ldo_top_VIA4 $T=312910 117780 0 0 $X=312660 $Y=117550
X7684 3 digital_ldo_top_VIA4 $T=312910 121860 0 0 $X=312660 $Y=121630
X7685 3 digital_ldo_top_VIA4 $T=312910 125940 0 0 $X=312660 $Y=125710
X7686 2 digital_ldo_top_VIA4 $T=314290 13060 0 0 $X=314040 $Y=12830
X7687 2 digital_ldo_top_VIA4 $T=314290 17140 0 0 $X=314040 $Y=16910
X7688 2 digital_ldo_top_VIA4 $T=314290 21220 0 0 $X=314040 $Y=20990
X7689 2 digital_ldo_top_VIA4 $T=314290 25300 0 0 $X=314040 $Y=25070
X7690 2 digital_ldo_top_VIA4 $T=314290 29380 0 0 $X=314040 $Y=29150
X7691 2 digital_ldo_top_VIA4 $T=314290 33460 0 0 $X=314040 $Y=33230
X7692 2 digital_ldo_top_VIA4 $T=314290 37540 0 0 $X=314040 $Y=37310
X7693 2 digital_ldo_top_VIA4 $T=314290 41620 0 0 $X=314040 $Y=41390
X7694 2 digital_ldo_top_VIA4 $T=314290 45700 0 0 $X=314040 $Y=45470
X7695 2 digital_ldo_top_VIA4 $T=314290 49780 0 0 $X=314040 $Y=49550
X7696 2 digital_ldo_top_VIA4 $T=314290 53860 0 0 $X=314040 $Y=53630
X7697 2 digital_ldo_top_VIA4 $T=314290 57940 0 0 $X=314040 $Y=57710
X7698 2 digital_ldo_top_VIA4 $T=314290 62020 0 0 $X=314040 $Y=61790
X7699 2 digital_ldo_top_VIA4 $T=314290 66100 0 0 $X=314040 $Y=65870
X7700 2 digital_ldo_top_VIA4 $T=314290 70180 0 0 $X=314040 $Y=69950
X7701 2 digital_ldo_top_VIA4 $T=314290 74260 0 0 $X=314040 $Y=74030
X7702 2 digital_ldo_top_VIA4 $T=314290 78340 0 0 $X=314040 $Y=78110
X7703 2 digital_ldo_top_VIA4 $T=314290 82420 0 0 $X=314040 $Y=82190
X7704 2 digital_ldo_top_VIA4 $T=314290 86500 0 0 $X=314040 $Y=86270
X7705 2 digital_ldo_top_VIA4 $T=314290 90580 0 0 $X=314040 $Y=90350
X7706 2 digital_ldo_top_VIA4 $T=314290 94660 0 0 $X=314040 $Y=94430
X7707 2 digital_ldo_top_VIA4 $T=314290 98740 0 0 $X=314040 $Y=98510
X7708 2 digital_ldo_top_VIA4 $T=314290 102820 0 0 $X=314040 $Y=102590
X7709 2 digital_ldo_top_VIA4 $T=314290 106900 0 0 $X=314040 $Y=106670
X7710 2 digital_ldo_top_VIA4 $T=314290 110980 0 0 $X=314040 $Y=110750
X7711 2 digital_ldo_top_VIA4 $T=314290 115060 0 0 $X=314040 $Y=114830
X7712 2 digital_ldo_top_VIA4 $T=314290 119140 0 0 $X=314040 $Y=118910
X7713 2 digital_ldo_top_VIA4 $T=314290 123220 0 0 $X=314040 $Y=122990
X7714 2 digital_ldo_top_VIA4 $T=314290 127300 0 0 $X=314040 $Y=127070
X7715 3 digital_ldo_top_VIA4 $T=316590 11700 0 0 $X=316340 $Y=11470
X7716 3 digital_ldo_top_VIA4 $T=316590 15780 0 0 $X=316340 $Y=15550
X7717 3 digital_ldo_top_VIA4 $T=316590 19860 0 0 $X=316340 $Y=19630
X7718 3 digital_ldo_top_VIA4 $T=316590 23940 0 0 $X=316340 $Y=23710
X7719 3 digital_ldo_top_VIA4 $T=316590 28020 0 0 $X=316340 $Y=27790
X7720 3 digital_ldo_top_VIA4 $T=316590 32100 0 0 $X=316340 $Y=31870
X7721 3 digital_ldo_top_VIA4 $T=316590 36180 0 0 $X=316340 $Y=35950
X7722 3 digital_ldo_top_VIA4 $T=316590 40260 0 0 $X=316340 $Y=40030
X7723 3 digital_ldo_top_VIA4 $T=316590 44340 0 0 $X=316340 $Y=44110
X7724 3 digital_ldo_top_VIA4 $T=316590 48420 0 0 $X=316340 $Y=48190
X7725 3 digital_ldo_top_VIA4 $T=316590 52500 0 0 $X=316340 $Y=52270
X7726 3 digital_ldo_top_VIA4 $T=316590 56580 0 0 $X=316340 $Y=56350
X7727 3 digital_ldo_top_VIA4 $T=316590 60660 0 0 $X=316340 $Y=60430
X7728 3 digital_ldo_top_VIA4 $T=316590 64740 0 0 $X=316340 $Y=64510
X7729 3 digital_ldo_top_VIA4 $T=316590 68820 0 0 $X=316340 $Y=68590
X7730 3 digital_ldo_top_VIA4 $T=316590 72900 0 0 $X=316340 $Y=72670
X7731 3 digital_ldo_top_VIA4 $T=316590 76980 0 0 $X=316340 $Y=76750
X7732 3 digital_ldo_top_VIA4 $T=316590 81060 0 0 $X=316340 $Y=80830
X7733 3 digital_ldo_top_VIA4 $T=316590 85140 0 0 $X=316340 $Y=84910
X7734 3 digital_ldo_top_VIA4 $T=316590 89220 0 0 $X=316340 $Y=88990
X7735 3 digital_ldo_top_VIA4 $T=316590 93300 0 0 $X=316340 $Y=93070
X7736 3 digital_ldo_top_VIA4 $T=316590 97380 0 0 $X=316340 $Y=97150
X7737 3 digital_ldo_top_VIA4 $T=316590 101460 0 0 $X=316340 $Y=101230
X7738 3 digital_ldo_top_VIA4 $T=316590 105540 0 0 $X=316340 $Y=105310
X7739 3 digital_ldo_top_VIA4 $T=316590 109620 0 0 $X=316340 $Y=109390
X7740 3 digital_ldo_top_VIA4 $T=316590 113700 0 0 $X=316340 $Y=113470
X7741 3 digital_ldo_top_VIA4 $T=316590 117780 0 0 $X=316340 $Y=117550
X7742 3 digital_ldo_top_VIA4 $T=316590 121860 0 0 $X=316340 $Y=121630
X7743 3 digital_ldo_top_VIA4 $T=316590 125940 0 0 $X=316340 $Y=125710
X7744 2 digital_ldo_top_VIA4 $T=317970 13060 0 0 $X=317720 $Y=12830
X7745 2 digital_ldo_top_VIA4 $T=317970 17140 0 0 $X=317720 $Y=16910
X7746 2 digital_ldo_top_VIA4 $T=317970 21220 0 0 $X=317720 $Y=20990
X7747 2 digital_ldo_top_VIA4 $T=317970 25300 0 0 $X=317720 $Y=25070
X7748 2 digital_ldo_top_VIA4 $T=317970 29380 0 0 $X=317720 $Y=29150
X7749 2 digital_ldo_top_VIA4 $T=317970 33460 0 0 $X=317720 $Y=33230
X7750 2 digital_ldo_top_VIA4 $T=317970 37540 0 0 $X=317720 $Y=37310
X7751 2 digital_ldo_top_VIA4 $T=317970 41620 0 0 $X=317720 $Y=41390
X7752 2 digital_ldo_top_VIA4 $T=317970 45700 0 0 $X=317720 $Y=45470
X7753 2 digital_ldo_top_VIA4 $T=317970 49780 0 0 $X=317720 $Y=49550
X7754 2 digital_ldo_top_VIA4 $T=317970 53860 0 0 $X=317720 $Y=53630
X7755 2 digital_ldo_top_VIA4 $T=317970 57940 0 0 $X=317720 $Y=57710
X7756 2 digital_ldo_top_VIA4 $T=317970 62020 0 0 $X=317720 $Y=61790
X7757 2 digital_ldo_top_VIA4 $T=317970 66100 0 0 $X=317720 $Y=65870
X7758 2 digital_ldo_top_VIA4 $T=317970 70180 0 0 $X=317720 $Y=69950
X7759 2 digital_ldo_top_VIA4 $T=317970 74260 0 0 $X=317720 $Y=74030
X7760 2 digital_ldo_top_VIA4 $T=317970 78340 0 0 $X=317720 $Y=78110
X7761 2 digital_ldo_top_VIA4 $T=317970 82420 0 0 $X=317720 $Y=82190
X7762 2 digital_ldo_top_VIA4 $T=317970 86500 0 0 $X=317720 $Y=86270
X7763 2 digital_ldo_top_VIA4 $T=317970 90580 0 0 $X=317720 $Y=90350
X7764 2 digital_ldo_top_VIA4 $T=317970 94660 0 0 $X=317720 $Y=94430
X7765 2 digital_ldo_top_VIA4 $T=317970 98740 0 0 $X=317720 $Y=98510
X7766 2 digital_ldo_top_VIA4 $T=317970 102820 0 0 $X=317720 $Y=102590
X7767 2 digital_ldo_top_VIA4 $T=317970 106900 0 0 $X=317720 $Y=106670
X7768 2 digital_ldo_top_VIA4 $T=317970 110980 0 0 $X=317720 $Y=110750
X7769 2 digital_ldo_top_VIA4 $T=317970 115060 0 0 $X=317720 $Y=114830
X7770 2 digital_ldo_top_VIA4 $T=317970 119140 0 0 $X=317720 $Y=118910
X7771 2 digital_ldo_top_VIA4 $T=317970 123220 0 0 $X=317720 $Y=122990
X7772 2 digital_ldo_top_VIA4 $T=317970 127300 0 0 $X=317720 $Y=127070
X7773 3 digital_ldo_top_VIA4 $T=320270 11700 0 0 $X=320020 $Y=11470
X7774 3 digital_ldo_top_VIA4 $T=320270 15780 0 0 $X=320020 $Y=15550
X7775 3 digital_ldo_top_VIA4 $T=320270 19860 0 0 $X=320020 $Y=19630
X7776 3 digital_ldo_top_VIA4 $T=320270 23940 0 0 $X=320020 $Y=23710
X7777 3 digital_ldo_top_VIA4 $T=320270 28020 0 0 $X=320020 $Y=27790
X7778 3 digital_ldo_top_VIA4 $T=320270 32100 0 0 $X=320020 $Y=31870
X7779 3 digital_ldo_top_VIA4 $T=320270 36180 0 0 $X=320020 $Y=35950
X7780 3 digital_ldo_top_VIA4 $T=320270 40260 0 0 $X=320020 $Y=40030
X7781 3 digital_ldo_top_VIA4 $T=320270 44340 0 0 $X=320020 $Y=44110
X7782 3 digital_ldo_top_VIA4 $T=320270 48420 0 0 $X=320020 $Y=48190
X7783 3 digital_ldo_top_VIA4 $T=320270 52500 0 0 $X=320020 $Y=52270
X7784 3 digital_ldo_top_VIA4 $T=320270 56580 0 0 $X=320020 $Y=56350
X7785 3 digital_ldo_top_VIA4 $T=320270 60660 0 0 $X=320020 $Y=60430
X7786 3 digital_ldo_top_VIA4 $T=320270 64740 0 0 $X=320020 $Y=64510
X7787 3 digital_ldo_top_VIA4 $T=320270 68820 0 0 $X=320020 $Y=68590
X7788 3 digital_ldo_top_VIA4 $T=320270 72900 0 0 $X=320020 $Y=72670
X7789 3 digital_ldo_top_VIA4 $T=320270 76980 0 0 $X=320020 $Y=76750
X7790 3 digital_ldo_top_VIA4 $T=320270 81060 0 0 $X=320020 $Y=80830
X7791 3 digital_ldo_top_VIA4 $T=320270 85140 0 0 $X=320020 $Y=84910
X7792 3 digital_ldo_top_VIA4 $T=320270 89220 0 0 $X=320020 $Y=88990
X7793 3 digital_ldo_top_VIA4 $T=320270 93300 0 0 $X=320020 $Y=93070
X7794 3 digital_ldo_top_VIA4 $T=320270 97380 0 0 $X=320020 $Y=97150
X7795 3 digital_ldo_top_VIA4 $T=320270 101460 0 0 $X=320020 $Y=101230
X7796 3 digital_ldo_top_VIA4 $T=320270 105540 0 0 $X=320020 $Y=105310
X7797 3 digital_ldo_top_VIA4 $T=320270 109620 0 0 $X=320020 $Y=109390
X7798 3 digital_ldo_top_VIA4 $T=320270 113700 0 0 $X=320020 $Y=113470
X7799 3 digital_ldo_top_VIA4 $T=320270 117780 0 0 $X=320020 $Y=117550
X7800 3 digital_ldo_top_VIA4 $T=320270 121860 0 0 $X=320020 $Y=121630
X7801 3 digital_ldo_top_VIA4 $T=320270 125940 0 0 $X=320020 $Y=125710
X7802 2 digital_ldo_top_VIA4 $T=321650 13060 0 0 $X=321400 $Y=12830
X7803 2 digital_ldo_top_VIA4 $T=321650 17140 0 0 $X=321400 $Y=16910
X7804 2 digital_ldo_top_VIA4 $T=321650 21220 0 0 $X=321400 $Y=20990
X7805 2 digital_ldo_top_VIA4 $T=321650 25300 0 0 $X=321400 $Y=25070
X7806 2 digital_ldo_top_VIA4 $T=321650 29380 0 0 $X=321400 $Y=29150
X7807 2 digital_ldo_top_VIA4 $T=321650 33460 0 0 $X=321400 $Y=33230
X7808 2 digital_ldo_top_VIA4 $T=321650 37540 0 0 $X=321400 $Y=37310
X7809 2 digital_ldo_top_VIA4 $T=321650 41620 0 0 $X=321400 $Y=41390
X7810 2 digital_ldo_top_VIA4 $T=321650 45700 0 0 $X=321400 $Y=45470
X7811 2 digital_ldo_top_VIA4 $T=321650 49780 0 0 $X=321400 $Y=49550
X7812 2 digital_ldo_top_VIA4 $T=321650 53860 0 0 $X=321400 $Y=53630
X7813 2 digital_ldo_top_VIA4 $T=321650 57940 0 0 $X=321400 $Y=57710
X7814 2 digital_ldo_top_VIA4 $T=321650 62020 0 0 $X=321400 $Y=61790
X7815 2 digital_ldo_top_VIA4 $T=321650 66100 0 0 $X=321400 $Y=65870
X7816 2 digital_ldo_top_VIA4 $T=321650 70180 0 0 $X=321400 $Y=69950
X7817 2 digital_ldo_top_VIA4 $T=321650 74260 0 0 $X=321400 $Y=74030
X7818 2 digital_ldo_top_VIA4 $T=321650 78340 0 0 $X=321400 $Y=78110
X7819 2 digital_ldo_top_VIA4 $T=321650 82420 0 0 $X=321400 $Y=82190
X7820 2 digital_ldo_top_VIA4 $T=321650 86500 0 0 $X=321400 $Y=86270
X7821 2 digital_ldo_top_VIA4 $T=321650 90580 0 0 $X=321400 $Y=90350
X7822 2 digital_ldo_top_VIA4 $T=321650 94660 0 0 $X=321400 $Y=94430
X7823 2 digital_ldo_top_VIA4 $T=321650 98740 0 0 $X=321400 $Y=98510
X7824 2 digital_ldo_top_VIA4 $T=321650 102820 0 0 $X=321400 $Y=102590
X7825 2 digital_ldo_top_VIA4 $T=321650 106900 0 0 $X=321400 $Y=106670
X7826 2 digital_ldo_top_VIA4 $T=321650 110980 0 0 $X=321400 $Y=110750
X7827 2 digital_ldo_top_VIA4 $T=321650 115060 0 0 $X=321400 $Y=114830
X7828 2 digital_ldo_top_VIA4 $T=321650 119140 0 0 $X=321400 $Y=118910
X7829 2 digital_ldo_top_VIA4 $T=321650 123220 0 0 $X=321400 $Y=122990
X7830 2 digital_ldo_top_VIA4 $T=321650 127300 0 0 $X=321400 $Y=127070
X7831 3 digital_ldo_top_VIA4 $T=323950 11700 0 0 $X=323700 $Y=11470
X7832 3 digital_ldo_top_VIA4 $T=323950 52500 0 0 $X=323700 $Y=52270
X7833 3 digital_ldo_top_VIA4 $T=323950 56580 0 0 $X=323700 $Y=56350
X7834 3 digital_ldo_top_VIA4 $T=323950 60660 0 0 $X=323700 $Y=60430
X7835 3 digital_ldo_top_VIA4 $T=323950 64740 0 0 $X=323700 $Y=64510
X7836 3 digital_ldo_top_VIA4 $T=323950 68820 0 0 $X=323700 $Y=68590
X7837 3 digital_ldo_top_VIA4 $T=323950 72900 0 0 $X=323700 $Y=72670
X7838 3 digital_ldo_top_VIA4 $T=323950 76980 0 0 $X=323700 $Y=76750
X7839 3 digital_ldo_top_VIA4 $T=323950 81060 0 0 $X=323700 $Y=80830
X7840 3 digital_ldo_top_VIA4 $T=323950 85140 0 0 $X=323700 $Y=84910
X7841 3 digital_ldo_top_VIA4 $T=323950 89220 0 0 $X=323700 $Y=88990
X7842 3 digital_ldo_top_VIA4 $T=323950 93300 0 0 $X=323700 $Y=93070
X7843 3 digital_ldo_top_VIA4 $T=323950 97380 0 0 $X=323700 $Y=97150
X7844 3 digital_ldo_top_VIA4 $T=323950 101460 0 0 $X=323700 $Y=101230
X7845 3 digital_ldo_top_VIA4 $T=323950 105540 0 0 $X=323700 $Y=105310
X7846 3 digital_ldo_top_VIA4 $T=323950 109620 0 0 $X=323700 $Y=109390
X7847 3 digital_ldo_top_VIA4 $T=323950 113700 0 0 $X=323700 $Y=113470
X7848 3 digital_ldo_top_VIA4 $T=323950 117780 0 0 $X=323700 $Y=117550
X7849 3 digital_ldo_top_VIA4 $T=323950 121860 0 0 $X=323700 $Y=121630
X7850 3 digital_ldo_top_VIA4 $T=323950 125940 0 0 $X=323700 $Y=125710
X7851 2 digital_ldo_top_VIA4 $T=325330 13060 0 0 $X=325080 $Y=12830
X7852 2 digital_ldo_top_VIA4 $T=325330 49780 0 0 $X=325080 $Y=49550
X7853 2 digital_ldo_top_VIA4 $T=325330 53860 0 0 $X=325080 $Y=53630
X7854 2 digital_ldo_top_VIA4 $T=325330 57940 0 0 $X=325080 $Y=57710
X7855 2 digital_ldo_top_VIA4 $T=325330 62020 0 0 $X=325080 $Y=61790
X7856 2 digital_ldo_top_VIA4 $T=325330 66100 0 0 $X=325080 $Y=65870
X7857 2 digital_ldo_top_VIA4 $T=325330 70180 0 0 $X=325080 $Y=69950
X7858 2 digital_ldo_top_VIA4 $T=325330 74260 0 0 $X=325080 $Y=74030
X7859 2 digital_ldo_top_VIA4 $T=325330 78340 0 0 $X=325080 $Y=78110
X7860 2 digital_ldo_top_VIA4 $T=325330 82420 0 0 $X=325080 $Y=82190
X7861 2 digital_ldo_top_VIA4 $T=325330 86500 0 0 $X=325080 $Y=86270
X7862 2 digital_ldo_top_VIA4 $T=325330 90580 0 0 $X=325080 $Y=90350
X7863 2 digital_ldo_top_VIA4 $T=325330 94660 0 0 $X=325080 $Y=94430
X7864 2 digital_ldo_top_VIA4 $T=325330 98740 0 0 $X=325080 $Y=98510
X7865 2 digital_ldo_top_VIA4 $T=325330 102820 0 0 $X=325080 $Y=102590
X7866 2 digital_ldo_top_VIA4 $T=325330 106900 0 0 $X=325080 $Y=106670
X7867 2 digital_ldo_top_VIA4 $T=325330 110980 0 0 $X=325080 $Y=110750
X7868 2 digital_ldo_top_VIA4 $T=325330 115060 0 0 $X=325080 $Y=114830
X7869 2 digital_ldo_top_VIA4 $T=325330 119140 0 0 $X=325080 $Y=118910
X7870 2 digital_ldo_top_VIA4 $T=325330 123220 0 0 $X=325080 $Y=122990
X7871 2 digital_ldo_top_VIA4 $T=325330 127300 0 0 $X=325080 $Y=127070
X7872 3 digital_ldo_top_VIA4 $T=327630 11700 0 0 $X=327380 $Y=11470
X7873 3 digital_ldo_top_VIA4 $T=327630 52500 0 0 $X=327380 $Y=52270
X7874 3 digital_ldo_top_VIA4 $T=327630 56580 0 0 $X=327380 $Y=56350
X7875 3 digital_ldo_top_VIA4 $T=327630 60660 0 0 $X=327380 $Y=60430
X7876 3 digital_ldo_top_VIA4 $T=327630 64740 0 0 $X=327380 $Y=64510
X7877 3 digital_ldo_top_VIA4 $T=327630 68820 0 0 $X=327380 $Y=68590
X7878 3 digital_ldo_top_VIA4 $T=327630 72900 0 0 $X=327380 $Y=72670
X7879 3 digital_ldo_top_VIA4 $T=327630 76980 0 0 $X=327380 $Y=76750
X7880 3 digital_ldo_top_VIA4 $T=327630 81060 0 0 $X=327380 $Y=80830
X7881 3 digital_ldo_top_VIA4 $T=327630 85140 0 0 $X=327380 $Y=84910
X7882 3 digital_ldo_top_VIA4 $T=327630 89220 0 0 $X=327380 $Y=88990
X7883 3 digital_ldo_top_VIA4 $T=327630 93300 0 0 $X=327380 $Y=93070
X7884 3 digital_ldo_top_VIA4 $T=327630 97380 0 0 $X=327380 $Y=97150
X7885 3 digital_ldo_top_VIA4 $T=327630 101460 0 0 $X=327380 $Y=101230
X7886 3 digital_ldo_top_VIA4 $T=327630 105540 0 0 $X=327380 $Y=105310
X7887 3 digital_ldo_top_VIA4 $T=327630 109620 0 0 $X=327380 $Y=109390
X7888 3 digital_ldo_top_VIA4 $T=327630 113700 0 0 $X=327380 $Y=113470
X7889 3 digital_ldo_top_VIA4 $T=327630 117780 0 0 $X=327380 $Y=117550
X7890 3 digital_ldo_top_VIA4 $T=327630 121860 0 0 $X=327380 $Y=121630
X7891 3 digital_ldo_top_VIA4 $T=327630 125940 0 0 $X=327380 $Y=125710
X7892 2 digital_ldo_top_VIA4 $T=329010 13060 0 0 $X=328760 $Y=12830
X7893 2 digital_ldo_top_VIA4 $T=329010 49780 0 0 $X=328760 $Y=49550
X7894 2 digital_ldo_top_VIA4 $T=329010 53860 0 0 $X=328760 $Y=53630
X7895 2 digital_ldo_top_VIA4 $T=329010 57940 0 0 $X=328760 $Y=57710
X7896 2 digital_ldo_top_VIA4 $T=329010 62020 0 0 $X=328760 $Y=61790
X7897 2 digital_ldo_top_VIA4 $T=329010 66100 0 0 $X=328760 $Y=65870
X7898 2 digital_ldo_top_VIA4 $T=329010 70180 0 0 $X=328760 $Y=69950
X7899 2 digital_ldo_top_VIA4 $T=329010 74260 0 0 $X=328760 $Y=74030
X7900 2 digital_ldo_top_VIA4 $T=329010 78340 0 0 $X=328760 $Y=78110
X7901 2 digital_ldo_top_VIA4 $T=329010 82420 0 0 $X=328760 $Y=82190
X7902 2 digital_ldo_top_VIA4 $T=329010 86500 0 0 $X=328760 $Y=86270
X7903 2 digital_ldo_top_VIA4 $T=329010 90580 0 0 $X=328760 $Y=90350
X7904 2 digital_ldo_top_VIA4 $T=329010 94660 0 0 $X=328760 $Y=94430
X7905 2 digital_ldo_top_VIA4 $T=329010 98740 0 0 $X=328760 $Y=98510
X7906 2 digital_ldo_top_VIA4 $T=329010 102820 0 0 $X=328760 $Y=102590
X7907 2 digital_ldo_top_VIA4 $T=329010 106900 0 0 $X=328760 $Y=106670
X7908 2 digital_ldo_top_VIA4 $T=329010 110980 0 0 $X=328760 $Y=110750
X7909 2 digital_ldo_top_VIA4 $T=329010 115060 0 0 $X=328760 $Y=114830
X7910 2 digital_ldo_top_VIA4 $T=329010 119140 0 0 $X=328760 $Y=118910
X7911 2 digital_ldo_top_VIA4 $T=329010 123220 0 0 $X=328760 $Y=122990
X7912 2 digital_ldo_top_VIA4 $T=329010 127300 0 0 $X=328760 $Y=127070
X7913 3 digital_ldo_top_VIA4 $T=331310 11700 0 0 $X=331060 $Y=11470
X7914 3 digital_ldo_top_VIA4 $T=331310 52500 0 0 $X=331060 $Y=52270
X7915 3 digital_ldo_top_VIA4 $T=331310 56580 0 0 $X=331060 $Y=56350
X7916 3 digital_ldo_top_VIA4 $T=331310 60660 0 0 $X=331060 $Y=60430
X7917 3 digital_ldo_top_VIA4 $T=331310 64740 0 0 $X=331060 $Y=64510
X7918 3 digital_ldo_top_VIA4 $T=331310 68820 0 0 $X=331060 $Y=68590
X7919 3 digital_ldo_top_VIA4 $T=331310 72900 0 0 $X=331060 $Y=72670
X7920 3 digital_ldo_top_VIA4 $T=331310 76980 0 0 $X=331060 $Y=76750
X7921 3 digital_ldo_top_VIA4 $T=331310 81060 0 0 $X=331060 $Y=80830
X7922 3 digital_ldo_top_VIA4 $T=331310 85140 0 0 $X=331060 $Y=84910
X7923 3 digital_ldo_top_VIA4 $T=331310 89220 0 0 $X=331060 $Y=88990
X7924 3 digital_ldo_top_VIA4 $T=331310 93300 0 0 $X=331060 $Y=93070
X7925 3 digital_ldo_top_VIA4 $T=331310 97380 0 0 $X=331060 $Y=97150
X7926 3 digital_ldo_top_VIA4 $T=331310 101460 0 0 $X=331060 $Y=101230
X7927 3 digital_ldo_top_VIA4 $T=331310 105540 0 0 $X=331060 $Y=105310
X7928 3 digital_ldo_top_VIA4 $T=331310 109620 0 0 $X=331060 $Y=109390
X7929 3 digital_ldo_top_VIA4 $T=331310 113700 0 0 $X=331060 $Y=113470
X7930 3 digital_ldo_top_VIA4 $T=331310 117780 0 0 $X=331060 $Y=117550
X7931 3 digital_ldo_top_VIA4 $T=331310 121860 0 0 $X=331060 $Y=121630
X7932 3 digital_ldo_top_VIA4 $T=331310 125940 0 0 $X=331060 $Y=125710
X7933 2 digital_ldo_top_VIA4 $T=332690 13060 0 0 $X=332440 $Y=12830
X7934 2 digital_ldo_top_VIA4 $T=332690 49780 0 0 $X=332440 $Y=49550
X7935 2 digital_ldo_top_VIA4 $T=332690 53860 0 0 $X=332440 $Y=53630
X7936 2 digital_ldo_top_VIA4 $T=332690 57940 0 0 $X=332440 $Y=57710
X7937 2 digital_ldo_top_VIA4 $T=332690 62020 0 0 $X=332440 $Y=61790
X7938 2 digital_ldo_top_VIA4 $T=332690 66100 0 0 $X=332440 $Y=65870
X7939 2 digital_ldo_top_VIA4 $T=332690 70180 0 0 $X=332440 $Y=69950
X7940 2 digital_ldo_top_VIA4 $T=332690 74260 0 0 $X=332440 $Y=74030
X7941 2 digital_ldo_top_VIA4 $T=332690 78340 0 0 $X=332440 $Y=78110
X7942 2 digital_ldo_top_VIA4 $T=332690 82420 0 0 $X=332440 $Y=82190
X7943 2 digital_ldo_top_VIA4 $T=332690 86500 0 0 $X=332440 $Y=86270
X7944 2 digital_ldo_top_VIA4 $T=332690 90580 0 0 $X=332440 $Y=90350
X7945 2 digital_ldo_top_VIA4 $T=332690 94660 0 0 $X=332440 $Y=94430
X7946 2 digital_ldo_top_VIA4 $T=332690 98740 0 0 $X=332440 $Y=98510
X7947 2 digital_ldo_top_VIA4 $T=332690 102820 0 0 $X=332440 $Y=102590
X7948 2 digital_ldo_top_VIA4 $T=332690 106900 0 0 $X=332440 $Y=106670
X7949 2 digital_ldo_top_VIA4 $T=332690 110980 0 0 $X=332440 $Y=110750
X7950 2 digital_ldo_top_VIA4 $T=332690 115060 0 0 $X=332440 $Y=114830
X7951 2 digital_ldo_top_VIA4 $T=332690 119140 0 0 $X=332440 $Y=118910
X7952 2 digital_ldo_top_VIA4 $T=332690 123220 0 0 $X=332440 $Y=122990
X7953 2 digital_ldo_top_VIA4 $T=332690 127300 0 0 $X=332440 $Y=127070
X7954 3 digital_ldo_top_VIA4 $T=334990 11700 0 0 $X=334740 $Y=11470
X7955 3 digital_ldo_top_VIA4 $T=334990 52500 0 0 $X=334740 $Y=52270
X7956 3 digital_ldo_top_VIA4 $T=334990 56580 0 0 $X=334740 $Y=56350
X7957 3 digital_ldo_top_VIA4 $T=334990 60660 0 0 $X=334740 $Y=60430
X7958 3 digital_ldo_top_VIA4 $T=334990 64740 0 0 $X=334740 $Y=64510
X7959 3 digital_ldo_top_VIA4 $T=334990 68820 0 0 $X=334740 $Y=68590
X7960 3 digital_ldo_top_VIA4 $T=334990 72900 0 0 $X=334740 $Y=72670
X7961 3 digital_ldo_top_VIA4 $T=334990 76980 0 0 $X=334740 $Y=76750
X7962 3 digital_ldo_top_VIA4 $T=334990 81060 0 0 $X=334740 $Y=80830
X7963 3 digital_ldo_top_VIA4 $T=334990 85140 0 0 $X=334740 $Y=84910
X7964 3 digital_ldo_top_VIA4 $T=334990 89220 0 0 $X=334740 $Y=88990
X7965 3 digital_ldo_top_VIA4 $T=334990 93300 0 0 $X=334740 $Y=93070
X7966 3 digital_ldo_top_VIA4 $T=334990 97380 0 0 $X=334740 $Y=97150
X7967 3 digital_ldo_top_VIA4 $T=334990 101460 0 0 $X=334740 $Y=101230
X7968 3 digital_ldo_top_VIA4 $T=334990 105540 0 0 $X=334740 $Y=105310
X7969 3 digital_ldo_top_VIA4 $T=334990 109620 0 0 $X=334740 $Y=109390
X7970 3 digital_ldo_top_VIA4 $T=334990 113700 0 0 $X=334740 $Y=113470
X7971 3 digital_ldo_top_VIA4 $T=334990 117780 0 0 $X=334740 $Y=117550
X7972 3 digital_ldo_top_VIA4 $T=334990 121860 0 0 $X=334740 $Y=121630
X7973 3 digital_ldo_top_VIA4 $T=334990 125940 0 0 $X=334740 $Y=125710
X7974 2 digital_ldo_top_VIA4 $T=336370 13060 0 0 $X=336120 $Y=12830
X7975 2 digital_ldo_top_VIA4 $T=336370 49780 0 0 $X=336120 $Y=49550
X7976 2 digital_ldo_top_VIA4 $T=336370 53860 0 0 $X=336120 $Y=53630
X7977 2 digital_ldo_top_VIA4 $T=336370 57940 0 0 $X=336120 $Y=57710
X7978 2 digital_ldo_top_VIA4 $T=336370 62020 0 0 $X=336120 $Y=61790
X7979 2 digital_ldo_top_VIA4 $T=336370 66100 0 0 $X=336120 $Y=65870
X7980 2 digital_ldo_top_VIA4 $T=336370 70180 0 0 $X=336120 $Y=69950
X7981 2 digital_ldo_top_VIA4 $T=336370 74260 0 0 $X=336120 $Y=74030
X7982 2 digital_ldo_top_VIA4 $T=336370 78340 0 0 $X=336120 $Y=78110
X7983 2 digital_ldo_top_VIA4 $T=336370 82420 0 0 $X=336120 $Y=82190
X7984 2 digital_ldo_top_VIA4 $T=336370 86500 0 0 $X=336120 $Y=86270
X7985 2 digital_ldo_top_VIA4 $T=336370 90580 0 0 $X=336120 $Y=90350
X7986 2 digital_ldo_top_VIA4 $T=336370 94660 0 0 $X=336120 $Y=94430
X7987 2 digital_ldo_top_VIA4 $T=336370 98740 0 0 $X=336120 $Y=98510
X7988 2 digital_ldo_top_VIA4 $T=336370 102820 0 0 $X=336120 $Y=102590
X7989 2 digital_ldo_top_VIA4 $T=336370 106900 0 0 $X=336120 $Y=106670
X7990 2 digital_ldo_top_VIA4 $T=336370 110980 0 0 $X=336120 $Y=110750
X7991 2 digital_ldo_top_VIA4 $T=336370 115060 0 0 $X=336120 $Y=114830
X7992 2 digital_ldo_top_VIA4 $T=336370 119140 0 0 $X=336120 $Y=118910
X7993 2 digital_ldo_top_VIA4 $T=336370 123220 0 0 $X=336120 $Y=122990
X7994 2 digital_ldo_top_VIA4 $T=336370 127300 0 0 $X=336120 $Y=127070
X7995 3 digital_ldo_top_VIA4 $T=338670 11700 0 0 $X=338420 $Y=11470
X7996 3 digital_ldo_top_VIA4 $T=338670 52500 0 0 $X=338420 $Y=52270
X7997 3 digital_ldo_top_VIA4 $T=338670 56580 0 0 $X=338420 $Y=56350
X7998 3 digital_ldo_top_VIA4 $T=338670 60660 0 0 $X=338420 $Y=60430
X7999 3 digital_ldo_top_VIA4 $T=338670 64740 0 0 $X=338420 $Y=64510
X8000 3 digital_ldo_top_VIA4 $T=338670 68820 0 0 $X=338420 $Y=68590
X8001 3 digital_ldo_top_VIA4 $T=338670 72900 0 0 $X=338420 $Y=72670
X8002 3 digital_ldo_top_VIA4 $T=338670 76980 0 0 $X=338420 $Y=76750
X8003 3 digital_ldo_top_VIA4 $T=338670 81060 0 0 $X=338420 $Y=80830
X8004 3 digital_ldo_top_VIA4 $T=338670 85140 0 0 $X=338420 $Y=84910
X8005 3 digital_ldo_top_VIA4 $T=338670 89220 0 0 $X=338420 $Y=88990
X8006 3 digital_ldo_top_VIA4 $T=338670 93300 0 0 $X=338420 $Y=93070
X8007 3 digital_ldo_top_VIA4 $T=338670 97380 0 0 $X=338420 $Y=97150
X8008 3 digital_ldo_top_VIA4 $T=338670 101460 0 0 $X=338420 $Y=101230
X8009 3 digital_ldo_top_VIA4 $T=338670 105540 0 0 $X=338420 $Y=105310
X8010 3 digital_ldo_top_VIA4 $T=338670 109620 0 0 $X=338420 $Y=109390
X8011 3 digital_ldo_top_VIA4 $T=338670 113700 0 0 $X=338420 $Y=113470
X8012 3 digital_ldo_top_VIA4 $T=338670 117780 0 0 $X=338420 $Y=117550
X8013 3 digital_ldo_top_VIA4 $T=338670 121860 0 0 $X=338420 $Y=121630
X8014 3 digital_ldo_top_VIA4 $T=338670 125940 0 0 $X=338420 $Y=125710
X8015 2 digital_ldo_top_VIA4 $T=340050 13060 0 0 $X=339800 $Y=12830
X8016 2 digital_ldo_top_VIA4 $T=340050 49780 0 0 $X=339800 $Y=49550
X8017 2 digital_ldo_top_VIA4 $T=340050 53860 0 0 $X=339800 $Y=53630
X8018 2 digital_ldo_top_VIA4 $T=340050 57940 0 0 $X=339800 $Y=57710
X8019 2 digital_ldo_top_VIA4 $T=340050 62020 0 0 $X=339800 $Y=61790
X8020 2 digital_ldo_top_VIA4 $T=340050 66100 0 0 $X=339800 $Y=65870
X8021 2 digital_ldo_top_VIA4 $T=340050 70180 0 0 $X=339800 $Y=69950
X8022 2 digital_ldo_top_VIA4 $T=340050 74260 0 0 $X=339800 $Y=74030
X8023 2 digital_ldo_top_VIA4 $T=340050 78340 0 0 $X=339800 $Y=78110
X8024 2 digital_ldo_top_VIA4 $T=340050 82420 0 0 $X=339800 $Y=82190
X8025 2 digital_ldo_top_VIA4 $T=340050 86500 0 0 $X=339800 $Y=86270
X8026 2 digital_ldo_top_VIA4 $T=340050 90580 0 0 $X=339800 $Y=90350
X8027 2 digital_ldo_top_VIA4 $T=340050 94660 0 0 $X=339800 $Y=94430
X8028 2 digital_ldo_top_VIA4 $T=340050 98740 0 0 $X=339800 $Y=98510
X8029 2 digital_ldo_top_VIA4 $T=340050 102820 0 0 $X=339800 $Y=102590
X8030 2 digital_ldo_top_VIA4 $T=340050 106900 0 0 $X=339800 $Y=106670
X8031 2 digital_ldo_top_VIA4 $T=340050 110980 0 0 $X=339800 $Y=110750
X8032 2 digital_ldo_top_VIA4 $T=340050 115060 0 0 $X=339800 $Y=114830
X8033 2 digital_ldo_top_VIA4 $T=340050 119140 0 0 $X=339800 $Y=118910
X8034 2 digital_ldo_top_VIA4 $T=340050 123220 0 0 $X=339800 $Y=122990
X8035 2 digital_ldo_top_VIA4 $T=340050 127300 0 0 $X=339800 $Y=127070
X8036 3 digital_ldo_top_VIA4 $T=342350 11700 0 0 $X=342100 $Y=11470
X8037 3 digital_ldo_top_VIA4 $T=342350 52500 0 0 $X=342100 $Y=52270
X8038 3 digital_ldo_top_VIA4 $T=342350 56580 0 0 $X=342100 $Y=56350
X8039 3 digital_ldo_top_VIA4 $T=342350 60660 0 0 $X=342100 $Y=60430
X8040 3 digital_ldo_top_VIA4 $T=342350 64740 0 0 $X=342100 $Y=64510
X8041 3 digital_ldo_top_VIA4 $T=342350 68820 0 0 $X=342100 $Y=68590
X8042 3 digital_ldo_top_VIA4 $T=342350 72900 0 0 $X=342100 $Y=72670
X8043 3 digital_ldo_top_VIA4 $T=342350 76980 0 0 $X=342100 $Y=76750
X8044 3 digital_ldo_top_VIA4 $T=342350 81060 0 0 $X=342100 $Y=80830
X8045 3 digital_ldo_top_VIA4 $T=342350 85140 0 0 $X=342100 $Y=84910
X8046 3 digital_ldo_top_VIA4 $T=342350 89220 0 0 $X=342100 $Y=88990
X8047 3 digital_ldo_top_VIA4 $T=342350 93300 0 0 $X=342100 $Y=93070
X8048 3 digital_ldo_top_VIA4 $T=342350 97380 0 0 $X=342100 $Y=97150
X8049 3 digital_ldo_top_VIA4 $T=342350 101460 0 0 $X=342100 $Y=101230
X8050 3 digital_ldo_top_VIA4 $T=342350 105540 0 0 $X=342100 $Y=105310
X8051 3 digital_ldo_top_VIA4 $T=342350 109620 0 0 $X=342100 $Y=109390
X8052 3 digital_ldo_top_VIA4 $T=342350 113700 0 0 $X=342100 $Y=113470
X8053 3 digital_ldo_top_VIA4 $T=342350 117780 0 0 $X=342100 $Y=117550
X8054 3 digital_ldo_top_VIA4 $T=342350 121860 0 0 $X=342100 $Y=121630
X8055 3 digital_ldo_top_VIA4 $T=342350 125940 0 0 $X=342100 $Y=125710
X8056 2 digital_ldo_top_VIA4 $T=343730 13060 0 0 $X=343480 $Y=12830
X8057 2 digital_ldo_top_VIA4 $T=343730 49780 0 0 $X=343480 $Y=49550
X8058 2 digital_ldo_top_VIA4 $T=343730 53860 0 0 $X=343480 $Y=53630
X8059 2 digital_ldo_top_VIA4 $T=343730 57940 0 0 $X=343480 $Y=57710
X8060 2 digital_ldo_top_VIA4 $T=343730 62020 0 0 $X=343480 $Y=61790
X8061 2 digital_ldo_top_VIA4 $T=343730 66100 0 0 $X=343480 $Y=65870
X8062 2 digital_ldo_top_VIA4 $T=343730 70180 0 0 $X=343480 $Y=69950
X8063 2 digital_ldo_top_VIA4 $T=343730 74260 0 0 $X=343480 $Y=74030
X8064 2 digital_ldo_top_VIA4 $T=343730 78340 0 0 $X=343480 $Y=78110
X8065 2 digital_ldo_top_VIA4 $T=343730 82420 0 0 $X=343480 $Y=82190
X8066 2 digital_ldo_top_VIA4 $T=343730 86500 0 0 $X=343480 $Y=86270
X8067 2 digital_ldo_top_VIA4 $T=343730 90580 0 0 $X=343480 $Y=90350
X8068 2 digital_ldo_top_VIA4 $T=343730 94660 0 0 $X=343480 $Y=94430
X8069 2 digital_ldo_top_VIA4 $T=343730 98740 0 0 $X=343480 $Y=98510
X8070 2 digital_ldo_top_VIA4 $T=343730 102820 0 0 $X=343480 $Y=102590
X8071 2 digital_ldo_top_VIA4 $T=343730 106900 0 0 $X=343480 $Y=106670
X8072 2 digital_ldo_top_VIA4 $T=343730 110980 0 0 $X=343480 $Y=110750
X8073 2 digital_ldo_top_VIA4 $T=343730 115060 0 0 $X=343480 $Y=114830
X8074 2 digital_ldo_top_VIA4 $T=343730 119140 0 0 $X=343480 $Y=118910
X8075 2 digital_ldo_top_VIA4 $T=343730 123220 0 0 $X=343480 $Y=122990
X8076 2 digital_ldo_top_VIA4 $T=343730 127300 0 0 $X=343480 $Y=127070
X8077 3 digital_ldo_top_VIA4 $T=346030 11700 0 0 $X=345780 $Y=11470
X8078 3 digital_ldo_top_VIA4 $T=346030 52500 0 0 $X=345780 $Y=52270
X8079 3 digital_ldo_top_VIA4 $T=346030 56580 0 0 $X=345780 $Y=56350
X8080 3 digital_ldo_top_VIA4 $T=346030 60660 0 0 $X=345780 $Y=60430
X8081 3 digital_ldo_top_VIA4 $T=346030 64740 0 0 $X=345780 $Y=64510
X8082 3 digital_ldo_top_VIA4 $T=346030 68820 0 0 $X=345780 $Y=68590
X8083 3 digital_ldo_top_VIA4 $T=346030 72900 0 0 $X=345780 $Y=72670
X8084 3 digital_ldo_top_VIA4 $T=346030 76980 0 0 $X=345780 $Y=76750
X8085 3 digital_ldo_top_VIA4 $T=346030 81060 0 0 $X=345780 $Y=80830
X8086 3 digital_ldo_top_VIA4 $T=346030 85140 0 0 $X=345780 $Y=84910
X8087 3 digital_ldo_top_VIA4 $T=346030 89220 0 0 $X=345780 $Y=88990
X8088 3 digital_ldo_top_VIA4 $T=346030 93300 0 0 $X=345780 $Y=93070
X8089 3 digital_ldo_top_VIA4 $T=346030 97380 0 0 $X=345780 $Y=97150
X8090 3 digital_ldo_top_VIA4 $T=346030 101460 0 0 $X=345780 $Y=101230
X8091 3 digital_ldo_top_VIA4 $T=346030 105540 0 0 $X=345780 $Y=105310
X8092 3 digital_ldo_top_VIA4 $T=346030 109620 0 0 $X=345780 $Y=109390
X8093 3 digital_ldo_top_VIA4 $T=346030 113700 0 0 $X=345780 $Y=113470
X8094 3 digital_ldo_top_VIA4 $T=346030 117780 0 0 $X=345780 $Y=117550
X8095 3 digital_ldo_top_VIA4 $T=346030 121860 0 0 $X=345780 $Y=121630
X8096 3 digital_ldo_top_VIA4 $T=346030 125940 0 0 $X=345780 $Y=125710
X8097 2 digital_ldo_top_VIA4 $T=347410 13060 0 0 $X=347160 $Y=12830
X8098 2 digital_ldo_top_VIA4 $T=347410 49780 0 0 $X=347160 $Y=49550
X8099 2 digital_ldo_top_VIA4 $T=347410 53860 0 0 $X=347160 $Y=53630
X8100 2 digital_ldo_top_VIA4 $T=347410 57940 0 0 $X=347160 $Y=57710
X8101 2 digital_ldo_top_VIA4 $T=347410 62020 0 0 $X=347160 $Y=61790
X8102 2 digital_ldo_top_VIA4 $T=347410 66100 0 0 $X=347160 $Y=65870
X8103 2 digital_ldo_top_VIA4 $T=347410 70180 0 0 $X=347160 $Y=69950
X8104 2 digital_ldo_top_VIA4 $T=347410 74260 0 0 $X=347160 $Y=74030
X8105 2 digital_ldo_top_VIA4 $T=347410 78340 0 0 $X=347160 $Y=78110
X8106 2 digital_ldo_top_VIA4 $T=347410 82420 0 0 $X=347160 $Y=82190
X8107 2 digital_ldo_top_VIA4 $T=347410 86500 0 0 $X=347160 $Y=86270
X8108 2 digital_ldo_top_VIA4 $T=347410 90580 0 0 $X=347160 $Y=90350
X8109 2 digital_ldo_top_VIA4 $T=347410 94660 0 0 $X=347160 $Y=94430
X8110 2 digital_ldo_top_VIA4 $T=347410 98740 0 0 $X=347160 $Y=98510
X8111 2 digital_ldo_top_VIA4 $T=347410 102820 0 0 $X=347160 $Y=102590
X8112 2 digital_ldo_top_VIA4 $T=347410 106900 0 0 $X=347160 $Y=106670
X8113 2 digital_ldo_top_VIA4 $T=347410 110980 0 0 $X=347160 $Y=110750
X8114 2 digital_ldo_top_VIA4 $T=347410 115060 0 0 $X=347160 $Y=114830
X8115 2 digital_ldo_top_VIA4 $T=347410 119140 0 0 $X=347160 $Y=118910
X8116 2 digital_ldo_top_VIA4 $T=347410 123220 0 0 $X=347160 $Y=122990
X8117 2 digital_ldo_top_VIA4 $T=347410 127300 0 0 $X=347160 $Y=127070
X8118 3 digital_ldo_top_VIA4 $T=349710 11700 0 0 $X=349460 $Y=11470
X8119 3 digital_ldo_top_VIA4 $T=349710 52500 0 0 $X=349460 $Y=52270
X8120 3 digital_ldo_top_VIA4 $T=349710 56580 0 0 $X=349460 $Y=56350
X8121 3 digital_ldo_top_VIA4 $T=349710 60660 0 0 $X=349460 $Y=60430
X8122 3 digital_ldo_top_VIA4 $T=349710 64740 0 0 $X=349460 $Y=64510
X8123 3 digital_ldo_top_VIA4 $T=349710 68820 0 0 $X=349460 $Y=68590
X8124 3 digital_ldo_top_VIA4 $T=349710 72900 0 0 $X=349460 $Y=72670
X8125 3 digital_ldo_top_VIA4 $T=349710 76980 0 0 $X=349460 $Y=76750
X8126 3 digital_ldo_top_VIA4 $T=349710 81060 0 0 $X=349460 $Y=80830
X8127 3 digital_ldo_top_VIA4 $T=349710 85140 0 0 $X=349460 $Y=84910
X8128 3 digital_ldo_top_VIA4 $T=349710 89220 0 0 $X=349460 $Y=88990
X8129 3 digital_ldo_top_VIA4 $T=349710 93300 0 0 $X=349460 $Y=93070
X8130 3 digital_ldo_top_VIA4 $T=349710 97380 0 0 $X=349460 $Y=97150
X8131 3 digital_ldo_top_VIA4 $T=349710 101460 0 0 $X=349460 $Y=101230
X8132 3 digital_ldo_top_VIA4 $T=349710 105540 0 0 $X=349460 $Y=105310
X8133 3 digital_ldo_top_VIA4 $T=349710 109620 0 0 $X=349460 $Y=109390
X8134 3 digital_ldo_top_VIA4 $T=349710 113700 0 0 $X=349460 $Y=113470
X8135 3 digital_ldo_top_VIA4 $T=349710 117780 0 0 $X=349460 $Y=117550
X8136 3 digital_ldo_top_VIA4 $T=349710 121860 0 0 $X=349460 $Y=121630
X8137 3 digital_ldo_top_VIA4 $T=349710 125940 0 0 $X=349460 $Y=125710
X8138 2 digital_ldo_top_VIA4 $T=351090 13060 0 0 $X=350840 $Y=12830
X8139 2 digital_ldo_top_VIA4 $T=351090 17140 0 0 $X=350840 $Y=16910
X8140 2 digital_ldo_top_VIA4 $T=351090 21220 0 0 $X=350840 $Y=20990
X8141 2 digital_ldo_top_VIA4 $T=351090 25300 0 0 $X=350840 $Y=25070
X8142 2 digital_ldo_top_VIA4 $T=351090 29380 0 0 $X=350840 $Y=29150
X8143 2 digital_ldo_top_VIA4 $T=351090 33460 0 0 $X=350840 $Y=33230
X8144 2 digital_ldo_top_VIA4 $T=351090 37540 0 0 $X=350840 $Y=37310
X8145 2 digital_ldo_top_VIA4 $T=351090 41620 0 0 $X=350840 $Y=41390
X8146 2 digital_ldo_top_VIA4 $T=351090 45700 0 0 $X=350840 $Y=45470
X8147 2 digital_ldo_top_VIA4 $T=351090 49780 0 0 $X=350840 $Y=49550
X8148 2 digital_ldo_top_VIA4 $T=351090 53860 0 0 $X=350840 $Y=53630
X8149 2 digital_ldo_top_VIA4 $T=351090 57940 0 0 $X=350840 $Y=57710
X8150 2 digital_ldo_top_VIA4 $T=351090 62020 0 0 $X=350840 $Y=61790
X8151 2 digital_ldo_top_VIA4 $T=351090 66100 0 0 $X=350840 $Y=65870
X8152 2 digital_ldo_top_VIA4 $T=351090 70180 0 0 $X=350840 $Y=69950
X8153 2 digital_ldo_top_VIA4 $T=351090 74260 0 0 $X=350840 $Y=74030
X8154 2 digital_ldo_top_VIA4 $T=351090 78340 0 0 $X=350840 $Y=78110
X8155 2 digital_ldo_top_VIA4 $T=351090 82420 0 0 $X=350840 $Y=82190
X8156 2 digital_ldo_top_VIA4 $T=351090 86500 0 0 $X=350840 $Y=86270
X8157 2 digital_ldo_top_VIA4 $T=351090 90580 0 0 $X=350840 $Y=90350
X8158 2 digital_ldo_top_VIA4 $T=351090 94660 0 0 $X=350840 $Y=94430
X8159 2 digital_ldo_top_VIA4 $T=351090 98740 0 0 $X=350840 $Y=98510
X8160 2 digital_ldo_top_VIA4 $T=351090 102820 0 0 $X=350840 $Y=102590
X8161 2 digital_ldo_top_VIA4 $T=351090 106900 0 0 $X=350840 $Y=106670
X8162 2 digital_ldo_top_VIA4 $T=351090 110980 0 0 $X=350840 $Y=110750
X8163 2 digital_ldo_top_VIA4 $T=351090 115060 0 0 $X=350840 $Y=114830
X8164 2 digital_ldo_top_VIA4 $T=351090 119140 0 0 $X=350840 $Y=118910
X8165 2 digital_ldo_top_VIA4 $T=351090 123220 0 0 $X=350840 $Y=122990
X8166 2 digital_ldo_top_VIA4 $T=351090 127300 0 0 $X=350840 $Y=127070
X8167 3 digital_ldo_top_VIA4 $T=353390 11700 0 0 $X=353140 $Y=11470
X8168 3 digital_ldo_top_VIA4 $T=353390 15780 0 0 $X=353140 $Y=15550
X8169 3 digital_ldo_top_VIA4 $T=353390 19860 0 0 $X=353140 $Y=19630
X8170 3 digital_ldo_top_VIA4 $T=353390 23940 0 0 $X=353140 $Y=23710
X8171 3 digital_ldo_top_VIA4 $T=353390 28020 0 0 $X=353140 $Y=27790
X8172 3 digital_ldo_top_VIA4 $T=353390 32100 0 0 $X=353140 $Y=31870
X8173 3 digital_ldo_top_VIA4 $T=353390 36180 0 0 $X=353140 $Y=35950
X8174 3 digital_ldo_top_VIA4 $T=353390 40260 0 0 $X=353140 $Y=40030
X8175 3 digital_ldo_top_VIA4 $T=353390 44340 0 0 $X=353140 $Y=44110
X8176 3 digital_ldo_top_VIA4 $T=353390 48420 0 0 $X=353140 $Y=48190
X8177 3 digital_ldo_top_VIA4 $T=353390 52500 0 0 $X=353140 $Y=52270
X8178 3 digital_ldo_top_VIA4 $T=353390 56580 0 0 $X=353140 $Y=56350
X8179 3 digital_ldo_top_VIA4 $T=353390 60660 0 0 $X=353140 $Y=60430
X8180 3 digital_ldo_top_VIA4 $T=353390 64740 0 0 $X=353140 $Y=64510
X8181 3 digital_ldo_top_VIA4 $T=353390 68820 0 0 $X=353140 $Y=68590
X8182 3 digital_ldo_top_VIA4 $T=353390 72900 0 0 $X=353140 $Y=72670
X8183 3 digital_ldo_top_VIA4 $T=353390 76980 0 0 $X=353140 $Y=76750
X8184 3 digital_ldo_top_VIA4 $T=353390 81060 0 0 $X=353140 $Y=80830
X8185 3 digital_ldo_top_VIA4 $T=353390 85140 0 0 $X=353140 $Y=84910
X8186 3 digital_ldo_top_VIA4 $T=353390 89220 0 0 $X=353140 $Y=88990
X8187 3 digital_ldo_top_VIA4 $T=353390 93300 0 0 $X=353140 $Y=93070
X8188 3 digital_ldo_top_VIA4 $T=353390 97380 0 0 $X=353140 $Y=97150
X8189 3 digital_ldo_top_VIA4 $T=353390 101460 0 0 $X=353140 $Y=101230
X8190 3 digital_ldo_top_VIA4 $T=353390 105540 0 0 $X=353140 $Y=105310
X8191 3 digital_ldo_top_VIA4 $T=353390 109620 0 0 $X=353140 $Y=109390
X8192 3 digital_ldo_top_VIA4 $T=353390 113700 0 0 $X=353140 $Y=113470
X8193 3 digital_ldo_top_VIA4 $T=353390 117780 0 0 $X=353140 $Y=117550
X8194 3 digital_ldo_top_VIA4 $T=353390 121860 0 0 $X=353140 $Y=121630
X8195 3 digital_ldo_top_VIA4 $T=353390 125940 0 0 $X=353140 $Y=125710
X8196 2 digital_ldo_top_VIA4 $T=354770 13060 0 0 $X=354520 $Y=12830
X8197 2 digital_ldo_top_VIA4 $T=354770 17140 0 0 $X=354520 $Y=16910
X8198 2 digital_ldo_top_VIA4 $T=354770 21220 0 0 $X=354520 $Y=20990
X8199 2 digital_ldo_top_VIA4 $T=354770 25300 0 0 $X=354520 $Y=25070
X8200 2 digital_ldo_top_VIA4 $T=354770 29380 0 0 $X=354520 $Y=29150
X8201 2 digital_ldo_top_VIA4 $T=354770 33460 0 0 $X=354520 $Y=33230
X8202 2 digital_ldo_top_VIA4 $T=354770 37540 0 0 $X=354520 $Y=37310
X8203 2 digital_ldo_top_VIA4 $T=354770 41620 0 0 $X=354520 $Y=41390
X8204 2 digital_ldo_top_VIA4 $T=354770 45700 0 0 $X=354520 $Y=45470
X8205 2 digital_ldo_top_VIA4 $T=354770 49780 0 0 $X=354520 $Y=49550
X8206 2 digital_ldo_top_VIA4 $T=354770 53860 0 0 $X=354520 $Y=53630
X8207 2 digital_ldo_top_VIA4 $T=354770 57940 0 0 $X=354520 $Y=57710
X8208 2 digital_ldo_top_VIA4 $T=354770 62020 0 0 $X=354520 $Y=61790
X8209 2 digital_ldo_top_VIA4 $T=354770 66100 0 0 $X=354520 $Y=65870
X8210 2 digital_ldo_top_VIA4 $T=354770 70180 0 0 $X=354520 $Y=69950
X8211 2 digital_ldo_top_VIA4 $T=354770 74260 0 0 $X=354520 $Y=74030
X8212 2 digital_ldo_top_VIA4 $T=354770 78340 0 0 $X=354520 $Y=78110
X8213 2 digital_ldo_top_VIA4 $T=354770 82420 0 0 $X=354520 $Y=82190
X8214 2 digital_ldo_top_VIA4 $T=354770 86500 0 0 $X=354520 $Y=86270
X8215 2 digital_ldo_top_VIA4 $T=354770 90580 0 0 $X=354520 $Y=90350
X8216 2 digital_ldo_top_VIA4 $T=354770 94660 0 0 $X=354520 $Y=94430
X8217 2 digital_ldo_top_VIA4 $T=354770 98740 0 0 $X=354520 $Y=98510
X8218 2 digital_ldo_top_VIA4 $T=354770 102820 0 0 $X=354520 $Y=102590
X8219 2 digital_ldo_top_VIA4 $T=354770 106900 0 0 $X=354520 $Y=106670
X8220 2 digital_ldo_top_VIA4 $T=354770 110980 0 0 $X=354520 $Y=110750
X8221 2 digital_ldo_top_VIA4 $T=354770 115060 0 0 $X=354520 $Y=114830
X8222 2 digital_ldo_top_VIA4 $T=354770 119140 0 0 $X=354520 $Y=118910
X8223 2 digital_ldo_top_VIA4 $T=354770 123220 0 0 $X=354520 $Y=122990
X8224 2 digital_ldo_top_VIA4 $T=354770 127300 0 0 $X=354520 $Y=127070
X8225 3 digital_ldo_top_VIA4 $T=357070 11700 0 0 $X=356820 $Y=11470
X8226 3 digital_ldo_top_VIA4 $T=357070 15780 0 0 $X=356820 $Y=15550
X8227 3 digital_ldo_top_VIA4 $T=357070 19860 0 0 $X=356820 $Y=19630
X8228 3 digital_ldo_top_VIA4 $T=357070 23940 0 0 $X=356820 $Y=23710
X8229 3 digital_ldo_top_VIA4 $T=357070 28020 0 0 $X=356820 $Y=27790
X8230 3 digital_ldo_top_VIA4 $T=357070 32100 0 0 $X=356820 $Y=31870
X8231 3 digital_ldo_top_VIA4 $T=357070 36180 0 0 $X=356820 $Y=35950
X8232 3 digital_ldo_top_VIA4 $T=357070 40260 0 0 $X=356820 $Y=40030
X8233 3 digital_ldo_top_VIA4 $T=357070 44340 0 0 $X=356820 $Y=44110
X8234 3 digital_ldo_top_VIA4 $T=357070 48420 0 0 $X=356820 $Y=48190
X8235 3 digital_ldo_top_VIA4 $T=357070 52500 0 0 $X=356820 $Y=52270
X8236 3 digital_ldo_top_VIA4 $T=357070 56580 0 0 $X=356820 $Y=56350
X8237 3 digital_ldo_top_VIA4 $T=357070 60660 0 0 $X=356820 $Y=60430
X8238 3 digital_ldo_top_VIA4 $T=357070 64740 0 0 $X=356820 $Y=64510
X8239 3 digital_ldo_top_VIA4 $T=357070 68820 0 0 $X=356820 $Y=68590
X8240 3 digital_ldo_top_VIA4 $T=357070 72900 0 0 $X=356820 $Y=72670
X8241 3 digital_ldo_top_VIA4 $T=357070 76980 0 0 $X=356820 $Y=76750
X8242 3 digital_ldo_top_VIA4 $T=357070 81060 0 0 $X=356820 $Y=80830
X8243 3 digital_ldo_top_VIA4 $T=357070 85140 0 0 $X=356820 $Y=84910
X8244 3 digital_ldo_top_VIA4 $T=357070 89220 0 0 $X=356820 $Y=88990
X8245 3 digital_ldo_top_VIA4 $T=357070 93300 0 0 $X=356820 $Y=93070
X8246 3 digital_ldo_top_VIA4 $T=357070 97380 0 0 $X=356820 $Y=97150
X8247 3 digital_ldo_top_VIA4 $T=357070 101460 0 0 $X=356820 $Y=101230
X8248 3 digital_ldo_top_VIA4 $T=357070 105540 0 0 $X=356820 $Y=105310
X8249 3 digital_ldo_top_VIA4 $T=357070 109620 0 0 $X=356820 $Y=109390
X8250 3 digital_ldo_top_VIA4 $T=357070 113700 0 0 $X=356820 $Y=113470
X8251 3 digital_ldo_top_VIA4 $T=357070 117780 0 0 $X=356820 $Y=117550
X8252 3 digital_ldo_top_VIA4 $T=357070 121860 0 0 $X=356820 $Y=121630
X8253 3 digital_ldo_top_VIA4 $T=357070 125940 0 0 $X=356820 $Y=125710
X8254 2 digital_ldo_top_VIA4 $T=358450 13060 0 0 $X=358200 $Y=12830
X8255 2 digital_ldo_top_VIA4 $T=358450 17140 0 0 $X=358200 $Y=16910
X8256 2 digital_ldo_top_VIA4 $T=358450 21220 0 0 $X=358200 $Y=20990
X8257 2 digital_ldo_top_VIA4 $T=358450 25300 0 0 $X=358200 $Y=25070
X8258 2 digital_ldo_top_VIA4 $T=358450 29380 0 0 $X=358200 $Y=29150
X8259 2 digital_ldo_top_VIA4 $T=358450 33460 0 0 $X=358200 $Y=33230
X8260 2 digital_ldo_top_VIA4 $T=358450 37540 0 0 $X=358200 $Y=37310
X8261 2 digital_ldo_top_VIA4 $T=358450 41620 0 0 $X=358200 $Y=41390
X8262 2 digital_ldo_top_VIA4 $T=358450 45700 0 0 $X=358200 $Y=45470
X8263 2 digital_ldo_top_VIA4 $T=358450 49780 0 0 $X=358200 $Y=49550
X8264 2 digital_ldo_top_VIA4 $T=358450 53860 0 0 $X=358200 $Y=53630
X8265 2 digital_ldo_top_VIA4 $T=358450 57940 0 0 $X=358200 $Y=57710
X8266 2 digital_ldo_top_VIA4 $T=358450 62020 0 0 $X=358200 $Y=61790
X8267 2 digital_ldo_top_VIA4 $T=358450 66100 0 0 $X=358200 $Y=65870
X8268 2 digital_ldo_top_VIA4 $T=358450 70180 0 0 $X=358200 $Y=69950
X8269 2 digital_ldo_top_VIA4 $T=358450 74260 0 0 $X=358200 $Y=74030
X8270 2 digital_ldo_top_VIA4 $T=358450 78340 0 0 $X=358200 $Y=78110
X8271 2 digital_ldo_top_VIA4 $T=358450 82420 0 0 $X=358200 $Y=82190
X8272 2 digital_ldo_top_VIA4 $T=358450 86500 0 0 $X=358200 $Y=86270
X8273 2 digital_ldo_top_VIA4 $T=358450 90580 0 0 $X=358200 $Y=90350
X8274 2 digital_ldo_top_VIA4 $T=358450 94660 0 0 $X=358200 $Y=94430
X8275 2 digital_ldo_top_VIA4 $T=358450 98740 0 0 $X=358200 $Y=98510
X8276 2 digital_ldo_top_VIA4 $T=358450 102820 0 0 $X=358200 $Y=102590
X8277 2 digital_ldo_top_VIA4 $T=358450 106900 0 0 $X=358200 $Y=106670
X8278 2 digital_ldo_top_VIA4 $T=358450 110980 0 0 $X=358200 $Y=110750
X8279 2 digital_ldo_top_VIA4 $T=358450 115060 0 0 $X=358200 $Y=114830
X8280 2 digital_ldo_top_VIA4 $T=358450 119140 0 0 $X=358200 $Y=118910
X8281 2 digital_ldo_top_VIA4 $T=358450 123220 0 0 $X=358200 $Y=122990
X8282 2 digital_ldo_top_VIA4 $T=358450 127300 0 0 $X=358200 $Y=127070
X8283 3 digital_ldo_top_VIA4 $T=360750 11700 0 0 $X=360500 $Y=11470
X8284 3 digital_ldo_top_VIA4 $T=360750 15780 0 0 $X=360500 $Y=15550
X8285 3 digital_ldo_top_VIA4 $T=360750 19860 0 0 $X=360500 $Y=19630
X8286 3 digital_ldo_top_VIA4 $T=360750 23940 0 0 $X=360500 $Y=23710
X8287 3 digital_ldo_top_VIA4 $T=360750 28020 0 0 $X=360500 $Y=27790
X8288 3 digital_ldo_top_VIA4 $T=360750 32100 0 0 $X=360500 $Y=31870
X8289 3 digital_ldo_top_VIA4 $T=360750 36180 0 0 $X=360500 $Y=35950
X8290 3 digital_ldo_top_VIA4 $T=360750 40260 0 0 $X=360500 $Y=40030
X8291 3 digital_ldo_top_VIA4 $T=360750 44340 0 0 $X=360500 $Y=44110
X8292 3 digital_ldo_top_VIA4 $T=360750 48420 0 0 $X=360500 $Y=48190
X8293 3 digital_ldo_top_VIA4 $T=360750 52500 0 0 $X=360500 $Y=52270
X8294 3 digital_ldo_top_VIA4 $T=360750 56580 0 0 $X=360500 $Y=56350
X8295 3 digital_ldo_top_VIA4 $T=360750 60660 0 0 $X=360500 $Y=60430
X8296 3 digital_ldo_top_VIA4 $T=360750 64740 0 0 $X=360500 $Y=64510
X8297 3 digital_ldo_top_VIA4 $T=360750 68820 0 0 $X=360500 $Y=68590
X8298 3 digital_ldo_top_VIA4 $T=360750 72900 0 0 $X=360500 $Y=72670
X8299 3 digital_ldo_top_VIA4 $T=360750 76980 0 0 $X=360500 $Y=76750
X8300 3 digital_ldo_top_VIA4 $T=360750 81060 0 0 $X=360500 $Y=80830
X8301 3 digital_ldo_top_VIA4 $T=360750 85140 0 0 $X=360500 $Y=84910
X8302 3 digital_ldo_top_VIA4 $T=360750 89220 0 0 $X=360500 $Y=88990
X8303 3 digital_ldo_top_VIA4 $T=360750 93300 0 0 $X=360500 $Y=93070
X8304 3 digital_ldo_top_VIA4 $T=360750 97380 0 0 $X=360500 $Y=97150
X8305 3 digital_ldo_top_VIA4 $T=360750 101460 0 0 $X=360500 $Y=101230
X8306 3 digital_ldo_top_VIA4 $T=360750 105540 0 0 $X=360500 $Y=105310
X8307 3 digital_ldo_top_VIA4 $T=360750 109620 0 0 $X=360500 $Y=109390
X8308 3 digital_ldo_top_VIA4 $T=360750 113700 0 0 $X=360500 $Y=113470
X8309 3 digital_ldo_top_VIA4 $T=360750 117780 0 0 $X=360500 $Y=117550
X8310 3 digital_ldo_top_VIA4 $T=360750 121860 0 0 $X=360500 $Y=121630
X8311 3 digital_ldo_top_VIA4 $T=360750 125940 0 0 $X=360500 $Y=125710
X8312 2 digital_ldo_top_VIA4 $T=362130 13060 0 0 $X=361880 $Y=12830
X8313 2 digital_ldo_top_VIA4 $T=362130 17140 0 0 $X=361880 $Y=16910
X8314 2 digital_ldo_top_VIA4 $T=362130 21220 0 0 $X=361880 $Y=20990
X8315 2 digital_ldo_top_VIA4 $T=362130 25300 0 0 $X=361880 $Y=25070
X8316 2 digital_ldo_top_VIA4 $T=362130 29380 0 0 $X=361880 $Y=29150
X8317 2 digital_ldo_top_VIA4 $T=362130 33460 0 0 $X=361880 $Y=33230
X8318 2 digital_ldo_top_VIA4 $T=362130 37540 0 0 $X=361880 $Y=37310
X8319 2 digital_ldo_top_VIA4 $T=362130 41620 0 0 $X=361880 $Y=41390
X8320 2 digital_ldo_top_VIA4 $T=362130 45700 0 0 $X=361880 $Y=45470
X8321 2 digital_ldo_top_VIA4 $T=362130 49780 0 0 $X=361880 $Y=49550
X8322 2 digital_ldo_top_VIA4 $T=362130 53860 0 0 $X=361880 $Y=53630
X8323 2 digital_ldo_top_VIA4 $T=362130 57940 0 0 $X=361880 $Y=57710
X8324 2 digital_ldo_top_VIA4 $T=362130 62020 0 0 $X=361880 $Y=61790
X8325 2 digital_ldo_top_VIA4 $T=362130 66100 0 0 $X=361880 $Y=65870
X8326 2 digital_ldo_top_VIA4 $T=362130 70180 0 0 $X=361880 $Y=69950
X8327 2 digital_ldo_top_VIA4 $T=362130 74260 0 0 $X=361880 $Y=74030
X8328 2 digital_ldo_top_VIA4 $T=362130 78340 0 0 $X=361880 $Y=78110
X8329 2 digital_ldo_top_VIA4 $T=362130 82420 0 0 $X=361880 $Y=82190
X8330 2 digital_ldo_top_VIA4 $T=362130 86500 0 0 $X=361880 $Y=86270
X8331 2 digital_ldo_top_VIA4 $T=362130 90580 0 0 $X=361880 $Y=90350
X8332 2 digital_ldo_top_VIA4 $T=362130 94660 0 0 $X=361880 $Y=94430
X8333 2 digital_ldo_top_VIA4 $T=362130 98740 0 0 $X=361880 $Y=98510
X8334 2 digital_ldo_top_VIA4 $T=362130 102820 0 0 $X=361880 $Y=102590
X8335 2 digital_ldo_top_VIA4 $T=362130 106900 0 0 $X=361880 $Y=106670
X8336 2 digital_ldo_top_VIA4 $T=362130 110980 0 0 $X=361880 $Y=110750
X8337 2 digital_ldo_top_VIA4 $T=362130 115060 0 0 $X=361880 $Y=114830
X8338 2 digital_ldo_top_VIA4 $T=362130 119140 0 0 $X=361880 $Y=118910
X8339 2 digital_ldo_top_VIA4 $T=362130 123220 0 0 $X=361880 $Y=122990
X8340 2 digital_ldo_top_VIA4 $T=362130 127300 0 0 $X=361880 $Y=127070
X8341 3 digital_ldo_top_VIA4 $T=364430 11700 0 0 $X=364180 $Y=11470
X8342 3 digital_ldo_top_VIA4 $T=364430 15780 0 0 $X=364180 $Y=15550
X8343 3 digital_ldo_top_VIA4 $T=364430 19860 0 0 $X=364180 $Y=19630
X8344 3 digital_ldo_top_VIA4 $T=364430 23940 0 0 $X=364180 $Y=23710
X8345 3 digital_ldo_top_VIA4 $T=364430 28020 0 0 $X=364180 $Y=27790
X8346 3 digital_ldo_top_VIA4 $T=364430 32100 0 0 $X=364180 $Y=31870
X8347 3 digital_ldo_top_VIA4 $T=364430 36180 0 0 $X=364180 $Y=35950
X8348 3 digital_ldo_top_VIA4 $T=364430 40260 0 0 $X=364180 $Y=40030
X8349 3 digital_ldo_top_VIA4 $T=364430 44340 0 0 $X=364180 $Y=44110
X8350 3 digital_ldo_top_VIA4 $T=364430 48420 0 0 $X=364180 $Y=48190
X8351 3 digital_ldo_top_VIA4 $T=364430 52500 0 0 $X=364180 $Y=52270
X8352 3 digital_ldo_top_VIA4 $T=364430 56580 0 0 $X=364180 $Y=56350
X8353 3 digital_ldo_top_VIA4 $T=364430 60660 0 0 $X=364180 $Y=60430
X8354 3 digital_ldo_top_VIA4 $T=364430 64740 0 0 $X=364180 $Y=64510
X8355 3 digital_ldo_top_VIA4 $T=364430 68820 0 0 $X=364180 $Y=68590
X8356 3 digital_ldo_top_VIA4 $T=364430 72900 0 0 $X=364180 $Y=72670
X8357 3 digital_ldo_top_VIA4 $T=364430 76980 0 0 $X=364180 $Y=76750
X8358 3 digital_ldo_top_VIA4 $T=364430 81060 0 0 $X=364180 $Y=80830
X8359 3 digital_ldo_top_VIA4 $T=364430 85140 0 0 $X=364180 $Y=84910
X8360 3 digital_ldo_top_VIA4 $T=364430 89220 0 0 $X=364180 $Y=88990
X8361 3 digital_ldo_top_VIA4 $T=364430 93300 0 0 $X=364180 $Y=93070
X8362 3 digital_ldo_top_VIA4 $T=364430 97380 0 0 $X=364180 $Y=97150
X8363 3 digital_ldo_top_VIA4 $T=364430 101460 0 0 $X=364180 $Y=101230
X8364 3 digital_ldo_top_VIA4 $T=364430 105540 0 0 $X=364180 $Y=105310
X8365 3 digital_ldo_top_VIA4 $T=364430 109620 0 0 $X=364180 $Y=109390
X8366 3 digital_ldo_top_VIA4 $T=364430 113700 0 0 $X=364180 $Y=113470
X8367 3 digital_ldo_top_VIA4 $T=364430 117780 0 0 $X=364180 $Y=117550
X8368 3 digital_ldo_top_VIA4 $T=364430 121860 0 0 $X=364180 $Y=121630
X8369 3 digital_ldo_top_VIA4 $T=364430 125940 0 0 $X=364180 $Y=125710
X8370 2 digital_ldo_top_VIA4 $T=365810 13060 0 0 $X=365560 $Y=12830
X8371 2 digital_ldo_top_VIA4 $T=365810 17140 0 0 $X=365560 $Y=16910
X8372 2 digital_ldo_top_VIA4 $T=365810 21220 0 0 $X=365560 $Y=20990
X8373 2 digital_ldo_top_VIA4 $T=365810 25300 0 0 $X=365560 $Y=25070
X8374 2 digital_ldo_top_VIA4 $T=365810 29380 0 0 $X=365560 $Y=29150
X8375 2 digital_ldo_top_VIA4 $T=365810 33460 0 0 $X=365560 $Y=33230
X8376 2 digital_ldo_top_VIA4 $T=365810 37540 0 0 $X=365560 $Y=37310
X8377 2 digital_ldo_top_VIA4 $T=365810 41620 0 0 $X=365560 $Y=41390
X8378 2 digital_ldo_top_VIA4 $T=365810 45700 0 0 $X=365560 $Y=45470
X8379 2 digital_ldo_top_VIA4 $T=365810 49780 0 0 $X=365560 $Y=49550
X8380 2 digital_ldo_top_VIA4 $T=365810 53860 0 0 $X=365560 $Y=53630
X8381 2 digital_ldo_top_VIA4 $T=365810 57940 0 0 $X=365560 $Y=57710
X8382 2 digital_ldo_top_VIA4 $T=365810 62020 0 0 $X=365560 $Y=61790
X8383 2 digital_ldo_top_VIA4 $T=365810 66100 0 0 $X=365560 $Y=65870
X8384 2 digital_ldo_top_VIA4 $T=365810 70180 0 0 $X=365560 $Y=69950
X8385 2 digital_ldo_top_VIA4 $T=365810 74260 0 0 $X=365560 $Y=74030
X8386 2 digital_ldo_top_VIA4 $T=365810 78340 0 0 $X=365560 $Y=78110
X8387 2 digital_ldo_top_VIA4 $T=365810 82420 0 0 $X=365560 $Y=82190
X8388 2 digital_ldo_top_VIA4 $T=365810 86500 0 0 $X=365560 $Y=86270
X8389 2 digital_ldo_top_VIA4 $T=365810 90580 0 0 $X=365560 $Y=90350
X8390 2 digital_ldo_top_VIA4 $T=365810 94660 0 0 $X=365560 $Y=94430
X8391 2 digital_ldo_top_VIA4 $T=365810 98740 0 0 $X=365560 $Y=98510
X8392 2 digital_ldo_top_VIA4 $T=365810 102820 0 0 $X=365560 $Y=102590
X8393 2 digital_ldo_top_VIA4 $T=365810 106900 0 0 $X=365560 $Y=106670
X8394 2 digital_ldo_top_VIA4 $T=365810 110980 0 0 $X=365560 $Y=110750
X8395 2 digital_ldo_top_VIA4 $T=365810 115060 0 0 $X=365560 $Y=114830
X8396 2 digital_ldo_top_VIA4 $T=365810 119140 0 0 $X=365560 $Y=118910
X8397 2 digital_ldo_top_VIA4 $T=365810 123220 0 0 $X=365560 $Y=122990
X8398 2 digital_ldo_top_VIA4 $T=365810 127300 0 0 $X=365560 $Y=127070
X8399 3 digital_ldo_top_VIA4 $T=368110 11700 0 0 $X=367860 $Y=11470
X8400 3 digital_ldo_top_VIA4 $T=368110 15780 0 0 $X=367860 $Y=15550
X8401 3 digital_ldo_top_VIA4 $T=368110 19860 0 0 $X=367860 $Y=19630
X8402 3 digital_ldo_top_VIA4 $T=368110 23940 0 0 $X=367860 $Y=23710
X8403 3 digital_ldo_top_VIA4 $T=368110 28020 0 0 $X=367860 $Y=27790
X8404 3 digital_ldo_top_VIA4 $T=368110 32100 0 0 $X=367860 $Y=31870
X8405 3 digital_ldo_top_VIA4 $T=368110 36180 0 0 $X=367860 $Y=35950
X8406 3 digital_ldo_top_VIA4 $T=368110 40260 0 0 $X=367860 $Y=40030
X8407 3 digital_ldo_top_VIA4 $T=368110 44340 0 0 $X=367860 $Y=44110
X8408 3 digital_ldo_top_VIA4 $T=368110 48420 0 0 $X=367860 $Y=48190
X8409 3 digital_ldo_top_VIA4 $T=368110 52500 0 0 $X=367860 $Y=52270
X8410 3 digital_ldo_top_VIA4 $T=368110 56580 0 0 $X=367860 $Y=56350
X8411 3 digital_ldo_top_VIA4 $T=368110 60660 0 0 $X=367860 $Y=60430
X8412 3 digital_ldo_top_VIA4 $T=368110 64740 0 0 $X=367860 $Y=64510
X8413 3 digital_ldo_top_VIA4 $T=368110 68820 0 0 $X=367860 $Y=68590
X8414 3 digital_ldo_top_VIA4 $T=368110 72900 0 0 $X=367860 $Y=72670
X8415 3 digital_ldo_top_VIA4 $T=368110 76980 0 0 $X=367860 $Y=76750
X8416 3 digital_ldo_top_VIA4 $T=368110 81060 0 0 $X=367860 $Y=80830
X8417 3 digital_ldo_top_VIA4 $T=368110 85140 0 0 $X=367860 $Y=84910
X8418 3 digital_ldo_top_VIA4 $T=368110 89220 0 0 $X=367860 $Y=88990
X8419 3 digital_ldo_top_VIA4 $T=368110 93300 0 0 $X=367860 $Y=93070
X8420 3 digital_ldo_top_VIA4 $T=368110 97380 0 0 $X=367860 $Y=97150
X8421 3 digital_ldo_top_VIA4 $T=368110 101460 0 0 $X=367860 $Y=101230
X8422 3 digital_ldo_top_VIA4 $T=368110 105540 0 0 $X=367860 $Y=105310
X8423 3 digital_ldo_top_VIA4 $T=368110 109620 0 0 $X=367860 $Y=109390
X8424 3 digital_ldo_top_VIA4 $T=368110 113700 0 0 $X=367860 $Y=113470
X8425 3 digital_ldo_top_VIA4 $T=368110 117780 0 0 $X=367860 $Y=117550
X8426 3 digital_ldo_top_VIA4 $T=368110 121860 0 0 $X=367860 $Y=121630
X8427 3 digital_ldo_top_VIA4 $T=368110 125940 0 0 $X=367860 $Y=125710
X8428 2 digital_ldo_top_VIA4 $T=369490 13060 0 0 $X=369240 $Y=12830
X8429 2 digital_ldo_top_VIA4 $T=369490 17140 0 0 $X=369240 $Y=16910
X8430 2 digital_ldo_top_VIA4 $T=369490 21220 0 0 $X=369240 $Y=20990
X8431 2 digital_ldo_top_VIA4 $T=369490 25300 0 0 $X=369240 $Y=25070
X8432 2 digital_ldo_top_VIA4 $T=369490 29380 0 0 $X=369240 $Y=29150
X8433 2 digital_ldo_top_VIA4 $T=369490 33460 0 0 $X=369240 $Y=33230
X8434 2 digital_ldo_top_VIA4 $T=369490 37540 0 0 $X=369240 $Y=37310
X8435 2 digital_ldo_top_VIA4 $T=369490 41620 0 0 $X=369240 $Y=41390
X8436 2 digital_ldo_top_VIA4 $T=369490 45700 0 0 $X=369240 $Y=45470
X8437 2 digital_ldo_top_VIA4 $T=369490 49780 0 0 $X=369240 $Y=49550
X8438 2 digital_ldo_top_VIA4 $T=369490 53860 0 0 $X=369240 $Y=53630
X8439 2 digital_ldo_top_VIA4 $T=369490 57940 0 0 $X=369240 $Y=57710
X8440 2 digital_ldo_top_VIA4 $T=369490 62020 0 0 $X=369240 $Y=61790
X8441 2 digital_ldo_top_VIA4 $T=369490 66100 0 0 $X=369240 $Y=65870
X8442 2 digital_ldo_top_VIA4 $T=369490 70180 0 0 $X=369240 $Y=69950
X8443 2 digital_ldo_top_VIA4 $T=369490 74260 0 0 $X=369240 $Y=74030
X8444 2 digital_ldo_top_VIA4 $T=369490 78340 0 0 $X=369240 $Y=78110
X8445 2 digital_ldo_top_VIA4 $T=369490 82420 0 0 $X=369240 $Y=82190
X8446 2 digital_ldo_top_VIA4 $T=369490 86500 0 0 $X=369240 $Y=86270
X8447 2 digital_ldo_top_VIA4 $T=369490 90580 0 0 $X=369240 $Y=90350
X8448 2 digital_ldo_top_VIA4 $T=369490 94660 0 0 $X=369240 $Y=94430
X8449 2 digital_ldo_top_VIA4 $T=369490 98740 0 0 $X=369240 $Y=98510
X8450 2 digital_ldo_top_VIA4 $T=369490 102820 0 0 $X=369240 $Y=102590
X8451 2 digital_ldo_top_VIA4 $T=369490 106900 0 0 $X=369240 $Y=106670
X8452 2 digital_ldo_top_VIA4 $T=369490 110980 0 0 $X=369240 $Y=110750
X8453 2 digital_ldo_top_VIA4 $T=369490 115060 0 0 $X=369240 $Y=114830
X8454 2 digital_ldo_top_VIA4 $T=369490 119140 0 0 $X=369240 $Y=118910
X8455 2 digital_ldo_top_VIA4 $T=369490 123220 0 0 $X=369240 $Y=122990
X8456 2 digital_ldo_top_VIA4 $T=369490 127300 0 0 $X=369240 $Y=127070
X8457 3 digital_ldo_top_VIA4 $T=371790 11700 0 0 $X=371540 $Y=11470
X8458 3 digital_ldo_top_VIA4 $T=371790 15780 0 0 $X=371540 $Y=15550
X8459 3 digital_ldo_top_VIA4 $T=371790 19860 0 0 $X=371540 $Y=19630
X8460 3 digital_ldo_top_VIA4 $T=371790 23940 0 0 $X=371540 $Y=23710
X8461 3 digital_ldo_top_VIA4 $T=371790 28020 0 0 $X=371540 $Y=27790
X8462 3 digital_ldo_top_VIA4 $T=371790 32100 0 0 $X=371540 $Y=31870
X8463 3 digital_ldo_top_VIA4 $T=371790 36180 0 0 $X=371540 $Y=35950
X8464 3 digital_ldo_top_VIA4 $T=371790 40260 0 0 $X=371540 $Y=40030
X8465 3 digital_ldo_top_VIA4 $T=371790 44340 0 0 $X=371540 $Y=44110
X8466 3 digital_ldo_top_VIA4 $T=371790 48420 0 0 $X=371540 $Y=48190
X8467 3 digital_ldo_top_VIA4 $T=371790 52500 0 0 $X=371540 $Y=52270
X8468 3 digital_ldo_top_VIA4 $T=371790 56580 0 0 $X=371540 $Y=56350
X8469 3 digital_ldo_top_VIA4 $T=371790 60660 0 0 $X=371540 $Y=60430
X8470 3 digital_ldo_top_VIA4 $T=371790 64740 0 0 $X=371540 $Y=64510
X8471 3 digital_ldo_top_VIA4 $T=371790 68820 0 0 $X=371540 $Y=68590
X8472 3 digital_ldo_top_VIA4 $T=371790 72900 0 0 $X=371540 $Y=72670
X8473 3 digital_ldo_top_VIA4 $T=371790 76980 0 0 $X=371540 $Y=76750
X8474 3 digital_ldo_top_VIA4 $T=371790 81060 0 0 $X=371540 $Y=80830
X8475 3 digital_ldo_top_VIA4 $T=371790 85140 0 0 $X=371540 $Y=84910
X8476 3 digital_ldo_top_VIA4 $T=371790 89220 0 0 $X=371540 $Y=88990
X8477 3 digital_ldo_top_VIA4 $T=371790 93300 0 0 $X=371540 $Y=93070
X8478 3 digital_ldo_top_VIA4 $T=371790 97380 0 0 $X=371540 $Y=97150
X8479 3 digital_ldo_top_VIA4 $T=371790 101460 0 0 $X=371540 $Y=101230
X8480 3 digital_ldo_top_VIA4 $T=371790 105540 0 0 $X=371540 $Y=105310
X8481 3 digital_ldo_top_VIA4 $T=371790 109620 0 0 $X=371540 $Y=109390
X8482 3 digital_ldo_top_VIA4 $T=371790 113700 0 0 $X=371540 $Y=113470
X8483 3 digital_ldo_top_VIA4 $T=371790 117780 0 0 $X=371540 $Y=117550
X8484 3 digital_ldo_top_VIA4 $T=371790 121860 0 0 $X=371540 $Y=121630
X8485 3 digital_ldo_top_VIA4 $T=371790 125940 0 0 $X=371540 $Y=125710
X8486 2 digital_ldo_top_VIA4 $T=373170 13060 0 0 $X=372920 $Y=12830
X8487 2 digital_ldo_top_VIA4 $T=373170 17140 0 0 $X=372920 $Y=16910
X8488 2 digital_ldo_top_VIA4 $T=373170 21220 0 0 $X=372920 $Y=20990
X8489 2 digital_ldo_top_VIA4 $T=373170 25300 0 0 $X=372920 $Y=25070
X8490 2 digital_ldo_top_VIA4 $T=373170 29380 0 0 $X=372920 $Y=29150
X8491 2 digital_ldo_top_VIA4 $T=373170 33460 0 0 $X=372920 $Y=33230
X8492 2 digital_ldo_top_VIA4 $T=373170 37540 0 0 $X=372920 $Y=37310
X8493 2 digital_ldo_top_VIA4 $T=373170 41620 0 0 $X=372920 $Y=41390
X8494 2 digital_ldo_top_VIA4 $T=373170 45700 0 0 $X=372920 $Y=45470
X8495 2 digital_ldo_top_VIA4 $T=373170 49780 0 0 $X=372920 $Y=49550
X8496 2 digital_ldo_top_VIA4 $T=373170 53860 0 0 $X=372920 $Y=53630
X8497 2 digital_ldo_top_VIA4 $T=373170 57940 0 0 $X=372920 $Y=57710
X8498 2 digital_ldo_top_VIA4 $T=373170 62020 0 0 $X=372920 $Y=61790
X8499 2 digital_ldo_top_VIA4 $T=373170 66100 0 0 $X=372920 $Y=65870
X8500 2 digital_ldo_top_VIA4 $T=373170 70180 0 0 $X=372920 $Y=69950
X8501 2 digital_ldo_top_VIA4 $T=373170 74260 0 0 $X=372920 $Y=74030
X8502 2 digital_ldo_top_VIA4 $T=373170 78340 0 0 $X=372920 $Y=78110
X8503 2 digital_ldo_top_VIA4 $T=373170 82420 0 0 $X=372920 $Y=82190
X8504 2 digital_ldo_top_VIA4 $T=373170 86500 0 0 $X=372920 $Y=86270
X8505 2 digital_ldo_top_VIA4 $T=373170 90580 0 0 $X=372920 $Y=90350
X8506 2 digital_ldo_top_VIA4 $T=373170 94660 0 0 $X=372920 $Y=94430
X8507 2 digital_ldo_top_VIA4 $T=373170 98740 0 0 $X=372920 $Y=98510
X8508 2 digital_ldo_top_VIA4 $T=373170 102820 0 0 $X=372920 $Y=102590
X8509 2 digital_ldo_top_VIA4 $T=373170 106900 0 0 $X=372920 $Y=106670
X8510 2 digital_ldo_top_VIA4 $T=373170 110980 0 0 $X=372920 $Y=110750
X8511 2 digital_ldo_top_VIA4 $T=373170 115060 0 0 $X=372920 $Y=114830
X8512 2 digital_ldo_top_VIA4 $T=373170 119140 0 0 $X=372920 $Y=118910
X8513 2 digital_ldo_top_VIA4 $T=373170 123220 0 0 $X=372920 $Y=122990
X8514 2 digital_ldo_top_VIA4 $T=373170 127300 0 0 $X=372920 $Y=127070
X8515 3 digital_ldo_top_VIA4 $T=375470 11700 0 0 $X=375220 $Y=11470
X8516 3 digital_ldo_top_VIA4 $T=375470 15780 0 0 $X=375220 $Y=15550
X8517 3 digital_ldo_top_VIA4 $T=375470 19860 0 0 $X=375220 $Y=19630
X8518 3 digital_ldo_top_VIA4 $T=375470 23940 0 0 $X=375220 $Y=23710
X8519 3 digital_ldo_top_VIA4 $T=375470 28020 0 0 $X=375220 $Y=27790
X8520 3 digital_ldo_top_VIA4 $T=375470 32100 0 0 $X=375220 $Y=31870
X8521 3 digital_ldo_top_VIA4 $T=375470 36180 0 0 $X=375220 $Y=35950
X8522 3 digital_ldo_top_VIA4 $T=375470 40260 0 0 $X=375220 $Y=40030
X8523 3 digital_ldo_top_VIA4 $T=375470 44340 0 0 $X=375220 $Y=44110
X8524 3 digital_ldo_top_VIA4 $T=375470 48420 0 0 $X=375220 $Y=48190
X8525 3 digital_ldo_top_VIA4 $T=375470 52500 0 0 $X=375220 $Y=52270
X8526 3 digital_ldo_top_VIA4 $T=375470 56580 0 0 $X=375220 $Y=56350
X8527 3 digital_ldo_top_VIA4 $T=375470 60660 0 0 $X=375220 $Y=60430
X8528 3 digital_ldo_top_VIA4 $T=375470 64740 0 0 $X=375220 $Y=64510
X8529 3 digital_ldo_top_VIA4 $T=375470 68820 0 0 $X=375220 $Y=68590
X8530 3 digital_ldo_top_VIA4 $T=375470 72900 0 0 $X=375220 $Y=72670
X8531 3 digital_ldo_top_VIA4 $T=375470 76980 0 0 $X=375220 $Y=76750
X8532 3 digital_ldo_top_VIA4 $T=375470 81060 0 0 $X=375220 $Y=80830
X8533 3 digital_ldo_top_VIA4 $T=375470 85140 0 0 $X=375220 $Y=84910
X8534 3 digital_ldo_top_VIA4 $T=375470 89220 0 0 $X=375220 $Y=88990
X8535 3 digital_ldo_top_VIA4 $T=375470 93300 0 0 $X=375220 $Y=93070
X8536 3 digital_ldo_top_VIA4 $T=375470 97380 0 0 $X=375220 $Y=97150
X8537 3 digital_ldo_top_VIA4 $T=375470 101460 0 0 $X=375220 $Y=101230
X8538 3 digital_ldo_top_VIA4 $T=375470 105540 0 0 $X=375220 $Y=105310
X8539 3 digital_ldo_top_VIA4 $T=375470 109620 0 0 $X=375220 $Y=109390
X8540 3 digital_ldo_top_VIA4 $T=375470 113700 0 0 $X=375220 $Y=113470
X8541 3 digital_ldo_top_VIA4 $T=375470 117780 0 0 $X=375220 $Y=117550
X8542 3 digital_ldo_top_VIA4 $T=375470 121860 0 0 $X=375220 $Y=121630
X8543 3 digital_ldo_top_VIA4 $T=375470 125940 0 0 $X=375220 $Y=125710
X8544 2 digital_ldo_top_VIA4 $T=376850 13060 0 0 $X=376600 $Y=12830
X8545 2 digital_ldo_top_VIA4 $T=376850 17140 0 0 $X=376600 $Y=16910
X8546 2 digital_ldo_top_VIA4 $T=376850 21220 0 0 $X=376600 $Y=20990
X8547 2 digital_ldo_top_VIA4 $T=376850 25300 0 0 $X=376600 $Y=25070
X8548 2 digital_ldo_top_VIA4 $T=376850 29380 0 0 $X=376600 $Y=29150
X8549 2 digital_ldo_top_VIA4 $T=376850 33460 0 0 $X=376600 $Y=33230
X8550 2 digital_ldo_top_VIA4 $T=376850 37540 0 0 $X=376600 $Y=37310
X8551 2 digital_ldo_top_VIA4 $T=376850 41620 0 0 $X=376600 $Y=41390
X8552 2 digital_ldo_top_VIA4 $T=376850 45700 0 0 $X=376600 $Y=45470
X8553 2 digital_ldo_top_VIA4 $T=376850 49780 0 0 $X=376600 $Y=49550
X8554 2 digital_ldo_top_VIA4 $T=376850 53860 0 0 $X=376600 $Y=53630
X8555 2 digital_ldo_top_VIA4 $T=376850 57940 0 0 $X=376600 $Y=57710
X8556 2 digital_ldo_top_VIA4 $T=376850 62020 0 0 $X=376600 $Y=61790
X8557 2 digital_ldo_top_VIA4 $T=376850 66100 0 0 $X=376600 $Y=65870
X8558 2 digital_ldo_top_VIA4 $T=376850 70180 0 0 $X=376600 $Y=69950
X8559 2 digital_ldo_top_VIA4 $T=376850 74260 0 0 $X=376600 $Y=74030
X8560 2 digital_ldo_top_VIA4 $T=376850 78340 0 0 $X=376600 $Y=78110
X8561 2 digital_ldo_top_VIA4 $T=376850 82420 0 0 $X=376600 $Y=82190
X8562 2 digital_ldo_top_VIA4 $T=376850 86500 0 0 $X=376600 $Y=86270
X8563 2 digital_ldo_top_VIA4 $T=376850 90580 0 0 $X=376600 $Y=90350
X8564 2 digital_ldo_top_VIA4 $T=376850 94660 0 0 $X=376600 $Y=94430
X8565 2 digital_ldo_top_VIA4 $T=376850 98740 0 0 $X=376600 $Y=98510
X8566 2 digital_ldo_top_VIA4 $T=376850 102820 0 0 $X=376600 $Y=102590
X8567 2 digital_ldo_top_VIA4 $T=376850 106900 0 0 $X=376600 $Y=106670
X8568 2 digital_ldo_top_VIA4 $T=376850 110980 0 0 $X=376600 $Y=110750
X8569 2 digital_ldo_top_VIA4 $T=376850 115060 0 0 $X=376600 $Y=114830
X8570 2 digital_ldo_top_VIA4 $T=376850 119140 0 0 $X=376600 $Y=118910
X8571 2 digital_ldo_top_VIA4 $T=376850 123220 0 0 $X=376600 $Y=122990
X8572 2 digital_ldo_top_VIA4 $T=376850 127300 0 0 $X=376600 $Y=127070
X8573 3 digital_ldo_top_VIA4 $T=379150 11700 0 0 $X=378900 $Y=11470
X8574 3 digital_ldo_top_VIA4 $T=379150 15780 0 0 $X=378900 $Y=15550
X8575 3 digital_ldo_top_VIA4 $T=379150 19860 0 0 $X=378900 $Y=19630
X8576 3 digital_ldo_top_VIA4 $T=379150 23940 0 0 $X=378900 $Y=23710
X8577 3 digital_ldo_top_VIA4 $T=379150 28020 0 0 $X=378900 $Y=27790
X8578 3 digital_ldo_top_VIA4 $T=379150 32100 0 0 $X=378900 $Y=31870
X8579 3 digital_ldo_top_VIA4 $T=379150 36180 0 0 $X=378900 $Y=35950
X8580 3 digital_ldo_top_VIA4 $T=379150 40260 0 0 $X=378900 $Y=40030
X8581 3 digital_ldo_top_VIA4 $T=379150 44340 0 0 $X=378900 $Y=44110
X8582 3 digital_ldo_top_VIA4 $T=379150 48420 0 0 $X=378900 $Y=48190
X8583 3 digital_ldo_top_VIA4 $T=379150 52500 0 0 $X=378900 $Y=52270
X8584 3 digital_ldo_top_VIA4 $T=379150 56580 0 0 $X=378900 $Y=56350
X8585 3 digital_ldo_top_VIA4 $T=379150 60660 0 0 $X=378900 $Y=60430
X8586 3 digital_ldo_top_VIA4 $T=379150 64740 0 0 $X=378900 $Y=64510
X8587 3 digital_ldo_top_VIA4 $T=379150 68820 0 0 $X=378900 $Y=68590
X8588 3 digital_ldo_top_VIA4 $T=379150 72900 0 0 $X=378900 $Y=72670
X8589 3 digital_ldo_top_VIA4 $T=379150 76980 0 0 $X=378900 $Y=76750
X8590 3 digital_ldo_top_VIA4 $T=379150 81060 0 0 $X=378900 $Y=80830
X8591 3 digital_ldo_top_VIA4 $T=379150 85140 0 0 $X=378900 $Y=84910
X8592 3 digital_ldo_top_VIA4 $T=379150 89220 0 0 $X=378900 $Y=88990
X8593 3 digital_ldo_top_VIA4 $T=379150 93300 0 0 $X=378900 $Y=93070
X8594 3 digital_ldo_top_VIA4 $T=379150 97380 0 0 $X=378900 $Y=97150
X8595 3 digital_ldo_top_VIA4 $T=379150 101460 0 0 $X=378900 $Y=101230
X8596 3 digital_ldo_top_VIA4 $T=379150 105540 0 0 $X=378900 $Y=105310
X8597 3 digital_ldo_top_VIA4 $T=379150 109620 0 0 $X=378900 $Y=109390
X8598 3 digital_ldo_top_VIA4 $T=379150 113700 0 0 $X=378900 $Y=113470
X8599 3 digital_ldo_top_VIA4 $T=379150 117780 0 0 $X=378900 $Y=117550
X8600 3 digital_ldo_top_VIA4 $T=379150 121860 0 0 $X=378900 $Y=121630
X8601 3 digital_ldo_top_VIA4 $T=379150 125940 0 0 $X=378900 $Y=125710
X8602 3 digital_ldo_top_VIA5 $T=103065 28020 0 0 $X=102900 $Y=27790
X8603 3 digital_ldo_top_VIA5 $T=103065 36180 0 0 $X=102900 $Y=35950
X8604 3 digital_ldo_top_VIA5 $T=103065 40260 0 0 $X=102900 $Y=40030
X8605 3 digital_ldo_top_VIA5 $T=103065 44340 0 0 $X=102900 $Y=44110
X8606 3 digital_ldo_top_VIA5 $T=103065 48420 0 0 $X=102900 $Y=48190
X8607 3 digital_ldo_top_VIA5 $T=103065 52500 0 0 $X=102900 $Y=52270
X8608 3 digital_ldo_top_VIA5 $T=103065 56580 0 0 $X=102900 $Y=56350
X8609 3 digital_ldo_top_VIA5 $T=103065 60660 0 0 $X=102900 $Y=60430
X8610 3 digital_ldo_top_VIA5 $T=103065 64740 0 0 $X=102900 $Y=64510
X8611 3 digital_ldo_top_VIA5 $T=103065 68820 0 0 $X=102900 $Y=68590
X8612 3 digital_ldo_top_VIA5 $T=103065 72900 0 0 $X=102900 $Y=72670
X8613 3 digital_ldo_top_VIA5 $T=103065 76980 0 0 $X=102900 $Y=76750
X8614 3 digital_ldo_top_VIA5 $T=103065 81060 0 0 $X=102900 $Y=80830
X8615 2 digital_ldo_top_VIA5 $T=307015 29380 0 0 $X=306850 $Y=29150
X8616 2 digital_ldo_top_VIA5 $T=307015 33460 0 0 $X=306850 $Y=33230
X8617 2 digital_ldo_top_VIA5 $T=307015 37540 0 0 $X=306850 $Y=37310
X8618 2 digital_ldo_top_VIA5 $T=307015 41620 0 0 $X=306850 $Y=41390
X8619 2 digital_ldo_top_VIA5 $T=307015 45700 0 0 $X=306850 $Y=45470
X8620 2 digital_ldo_top_VIA5 $T=307015 49780 0 0 $X=306850 $Y=49550
X8621 2 digital_ldo_top_VIA5 $T=307015 53860 0 0 $X=306850 $Y=53630
X8622 2 digital_ldo_top_VIA5 $T=307015 57940 0 0 $X=306850 $Y=57710
X8623 2 digital_ldo_top_VIA5 $T=307015 62020 0 0 $X=306850 $Y=61790
X8624 2 digital_ldo_top_VIA5 $T=307015 66100 0 0 $X=306850 $Y=65870
X8625 2 digital_ldo_top_VIA5 $T=307015 70180 0 0 $X=306850 $Y=69950
X8626 2 digital_ldo_top_VIA5 $T=307015 74260 0 0 $X=306850 $Y=74030
X8627 2 digital_ldo_top_VIA5 $T=307015 78340 0 0 $X=306850 $Y=78110
X8628 2 digital_ldo_top_VIA5 $T=307015 82420 0 0 $X=306850 $Y=82190
X8629 2 digital_ldo_top_VIA7 $T=20305 21220 0 0 $X=20020 $Y=20990
X8630 2 digital_ldo_top_VIA7 $T=20305 25300 0 0 $X=20020 $Y=25070
X8631 2 digital_ldo_top_VIA7 $T=80305 21220 0 0 $X=80020 $Y=20990
X8632 2 digital_ldo_top_VIA7 $T=80305 25300 0 0 $X=80020 $Y=25070
X8633 2 digital_ldo_top_VIA7 $T=80305 33460 0 0 $X=80020 $Y=33230
X8634 2 digital_ldo_top_VIA7 $T=80305 37540 0 0 $X=80020 $Y=37310
X8635 2 digital_ldo_top_VIA8 $T=325180 33460 0 0 $X=325000 $Y=33230
X8636 2 digital_ldo_top_VIA8 $T=325180 37540 0 0 $X=325000 $Y=37310
X8637 2 digital_ldo_top_VIA8 $T=325180 41620 0 0 $X=325000 $Y=41390
X8638 2 digital_ldo_top_VIA9 $T=60225 21220 0 0 $X=60000 $Y=20990
X8639 2 digital_ldo_top_VIA9 $T=60225 25300 0 0 $X=60000 $Y=25070
X8640 3 digital_ldo_top_VIA10 $T=12300 11700 0 0 $X=11830 $Y=11470
X8641 3 digital_ldo_top_VIA10 $T=12300 15780 0 0 $X=11830 $Y=15550
X8642 3 digital_ldo_top_VIA10 $T=12300 19860 0 0 $X=11830 $Y=19630
X8643 3 digital_ldo_top_VIA10 $T=12300 23940 0 0 $X=11830 $Y=23710
X8644 3 digital_ldo_top_VIA10 $T=12300 28020 0 0 $X=11830 $Y=27790
X8645 3 digital_ldo_top_VIA10 $T=12300 32100 0 0 $X=11830 $Y=31870
X8646 3 digital_ldo_top_VIA10 $T=12300 36180 0 0 $X=11830 $Y=35950
X8647 3 digital_ldo_top_VIA10 $T=12300 40260 0 0 $X=11830 $Y=40030
X8648 3 digital_ldo_top_VIA10 $T=12300 44340 0 0 $X=11830 $Y=44110
X8649 3 digital_ldo_top_VIA10 $T=12300 48420 0 0 $X=11830 $Y=48190
X8650 3 digital_ldo_top_VIA10 $T=12300 52500 0 0 $X=11830 $Y=52270
X8651 3 digital_ldo_top_VIA10 $T=12300 56580 0 0 $X=11830 $Y=56350
X8652 3 digital_ldo_top_VIA10 $T=12300 60660 0 0 $X=11830 $Y=60430
X8653 3 digital_ldo_top_VIA10 $T=12300 64740 0 0 $X=11830 $Y=64510
X8654 3 digital_ldo_top_VIA10 $T=12300 68820 0 0 $X=11830 $Y=68590
X8655 3 digital_ldo_top_VIA10 $T=12300 72900 0 0 $X=11830 $Y=72670
X8656 3 digital_ldo_top_VIA10 $T=12300 76980 0 0 $X=11830 $Y=76750
X8657 3 digital_ldo_top_VIA10 $T=12300 81060 0 0 $X=11830 $Y=80830
X8658 3 digital_ldo_top_VIA10 $T=12300 85140 0 0 $X=11830 $Y=84910
X8659 3 digital_ldo_top_VIA10 $T=12300 89220 0 0 $X=11830 $Y=88990
X8660 3 digital_ldo_top_VIA10 $T=12300 93300 0 0 $X=11830 $Y=93070
X8661 3 digital_ldo_top_VIA10 $T=12300 97380 0 0 $X=11830 $Y=97150
X8662 3 digital_ldo_top_VIA10 $T=12300 101460 0 0 $X=11830 $Y=101230
X8663 3 digital_ldo_top_VIA10 $T=12300 105540 0 0 $X=11830 $Y=105310
X8664 3 digital_ldo_top_VIA10 $T=12300 109620 0 0 $X=11830 $Y=109390
X8665 3 digital_ldo_top_VIA10 $T=12300 113700 0 0 $X=11830 $Y=113470
X8666 3 digital_ldo_top_VIA10 $T=12300 117780 0 0 $X=11830 $Y=117550
X8667 3 digital_ldo_top_VIA10 $T=12300 121860 0 0 $X=11830 $Y=121630
X8668 3 digital_ldo_top_VIA10 $T=12300 125940 0 0 $X=11830 $Y=125710
X8669 2 digital_ldo_top_VIA10 $T=14140 13060 0 0 $X=13670 $Y=12830
X8670 2 digital_ldo_top_VIA10 $T=14140 17140 0 0 $X=13670 $Y=16910
X8671 2 digital_ldo_top_VIA10 $T=14140 21220 0 0 $X=13670 $Y=20990
X8672 2 digital_ldo_top_VIA10 $T=14140 25300 0 0 $X=13670 $Y=25070
X8673 2 digital_ldo_top_VIA10 $T=14140 29380 0 0 $X=13670 $Y=29150
X8674 2 digital_ldo_top_VIA10 $T=14140 33460 0 0 $X=13670 $Y=33230
X8675 2 digital_ldo_top_VIA10 $T=14140 37540 0 0 $X=13670 $Y=37310
X8676 2 digital_ldo_top_VIA10 $T=14140 41620 0 0 $X=13670 $Y=41390
X8677 2 digital_ldo_top_VIA10 $T=14140 45700 0 0 $X=13670 $Y=45470
X8678 2 digital_ldo_top_VIA10 $T=14140 49780 0 0 $X=13670 $Y=49550
X8679 2 digital_ldo_top_VIA10 $T=14140 53860 0 0 $X=13670 $Y=53630
X8680 2 digital_ldo_top_VIA10 $T=14140 57940 0 0 $X=13670 $Y=57710
X8681 2 digital_ldo_top_VIA10 $T=14140 62020 0 0 $X=13670 $Y=61790
X8682 2 digital_ldo_top_VIA10 $T=14140 66100 0 0 $X=13670 $Y=65870
X8683 2 digital_ldo_top_VIA10 $T=14140 70180 0 0 $X=13670 $Y=69950
X8684 2 digital_ldo_top_VIA10 $T=14140 74260 0 0 $X=13670 $Y=74030
X8685 2 digital_ldo_top_VIA10 $T=14140 78340 0 0 $X=13670 $Y=78110
X8686 2 digital_ldo_top_VIA10 $T=14140 82420 0 0 $X=13670 $Y=82190
X8687 2 digital_ldo_top_VIA10 $T=14140 86500 0 0 $X=13670 $Y=86270
X8688 2 digital_ldo_top_VIA10 $T=14140 90580 0 0 $X=13670 $Y=90350
X8689 2 digital_ldo_top_VIA10 $T=14140 94660 0 0 $X=13670 $Y=94430
X8690 2 digital_ldo_top_VIA10 $T=14140 98740 0 0 $X=13670 $Y=98510
X8691 2 digital_ldo_top_VIA10 $T=14140 102820 0 0 $X=13670 $Y=102590
X8692 2 digital_ldo_top_VIA10 $T=14140 106900 0 0 $X=13670 $Y=106670
X8693 2 digital_ldo_top_VIA10 $T=14140 110980 0 0 $X=13670 $Y=110750
X8694 2 digital_ldo_top_VIA10 $T=14140 115060 0 0 $X=13670 $Y=114830
X8695 2 digital_ldo_top_VIA10 $T=14140 119140 0 0 $X=13670 $Y=118910
X8696 2 digital_ldo_top_VIA10 $T=14140 123220 0 0 $X=13670 $Y=122990
X8697 2 digital_ldo_top_VIA10 $T=14140 127300 0 0 $X=13670 $Y=127070
X8698 3 digital_ldo_top_VIA10 $T=17820 11700 0 0 $X=17350 $Y=11470
X8699 3 digital_ldo_top_VIA10 $T=17820 15780 0 0 $X=17350 $Y=15550
X8700 3 digital_ldo_top_VIA10 $T=17820 19860 0 0 $X=17350 $Y=19630
X8701 3 digital_ldo_top_VIA10 $T=17820 23940 0 0 $X=17350 $Y=23710
X8702 3 digital_ldo_top_VIA10 $T=17820 28020 0 0 $X=17350 $Y=27790
X8703 3 digital_ldo_top_VIA10 $T=17820 32100 0 0 $X=17350 $Y=31870
X8704 3 digital_ldo_top_VIA10 $T=17820 36180 0 0 $X=17350 $Y=35950
X8705 3 digital_ldo_top_VIA10 $T=17820 40260 0 0 $X=17350 $Y=40030
X8706 3 digital_ldo_top_VIA10 $T=17820 44340 0 0 $X=17350 $Y=44110
X8707 3 digital_ldo_top_VIA10 $T=17820 48420 0 0 $X=17350 $Y=48190
X8708 3 digital_ldo_top_VIA10 $T=17820 52500 0 0 $X=17350 $Y=52270
X8709 3 digital_ldo_top_VIA10 $T=17820 56580 0 0 $X=17350 $Y=56350
X8710 3 digital_ldo_top_VIA10 $T=17820 60660 0 0 $X=17350 $Y=60430
X8711 3 digital_ldo_top_VIA10 $T=17820 64740 0 0 $X=17350 $Y=64510
X8712 3 digital_ldo_top_VIA10 $T=17820 68820 0 0 $X=17350 $Y=68590
X8713 3 digital_ldo_top_VIA10 $T=17820 72900 0 0 $X=17350 $Y=72670
X8714 3 digital_ldo_top_VIA10 $T=17820 76980 0 0 $X=17350 $Y=76750
X8715 3 digital_ldo_top_VIA10 $T=17820 81060 0 0 $X=17350 $Y=80830
X8716 3 digital_ldo_top_VIA10 $T=17820 85140 0 0 $X=17350 $Y=84910
X8717 3 digital_ldo_top_VIA10 $T=17820 89220 0 0 $X=17350 $Y=88990
X8718 3 digital_ldo_top_VIA10 $T=17820 93300 0 0 $X=17350 $Y=93070
X8719 3 digital_ldo_top_VIA10 $T=17820 97380 0 0 $X=17350 $Y=97150
X8720 3 digital_ldo_top_VIA10 $T=17820 101460 0 0 $X=17350 $Y=101230
X8721 3 digital_ldo_top_VIA10 $T=17820 105540 0 0 $X=17350 $Y=105310
X8722 3 digital_ldo_top_VIA10 $T=17820 109620 0 0 $X=17350 $Y=109390
X8723 3 digital_ldo_top_VIA10 $T=17820 113700 0 0 $X=17350 $Y=113470
X8724 3 digital_ldo_top_VIA10 $T=17820 117780 0 0 $X=17350 $Y=117550
X8725 3 digital_ldo_top_VIA10 $T=17820 121860 0 0 $X=17350 $Y=121630
X8726 3 digital_ldo_top_VIA10 $T=17820 125940 0 0 $X=17350 $Y=125710
X8727 2 digital_ldo_top_VIA10 $T=19660 13060 0 0 $X=19190 $Y=12830
X8728 2 digital_ldo_top_VIA10 $T=19660 17140 0 0 $X=19190 $Y=16910
X8729 2 digital_ldo_top_VIA10 $T=19660 21220 0 0 $X=19190 $Y=20990
X8730 2 digital_ldo_top_VIA10 $T=19660 25300 0 0 $X=19190 $Y=25070
X8731 2 digital_ldo_top_VIA10 $T=19660 29380 0 0 $X=19190 $Y=29150
X8732 2 digital_ldo_top_VIA10 $T=19660 33460 0 0 $X=19190 $Y=33230
X8733 2 digital_ldo_top_VIA10 $T=19660 37540 0 0 $X=19190 $Y=37310
X8734 2 digital_ldo_top_VIA10 $T=19660 41620 0 0 $X=19190 $Y=41390
X8735 2 digital_ldo_top_VIA10 $T=19660 45700 0 0 $X=19190 $Y=45470
X8736 2 digital_ldo_top_VIA10 $T=19660 49780 0 0 $X=19190 $Y=49550
X8737 2 digital_ldo_top_VIA10 $T=19660 53860 0 0 $X=19190 $Y=53630
X8738 2 digital_ldo_top_VIA10 $T=19660 57940 0 0 $X=19190 $Y=57710
X8739 2 digital_ldo_top_VIA10 $T=19660 62020 0 0 $X=19190 $Y=61790
X8740 2 digital_ldo_top_VIA10 $T=19660 66100 0 0 $X=19190 $Y=65870
X8741 2 digital_ldo_top_VIA10 $T=19660 70180 0 0 $X=19190 $Y=69950
X8742 2 digital_ldo_top_VIA10 $T=19660 74260 0 0 $X=19190 $Y=74030
X8743 2 digital_ldo_top_VIA10 $T=19660 78340 0 0 $X=19190 $Y=78110
X8744 2 digital_ldo_top_VIA10 $T=19660 82420 0 0 $X=19190 $Y=82190
X8745 2 digital_ldo_top_VIA10 $T=19660 86500 0 0 $X=19190 $Y=86270
X8746 2 digital_ldo_top_VIA10 $T=19660 90580 0 0 $X=19190 $Y=90350
X8747 2 digital_ldo_top_VIA10 $T=19660 94660 0 0 $X=19190 $Y=94430
X8748 2 digital_ldo_top_VIA10 $T=19660 98740 0 0 $X=19190 $Y=98510
X8749 2 digital_ldo_top_VIA10 $T=19660 102820 0 0 $X=19190 $Y=102590
X8750 2 digital_ldo_top_VIA10 $T=19660 106900 0 0 $X=19190 $Y=106670
X8751 2 digital_ldo_top_VIA10 $T=19660 110980 0 0 $X=19190 $Y=110750
X8752 2 digital_ldo_top_VIA10 $T=19660 115060 0 0 $X=19190 $Y=114830
X8753 2 digital_ldo_top_VIA10 $T=19660 119140 0 0 $X=19190 $Y=118910
X8754 2 digital_ldo_top_VIA10 $T=19660 123220 0 0 $X=19190 $Y=122990
X8755 2 digital_ldo_top_VIA10 $T=19660 127300 0 0 $X=19190 $Y=127070
X8756 3 digital_ldo_top_VIA10 $T=23340 11700 0 0 $X=22870 $Y=11470
X8757 3 digital_ldo_top_VIA10 $T=23340 15780 0 0 $X=22870 $Y=15550
X8758 3 digital_ldo_top_VIA10 $T=23340 19860 0 0 $X=22870 $Y=19630
X8759 3 digital_ldo_top_VIA10 $T=23340 23940 0 0 $X=22870 $Y=23710
X8760 3 digital_ldo_top_VIA10 $T=23340 28020 0 0 $X=22870 $Y=27790
X8761 3 digital_ldo_top_VIA10 $T=23340 32100 0 0 $X=22870 $Y=31870
X8762 3 digital_ldo_top_VIA10 $T=23340 36180 0 0 $X=22870 $Y=35950
X8763 3 digital_ldo_top_VIA10 $T=23340 40260 0 0 $X=22870 $Y=40030
X8764 3 digital_ldo_top_VIA10 $T=23340 44340 0 0 $X=22870 $Y=44110
X8765 3 digital_ldo_top_VIA10 $T=23340 48420 0 0 $X=22870 $Y=48190
X8766 3 digital_ldo_top_VIA10 $T=23340 52500 0 0 $X=22870 $Y=52270
X8767 3 digital_ldo_top_VIA10 $T=23340 56580 0 0 $X=22870 $Y=56350
X8768 3 digital_ldo_top_VIA10 $T=23340 60660 0 0 $X=22870 $Y=60430
X8769 3 digital_ldo_top_VIA10 $T=23340 64740 0 0 $X=22870 $Y=64510
X8770 3 digital_ldo_top_VIA10 $T=23340 68820 0 0 $X=22870 $Y=68590
X8771 3 digital_ldo_top_VIA10 $T=23340 72900 0 0 $X=22870 $Y=72670
X8772 3 digital_ldo_top_VIA10 $T=23340 76980 0 0 $X=22870 $Y=76750
X8773 3 digital_ldo_top_VIA10 $T=23340 81060 0 0 $X=22870 $Y=80830
X8774 3 digital_ldo_top_VIA10 $T=23340 85140 0 0 $X=22870 $Y=84910
X8775 3 digital_ldo_top_VIA10 $T=23340 89220 0 0 $X=22870 $Y=88990
X8776 3 digital_ldo_top_VIA10 $T=23340 93300 0 0 $X=22870 $Y=93070
X8777 3 digital_ldo_top_VIA10 $T=23340 97380 0 0 $X=22870 $Y=97150
X8778 3 digital_ldo_top_VIA10 $T=23340 101460 0 0 $X=22870 $Y=101230
X8779 3 digital_ldo_top_VIA10 $T=23340 105540 0 0 $X=22870 $Y=105310
X8780 3 digital_ldo_top_VIA10 $T=23340 109620 0 0 $X=22870 $Y=109390
X8781 3 digital_ldo_top_VIA10 $T=23340 113700 0 0 $X=22870 $Y=113470
X8782 3 digital_ldo_top_VIA10 $T=23340 117780 0 0 $X=22870 $Y=117550
X8783 3 digital_ldo_top_VIA10 $T=23340 121860 0 0 $X=22870 $Y=121630
X8784 3 digital_ldo_top_VIA10 $T=23340 125940 0 0 $X=22870 $Y=125710
X8785 2 digital_ldo_top_VIA10 $T=25180 13060 0 0 $X=24710 $Y=12830
X8786 2 digital_ldo_top_VIA10 $T=25180 17140 0 0 $X=24710 $Y=16910
X8787 2 digital_ldo_top_VIA10 $T=25180 21220 0 0 $X=24710 $Y=20990
X8788 2 digital_ldo_top_VIA10 $T=25180 25300 0 0 $X=24710 $Y=25070
X8789 2 digital_ldo_top_VIA10 $T=25180 29380 0 0 $X=24710 $Y=29150
X8790 2 digital_ldo_top_VIA10 $T=25180 33460 0 0 $X=24710 $Y=33230
X8791 2 digital_ldo_top_VIA10 $T=25180 37540 0 0 $X=24710 $Y=37310
X8792 2 digital_ldo_top_VIA10 $T=25180 41620 0 0 $X=24710 $Y=41390
X8793 2 digital_ldo_top_VIA10 $T=25180 45700 0 0 $X=24710 $Y=45470
X8794 2 digital_ldo_top_VIA10 $T=25180 49780 0 0 $X=24710 $Y=49550
X8795 2 digital_ldo_top_VIA10 $T=25180 53860 0 0 $X=24710 $Y=53630
X8796 2 digital_ldo_top_VIA10 $T=25180 57940 0 0 $X=24710 $Y=57710
X8797 2 digital_ldo_top_VIA10 $T=25180 62020 0 0 $X=24710 $Y=61790
X8798 2 digital_ldo_top_VIA10 $T=25180 66100 0 0 $X=24710 $Y=65870
X8799 2 digital_ldo_top_VIA10 $T=25180 70180 0 0 $X=24710 $Y=69950
X8800 2 digital_ldo_top_VIA10 $T=25180 74260 0 0 $X=24710 $Y=74030
X8801 2 digital_ldo_top_VIA10 $T=25180 78340 0 0 $X=24710 $Y=78110
X8802 2 digital_ldo_top_VIA10 $T=25180 82420 0 0 $X=24710 $Y=82190
X8803 2 digital_ldo_top_VIA10 $T=25180 86500 0 0 $X=24710 $Y=86270
X8804 2 digital_ldo_top_VIA10 $T=25180 90580 0 0 $X=24710 $Y=90350
X8805 2 digital_ldo_top_VIA10 $T=25180 94660 0 0 $X=24710 $Y=94430
X8806 2 digital_ldo_top_VIA10 $T=25180 98740 0 0 $X=24710 $Y=98510
X8807 2 digital_ldo_top_VIA10 $T=25180 102820 0 0 $X=24710 $Y=102590
X8808 2 digital_ldo_top_VIA10 $T=25180 106900 0 0 $X=24710 $Y=106670
X8809 2 digital_ldo_top_VIA10 $T=25180 110980 0 0 $X=24710 $Y=110750
X8810 2 digital_ldo_top_VIA10 $T=25180 115060 0 0 $X=24710 $Y=114830
X8811 2 digital_ldo_top_VIA10 $T=25180 119140 0 0 $X=24710 $Y=118910
X8812 2 digital_ldo_top_VIA10 $T=25180 123220 0 0 $X=24710 $Y=122990
X8813 2 digital_ldo_top_VIA10 $T=25180 127300 0 0 $X=24710 $Y=127070
X8814 3 digital_ldo_top_VIA10 $T=28860 11700 0 0 $X=28390 $Y=11470
X8815 3 digital_ldo_top_VIA10 $T=28860 15780 0 0 $X=28390 $Y=15550
X8816 3 digital_ldo_top_VIA10 $T=28860 19860 0 0 $X=28390 $Y=19630
X8817 3 digital_ldo_top_VIA10 $T=28860 23940 0 0 $X=28390 $Y=23710
X8818 3 digital_ldo_top_VIA10 $T=28860 28020 0 0 $X=28390 $Y=27790
X8819 3 digital_ldo_top_VIA10 $T=28860 32100 0 0 $X=28390 $Y=31870
X8820 3 digital_ldo_top_VIA10 $T=28860 36180 0 0 $X=28390 $Y=35950
X8821 3 digital_ldo_top_VIA10 $T=28860 40260 0 0 $X=28390 $Y=40030
X8822 3 digital_ldo_top_VIA10 $T=28860 44340 0 0 $X=28390 $Y=44110
X8823 3 digital_ldo_top_VIA10 $T=28860 48420 0 0 $X=28390 $Y=48190
X8824 3 digital_ldo_top_VIA10 $T=28860 52500 0 0 $X=28390 $Y=52270
X8825 3 digital_ldo_top_VIA10 $T=28860 56580 0 0 $X=28390 $Y=56350
X8826 3 digital_ldo_top_VIA10 $T=28860 60660 0 0 $X=28390 $Y=60430
X8827 3 digital_ldo_top_VIA10 $T=28860 64740 0 0 $X=28390 $Y=64510
X8828 3 digital_ldo_top_VIA10 $T=28860 68820 0 0 $X=28390 $Y=68590
X8829 3 digital_ldo_top_VIA10 $T=28860 72900 0 0 $X=28390 $Y=72670
X8830 3 digital_ldo_top_VIA10 $T=28860 76980 0 0 $X=28390 $Y=76750
X8831 3 digital_ldo_top_VIA10 $T=28860 81060 0 0 $X=28390 $Y=80830
X8832 3 digital_ldo_top_VIA10 $T=28860 85140 0 0 $X=28390 $Y=84910
X8833 3 digital_ldo_top_VIA10 $T=28860 89220 0 0 $X=28390 $Y=88990
X8834 3 digital_ldo_top_VIA10 $T=28860 93300 0 0 $X=28390 $Y=93070
X8835 3 digital_ldo_top_VIA10 $T=28860 97380 0 0 $X=28390 $Y=97150
X8836 3 digital_ldo_top_VIA10 $T=28860 101460 0 0 $X=28390 $Y=101230
X8837 3 digital_ldo_top_VIA10 $T=28860 105540 0 0 $X=28390 $Y=105310
X8838 3 digital_ldo_top_VIA10 $T=28860 109620 0 0 $X=28390 $Y=109390
X8839 3 digital_ldo_top_VIA10 $T=28860 113700 0 0 $X=28390 $Y=113470
X8840 3 digital_ldo_top_VIA10 $T=28860 117780 0 0 $X=28390 $Y=117550
X8841 3 digital_ldo_top_VIA10 $T=28860 121860 0 0 $X=28390 $Y=121630
X8842 3 digital_ldo_top_VIA10 $T=28860 125940 0 0 $X=28390 $Y=125710
X8843 2 digital_ldo_top_VIA10 $T=30700 13060 0 0 $X=30230 $Y=12830
X8844 2 digital_ldo_top_VIA10 $T=30700 17140 0 0 $X=30230 $Y=16910
X8845 2 digital_ldo_top_VIA10 $T=30700 21220 0 0 $X=30230 $Y=20990
X8846 2 digital_ldo_top_VIA10 $T=30700 25300 0 0 $X=30230 $Y=25070
X8847 2 digital_ldo_top_VIA10 $T=30700 29380 0 0 $X=30230 $Y=29150
X8848 2 digital_ldo_top_VIA10 $T=30700 33460 0 0 $X=30230 $Y=33230
X8849 2 digital_ldo_top_VIA10 $T=30700 37540 0 0 $X=30230 $Y=37310
X8850 2 digital_ldo_top_VIA10 $T=30700 41620 0 0 $X=30230 $Y=41390
X8851 2 digital_ldo_top_VIA10 $T=30700 45700 0 0 $X=30230 $Y=45470
X8852 2 digital_ldo_top_VIA10 $T=30700 49780 0 0 $X=30230 $Y=49550
X8853 2 digital_ldo_top_VIA10 $T=30700 53860 0 0 $X=30230 $Y=53630
X8854 2 digital_ldo_top_VIA10 $T=30700 57940 0 0 $X=30230 $Y=57710
X8855 2 digital_ldo_top_VIA10 $T=30700 62020 0 0 $X=30230 $Y=61790
X8856 2 digital_ldo_top_VIA10 $T=30700 66100 0 0 $X=30230 $Y=65870
X8857 2 digital_ldo_top_VIA10 $T=30700 70180 0 0 $X=30230 $Y=69950
X8858 2 digital_ldo_top_VIA10 $T=30700 74260 0 0 $X=30230 $Y=74030
X8859 2 digital_ldo_top_VIA10 $T=30700 78340 0 0 $X=30230 $Y=78110
X8860 2 digital_ldo_top_VIA10 $T=30700 82420 0 0 $X=30230 $Y=82190
X8861 2 digital_ldo_top_VIA10 $T=30700 86500 0 0 $X=30230 $Y=86270
X8862 2 digital_ldo_top_VIA10 $T=30700 90580 0 0 $X=30230 $Y=90350
X8863 2 digital_ldo_top_VIA10 $T=30700 94660 0 0 $X=30230 $Y=94430
X8864 2 digital_ldo_top_VIA10 $T=30700 98740 0 0 $X=30230 $Y=98510
X8865 2 digital_ldo_top_VIA10 $T=30700 102820 0 0 $X=30230 $Y=102590
X8866 2 digital_ldo_top_VIA10 $T=30700 106900 0 0 $X=30230 $Y=106670
X8867 2 digital_ldo_top_VIA10 $T=30700 110980 0 0 $X=30230 $Y=110750
X8868 2 digital_ldo_top_VIA10 $T=30700 115060 0 0 $X=30230 $Y=114830
X8869 2 digital_ldo_top_VIA10 $T=30700 119140 0 0 $X=30230 $Y=118910
X8870 2 digital_ldo_top_VIA10 $T=30700 123220 0 0 $X=30230 $Y=122990
X8871 2 digital_ldo_top_VIA10 $T=30700 127300 0 0 $X=30230 $Y=127070
X8872 3 digital_ldo_top_VIA10 $T=34380 11700 0 0 $X=33910 $Y=11470
X8873 3 digital_ldo_top_VIA10 $T=34380 15780 0 0 $X=33910 $Y=15550
X8874 3 digital_ldo_top_VIA10 $T=34380 19860 0 0 $X=33910 $Y=19630
X8875 3 digital_ldo_top_VIA10 $T=34380 23940 0 0 $X=33910 $Y=23710
X8876 3 digital_ldo_top_VIA10 $T=34380 28020 0 0 $X=33910 $Y=27790
X8877 3 digital_ldo_top_VIA10 $T=34380 32100 0 0 $X=33910 $Y=31870
X8878 3 digital_ldo_top_VIA10 $T=34380 36180 0 0 $X=33910 $Y=35950
X8879 3 digital_ldo_top_VIA10 $T=34380 40260 0 0 $X=33910 $Y=40030
X8880 3 digital_ldo_top_VIA10 $T=34380 44340 0 0 $X=33910 $Y=44110
X8881 3 digital_ldo_top_VIA10 $T=34380 48420 0 0 $X=33910 $Y=48190
X8882 3 digital_ldo_top_VIA10 $T=34380 52500 0 0 $X=33910 $Y=52270
X8883 3 digital_ldo_top_VIA10 $T=34380 56580 0 0 $X=33910 $Y=56350
X8884 3 digital_ldo_top_VIA10 $T=34380 60660 0 0 $X=33910 $Y=60430
X8885 3 digital_ldo_top_VIA10 $T=34380 64740 0 0 $X=33910 $Y=64510
X8886 3 digital_ldo_top_VIA10 $T=34380 68820 0 0 $X=33910 $Y=68590
X8887 3 digital_ldo_top_VIA10 $T=34380 72900 0 0 $X=33910 $Y=72670
X8888 3 digital_ldo_top_VIA10 $T=34380 76980 0 0 $X=33910 $Y=76750
X8889 3 digital_ldo_top_VIA10 $T=34380 81060 0 0 $X=33910 $Y=80830
X8890 3 digital_ldo_top_VIA10 $T=34380 85140 0 0 $X=33910 $Y=84910
X8891 3 digital_ldo_top_VIA10 $T=34380 89220 0 0 $X=33910 $Y=88990
X8892 3 digital_ldo_top_VIA10 $T=34380 93300 0 0 $X=33910 $Y=93070
X8893 3 digital_ldo_top_VIA10 $T=34380 97380 0 0 $X=33910 $Y=97150
X8894 3 digital_ldo_top_VIA10 $T=34380 101460 0 0 $X=33910 $Y=101230
X8895 3 digital_ldo_top_VIA10 $T=34380 105540 0 0 $X=33910 $Y=105310
X8896 3 digital_ldo_top_VIA10 $T=34380 109620 0 0 $X=33910 $Y=109390
X8897 3 digital_ldo_top_VIA10 $T=34380 113700 0 0 $X=33910 $Y=113470
X8898 3 digital_ldo_top_VIA10 $T=34380 117780 0 0 $X=33910 $Y=117550
X8899 3 digital_ldo_top_VIA10 $T=34380 121860 0 0 $X=33910 $Y=121630
X8900 3 digital_ldo_top_VIA10 $T=34380 125940 0 0 $X=33910 $Y=125710
X8901 2 digital_ldo_top_VIA10 $T=36220 13060 0 0 $X=35750 $Y=12830
X8902 2 digital_ldo_top_VIA10 $T=36220 17140 0 0 $X=35750 $Y=16910
X8903 2 digital_ldo_top_VIA10 $T=36220 21220 0 0 $X=35750 $Y=20990
X8904 2 digital_ldo_top_VIA10 $T=36220 25300 0 0 $X=35750 $Y=25070
X8905 2 digital_ldo_top_VIA10 $T=36220 29380 0 0 $X=35750 $Y=29150
X8906 2 digital_ldo_top_VIA10 $T=36220 33460 0 0 $X=35750 $Y=33230
X8907 2 digital_ldo_top_VIA10 $T=36220 37540 0 0 $X=35750 $Y=37310
X8908 2 digital_ldo_top_VIA10 $T=36220 41620 0 0 $X=35750 $Y=41390
X8909 2 digital_ldo_top_VIA10 $T=36220 45700 0 0 $X=35750 $Y=45470
X8910 2 digital_ldo_top_VIA10 $T=36220 49780 0 0 $X=35750 $Y=49550
X8911 2 digital_ldo_top_VIA10 $T=36220 53860 0 0 $X=35750 $Y=53630
X8912 2 digital_ldo_top_VIA10 $T=36220 57940 0 0 $X=35750 $Y=57710
X8913 2 digital_ldo_top_VIA10 $T=36220 62020 0 0 $X=35750 $Y=61790
X8914 2 digital_ldo_top_VIA10 $T=36220 66100 0 0 $X=35750 $Y=65870
X8915 2 digital_ldo_top_VIA10 $T=36220 70180 0 0 $X=35750 $Y=69950
X8916 2 digital_ldo_top_VIA10 $T=36220 74260 0 0 $X=35750 $Y=74030
X8917 2 digital_ldo_top_VIA10 $T=36220 78340 0 0 $X=35750 $Y=78110
X8918 2 digital_ldo_top_VIA10 $T=36220 82420 0 0 $X=35750 $Y=82190
X8919 2 digital_ldo_top_VIA10 $T=36220 86500 0 0 $X=35750 $Y=86270
X8920 2 digital_ldo_top_VIA10 $T=36220 90580 0 0 $X=35750 $Y=90350
X8921 2 digital_ldo_top_VIA10 $T=36220 94660 0 0 $X=35750 $Y=94430
X8922 2 digital_ldo_top_VIA10 $T=36220 98740 0 0 $X=35750 $Y=98510
X8923 2 digital_ldo_top_VIA10 $T=36220 102820 0 0 $X=35750 $Y=102590
X8924 2 digital_ldo_top_VIA10 $T=36220 106900 0 0 $X=35750 $Y=106670
X8925 2 digital_ldo_top_VIA10 $T=36220 110980 0 0 $X=35750 $Y=110750
X8926 2 digital_ldo_top_VIA10 $T=36220 115060 0 0 $X=35750 $Y=114830
X8927 2 digital_ldo_top_VIA10 $T=36220 119140 0 0 $X=35750 $Y=118910
X8928 2 digital_ldo_top_VIA10 $T=36220 123220 0 0 $X=35750 $Y=122990
X8929 2 digital_ldo_top_VIA10 $T=36220 127300 0 0 $X=35750 $Y=127070
X8930 3 digital_ldo_top_VIA10 $T=39900 11700 0 0 $X=39430 $Y=11470
X8931 3 digital_ldo_top_VIA10 $T=39900 15780 0 0 $X=39430 $Y=15550
X8932 3 digital_ldo_top_VIA10 $T=39900 19860 0 0 $X=39430 $Y=19630
X8933 3 digital_ldo_top_VIA10 $T=39900 23940 0 0 $X=39430 $Y=23710
X8934 3 digital_ldo_top_VIA10 $T=39900 28020 0 0 $X=39430 $Y=27790
X8935 3 digital_ldo_top_VIA10 $T=39900 32100 0 0 $X=39430 $Y=31870
X8936 3 digital_ldo_top_VIA10 $T=39900 36180 0 0 $X=39430 $Y=35950
X8937 3 digital_ldo_top_VIA10 $T=39900 40260 0 0 $X=39430 $Y=40030
X8938 3 digital_ldo_top_VIA10 $T=39900 44340 0 0 $X=39430 $Y=44110
X8939 3 digital_ldo_top_VIA10 $T=39900 48420 0 0 $X=39430 $Y=48190
X8940 3 digital_ldo_top_VIA10 $T=39900 52500 0 0 $X=39430 $Y=52270
X8941 3 digital_ldo_top_VIA10 $T=39900 56580 0 0 $X=39430 $Y=56350
X8942 3 digital_ldo_top_VIA10 $T=39900 60660 0 0 $X=39430 $Y=60430
X8943 3 digital_ldo_top_VIA10 $T=39900 64740 0 0 $X=39430 $Y=64510
X8944 3 digital_ldo_top_VIA10 $T=39900 68820 0 0 $X=39430 $Y=68590
X8945 3 digital_ldo_top_VIA10 $T=39900 72900 0 0 $X=39430 $Y=72670
X8946 3 digital_ldo_top_VIA10 $T=39900 76980 0 0 $X=39430 $Y=76750
X8947 3 digital_ldo_top_VIA10 $T=39900 81060 0 0 $X=39430 $Y=80830
X8948 3 digital_ldo_top_VIA10 $T=39900 85140 0 0 $X=39430 $Y=84910
X8949 3 digital_ldo_top_VIA10 $T=39900 89220 0 0 $X=39430 $Y=88990
X8950 3 digital_ldo_top_VIA10 $T=39900 93300 0 0 $X=39430 $Y=93070
X8951 3 digital_ldo_top_VIA10 $T=39900 97380 0 0 $X=39430 $Y=97150
X8952 3 digital_ldo_top_VIA10 $T=39900 101460 0 0 $X=39430 $Y=101230
X8953 3 digital_ldo_top_VIA10 $T=39900 105540 0 0 $X=39430 $Y=105310
X8954 3 digital_ldo_top_VIA10 $T=39900 109620 0 0 $X=39430 $Y=109390
X8955 3 digital_ldo_top_VIA10 $T=39900 113700 0 0 $X=39430 $Y=113470
X8956 3 digital_ldo_top_VIA10 $T=39900 117780 0 0 $X=39430 $Y=117550
X8957 3 digital_ldo_top_VIA10 $T=39900 121860 0 0 $X=39430 $Y=121630
X8958 3 digital_ldo_top_VIA10 $T=39900 125940 0 0 $X=39430 $Y=125710
X8959 2 digital_ldo_top_VIA10 $T=41740 13060 0 0 $X=41270 $Y=12830
X8960 2 digital_ldo_top_VIA10 $T=41740 17140 0 0 $X=41270 $Y=16910
X8961 2 digital_ldo_top_VIA10 $T=41740 21220 0 0 $X=41270 $Y=20990
X8962 2 digital_ldo_top_VIA10 $T=41740 25300 0 0 $X=41270 $Y=25070
X8963 2 digital_ldo_top_VIA10 $T=41740 29380 0 0 $X=41270 $Y=29150
X8964 2 digital_ldo_top_VIA10 $T=41740 33460 0 0 $X=41270 $Y=33230
X8965 2 digital_ldo_top_VIA10 $T=41740 37540 0 0 $X=41270 $Y=37310
X8966 2 digital_ldo_top_VIA10 $T=41740 41620 0 0 $X=41270 $Y=41390
X8967 2 digital_ldo_top_VIA10 $T=41740 45700 0 0 $X=41270 $Y=45470
X8968 2 digital_ldo_top_VIA10 $T=41740 49780 0 0 $X=41270 $Y=49550
X8969 2 digital_ldo_top_VIA10 $T=41740 53860 0 0 $X=41270 $Y=53630
X8970 2 digital_ldo_top_VIA10 $T=41740 57940 0 0 $X=41270 $Y=57710
X8971 2 digital_ldo_top_VIA10 $T=41740 62020 0 0 $X=41270 $Y=61790
X8972 2 digital_ldo_top_VIA10 $T=41740 66100 0 0 $X=41270 $Y=65870
X8973 2 digital_ldo_top_VIA10 $T=41740 70180 0 0 $X=41270 $Y=69950
X8974 2 digital_ldo_top_VIA10 $T=41740 74260 0 0 $X=41270 $Y=74030
X8975 2 digital_ldo_top_VIA10 $T=41740 78340 0 0 $X=41270 $Y=78110
X8976 2 digital_ldo_top_VIA10 $T=41740 82420 0 0 $X=41270 $Y=82190
X8977 2 digital_ldo_top_VIA10 $T=41740 86500 0 0 $X=41270 $Y=86270
X8978 2 digital_ldo_top_VIA10 $T=41740 90580 0 0 $X=41270 $Y=90350
X8979 2 digital_ldo_top_VIA10 $T=41740 94660 0 0 $X=41270 $Y=94430
X8980 2 digital_ldo_top_VIA10 $T=41740 98740 0 0 $X=41270 $Y=98510
X8981 2 digital_ldo_top_VIA10 $T=41740 102820 0 0 $X=41270 $Y=102590
X8982 2 digital_ldo_top_VIA10 $T=41740 106900 0 0 $X=41270 $Y=106670
X8983 2 digital_ldo_top_VIA10 $T=41740 110980 0 0 $X=41270 $Y=110750
X8984 2 digital_ldo_top_VIA10 $T=41740 115060 0 0 $X=41270 $Y=114830
X8985 2 digital_ldo_top_VIA10 $T=41740 119140 0 0 $X=41270 $Y=118910
X8986 2 digital_ldo_top_VIA10 $T=41740 123220 0 0 $X=41270 $Y=122990
X8987 2 digital_ldo_top_VIA10 $T=41740 127300 0 0 $X=41270 $Y=127070
X8988 3 digital_ldo_top_VIA10 $T=45420 11700 0 0 $X=44950 $Y=11470
X8989 3 digital_ldo_top_VIA10 $T=45420 15780 0 0 $X=44950 $Y=15550
X8990 3 digital_ldo_top_VIA10 $T=45420 19860 0 0 $X=44950 $Y=19630
X8991 3 digital_ldo_top_VIA10 $T=45420 23940 0 0 $X=44950 $Y=23710
X8992 3 digital_ldo_top_VIA10 $T=45420 28020 0 0 $X=44950 $Y=27790
X8993 3 digital_ldo_top_VIA10 $T=45420 32100 0 0 $X=44950 $Y=31870
X8994 3 digital_ldo_top_VIA10 $T=45420 36180 0 0 $X=44950 $Y=35950
X8995 3 digital_ldo_top_VIA10 $T=45420 40260 0 0 $X=44950 $Y=40030
X8996 3 digital_ldo_top_VIA10 $T=45420 44340 0 0 $X=44950 $Y=44110
X8997 3 digital_ldo_top_VIA10 $T=45420 48420 0 0 $X=44950 $Y=48190
X8998 3 digital_ldo_top_VIA10 $T=45420 52500 0 0 $X=44950 $Y=52270
X8999 3 digital_ldo_top_VIA10 $T=45420 56580 0 0 $X=44950 $Y=56350
X9000 3 digital_ldo_top_VIA10 $T=45420 60660 0 0 $X=44950 $Y=60430
X9001 3 digital_ldo_top_VIA10 $T=45420 64740 0 0 $X=44950 $Y=64510
X9002 3 digital_ldo_top_VIA10 $T=45420 68820 0 0 $X=44950 $Y=68590
X9003 3 digital_ldo_top_VIA10 $T=45420 72900 0 0 $X=44950 $Y=72670
X9004 3 digital_ldo_top_VIA10 $T=45420 76980 0 0 $X=44950 $Y=76750
X9005 3 digital_ldo_top_VIA10 $T=45420 81060 0 0 $X=44950 $Y=80830
X9006 3 digital_ldo_top_VIA10 $T=45420 85140 0 0 $X=44950 $Y=84910
X9007 3 digital_ldo_top_VIA10 $T=45420 89220 0 0 $X=44950 $Y=88990
X9008 3 digital_ldo_top_VIA10 $T=45420 93300 0 0 $X=44950 $Y=93070
X9009 3 digital_ldo_top_VIA10 $T=45420 97380 0 0 $X=44950 $Y=97150
X9010 3 digital_ldo_top_VIA10 $T=45420 101460 0 0 $X=44950 $Y=101230
X9011 3 digital_ldo_top_VIA10 $T=45420 105540 0 0 $X=44950 $Y=105310
X9012 3 digital_ldo_top_VIA10 $T=45420 109620 0 0 $X=44950 $Y=109390
X9013 3 digital_ldo_top_VIA10 $T=45420 113700 0 0 $X=44950 $Y=113470
X9014 3 digital_ldo_top_VIA10 $T=45420 117780 0 0 $X=44950 $Y=117550
X9015 3 digital_ldo_top_VIA10 $T=45420 121860 0 0 $X=44950 $Y=121630
X9016 3 digital_ldo_top_VIA10 $T=45420 125940 0 0 $X=44950 $Y=125710
X9017 2 digital_ldo_top_VIA10 $T=47260 13060 0 0 $X=46790 $Y=12830
X9018 2 digital_ldo_top_VIA10 $T=47260 17140 0 0 $X=46790 $Y=16910
X9019 2 digital_ldo_top_VIA10 $T=47260 21220 0 0 $X=46790 $Y=20990
X9020 2 digital_ldo_top_VIA10 $T=47260 25300 0 0 $X=46790 $Y=25070
X9021 2 digital_ldo_top_VIA10 $T=47260 29380 0 0 $X=46790 $Y=29150
X9022 2 digital_ldo_top_VIA10 $T=47260 33460 0 0 $X=46790 $Y=33230
X9023 2 digital_ldo_top_VIA10 $T=47260 37540 0 0 $X=46790 $Y=37310
X9024 2 digital_ldo_top_VIA10 $T=47260 41620 0 0 $X=46790 $Y=41390
X9025 2 digital_ldo_top_VIA10 $T=47260 45700 0 0 $X=46790 $Y=45470
X9026 2 digital_ldo_top_VIA10 $T=47260 49780 0 0 $X=46790 $Y=49550
X9027 2 digital_ldo_top_VIA10 $T=47260 53860 0 0 $X=46790 $Y=53630
X9028 2 digital_ldo_top_VIA10 $T=47260 57940 0 0 $X=46790 $Y=57710
X9029 2 digital_ldo_top_VIA10 $T=47260 62020 0 0 $X=46790 $Y=61790
X9030 2 digital_ldo_top_VIA10 $T=47260 66100 0 0 $X=46790 $Y=65870
X9031 2 digital_ldo_top_VIA10 $T=47260 70180 0 0 $X=46790 $Y=69950
X9032 2 digital_ldo_top_VIA10 $T=47260 74260 0 0 $X=46790 $Y=74030
X9033 2 digital_ldo_top_VIA10 $T=47260 78340 0 0 $X=46790 $Y=78110
X9034 2 digital_ldo_top_VIA10 $T=47260 82420 0 0 $X=46790 $Y=82190
X9035 2 digital_ldo_top_VIA10 $T=47260 86500 0 0 $X=46790 $Y=86270
X9036 2 digital_ldo_top_VIA10 $T=47260 90580 0 0 $X=46790 $Y=90350
X9037 2 digital_ldo_top_VIA10 $T=47260 94660 0 0 $X=46790 $Y=94430
X9038 2 digital_ldo_top_VIA10 $T=47260 98740 0 0 $X=46790 $Y=98510
X9039 2 digital_ldo_top_VIA10 $T=47260 102820 0 0 $X=46790 $Y=102590
X9040 2 digital_ldo_top_VIA10 $T=47260 106900 0 0 $X=46790 $Y=106670
X9041 2 digital_ldo_top_VIA10 $T=47260 110980 0 0 $X=46790 $Y=110750
X9042 2 digital_ldo_top_VIA10 $T=47260 115060 0 0 $X=46790 $Y=114830
X9043 2 digital_ldo_top_VIA10 $T=47260 119140 0 0 $X=46790 $Y=118910
X9044 2 digital_ldo_top_VIA10 $T=47260 123220 0 0 $X=46790 $Y=122990
X9045 2 digital_ldo_top_VIA10 $T=47260 127300 0 0 $X=46790 $Y=127070
X9046 3 digital_ldo_top_VIA10 $T=50940 11700 0 0 $X=50470 $Y=11470
X9047 3 digital_ldo_top_VIA10 $T=50940 15780 0 0 $X=50470 $Y=15550
X9048 3 digital_ldo_top_VIA10 $T=50940 19860 0 0 $X=50470 $Y=19630
X9049 3 digital_ldo_top_VIA10 $T=50940 23940 0 0 $X=50470 $Y=23710
X9050 3 digital_ldo_top_VIA10 $T=50940 28020 0 0 $X=50470 $Y=27790
X9051 3 digital_ldo_top_VIA10 $T=50940 32100 0 0 $X=50470 $Y=31870
X9052 3 digital_ldo_top_VIA10 $T=50940 36180 0 0 $X=50470 $Y=35950
X9053 3 digital_ldo_top_VIA10 $T=50940 40260 0 0 $X=50470 $Y=40030
X9054 3 digital_ldo_top_VIA10 $T=50940 44340 0 0 $X=50470 $Y=44110
X9055 3 digital_ldo_top_VIA10 $T=50940 48420 0 0 $X=50470 $Y=48190
X9056 3 digital_ldo_top_VIA10 $T=50940 52500 0 0 $X=50470 $Y=52270
X9057 3 digital_ldo_top_VIA10 $T=50940 56580 0 0 $X=50470 $Y=56350
X9058 3 digital_ldo_top_VIA10 $T=50940 60660 0 0 $X=50470 $Y=60430
X9059 3 digital_ldo_top_VIA10 $T=50940 64740 0 0 $X=50470 $Y=64510
X9060 3 digital_ldo_top_VIA10 $T=50940 68820 0 0 $X=50470 $Y=68590
X9061 3 digital_ldo_top_VIA10 $T=50940 72900 0 0 $X=50470 $Y=72670
X9062 3 digital_ldo_top_VIA10 $T=50940 76980 0 0 $X=50470 $Y=76750
X9063 3 digital_ldo_top_VIA10 $T=50940 81060 0 0 $X=50470 $Y=80830
X9064 3 digital_ldo_top_VIA10 $T=50940 85140 0 0 $X=50470 $Y=84910
X9065 3 digital_ldo_top_VIA10 $T=50940 89220 0 0 $X=50470 $Y=88990
X9066 3 digital_ldo_top_VIA10 $T=50940 93300 0 0 $X=50470 $Y=93070
X9067 3 digital_ldo_top_VIA10 $T=50940 97380 0 0 $X=50470 $Y=97150
X9068 3 digital_ldo_top_VIA10 $T=50940 101460 0 0 $X=50470 $Y=101230
X9069 3 digital_ldo_top_VIA10 $T=50940 105540 0 0 $X=50470 $Y=105310
X9070 3 digital_ldo_top_VIA10 $T=50940 109620 0 0 $X=50470 $Y=109390
X9071 3 digital_ldo_top_VIA10 $T=50940 113700 0 0 $X=50470 $Y=113470
X9072 3 digital_ldo_top_VIA10 $T=50940 117780 0 0 $X=50470 $Y=117550
X9073 3 digital_ldo_top_VIA10 $T=50940 121860 0 0 $X=50470 $Y=121630
X9074 3 digital_ldo_top_VIA10 $T=50940 125940 0 0 $X=50470 $Y=125710
X9075 2 digital_ldo_top_VIA10 $T=52780 13060 0 0 $X=52310 $Y=12830
X9076 2 digital_ldo_top_VIA10 $T=52780 17140 0 0 $X=52310 $Y=16910
X9077 2 digital_ldo_top_VIA10 $T=52780 21220 0 0 $X=52310 $Y=20990
X9078 2 digital_ldo_top_VIA10 $T=52780 25300 0 0 $X=52310 $Y=25070
X9079 2 digital_ldo_top_VIA10 $T=52780 29380 0 0 $X=52310 $Y=29150
X9080 2 digital_ldo_top_VIA10 $T=52780 33460 0 0 $X=52310 $Y=33230
X9081 2 digital_ldo_top_VIA10 $T=52780 37540 0 0 $X=52310 $Y=37310
X9082 2 digital_ldo_top_VIA10 $T=52780 41620 0 0 $X=52310 $Y=41390
X9083 2 digital_ldo_top_VIA10 $T=52780 45700 0 0 $X=52310 $Y=45470
X9084 2 digital_ldo_top_VIA10 $T=52780 49780 0 0 $X=52310 $Y=49550
X9085 2 digital_ldo_top_VIA10 $T=52780 53860 0 0 $X=52310 $Y=53630
X9086 2 digital_ldo_top_VIA10 $T=52780 57940 0 0 $X=52310 $Y=57710
X9087 2 digital_ldo_top_VIA10 $T=52780 62020 0 0 $X=52310 $Y=61790
X9088 2 digital_ldo_top_VIA10 $T=52780 66100 0 0 $X=52310 $Y=65870
X9089 2 digital_ldo_top_VIA10 $T=52780 70180 0 0 $X=52310 $Y=69950
X9090 2 digital_ldo_top_VIA10 $T=52780 74260 0 0 $X=52310 $Y=74030
X9091 2 digital_ldo_top_VIA10 $T=52780 78340 0 0 $X=52310 $Y=78110
X9092 2 digital_ldo_top_VIA10 $T=52780 82420 0 0 $X=52310 $Y=82190
X9093 2 digital_ldo_top_VIA10 $T=52780 86500 0 0 $X=52310 $Y=86270
X9094 2 digital_ldo_top_VIA10 $T=52780 90580 0 0 $X=52310 $Y=90350
X9095 2 digital_ldo_top_VIA10 $T=52780 94660 0 0 $X=52310 $Y=94430
X9096 2 digital_ldo_top_VIA10 $T=52780 98740 0 0 $X=52310 $Y=98510
X9097 2 digital_ldo_top_VIA10 $T=52780 102820 0 0 $X=52310 $Y=102590
X9098 2 digital_ldo_top_VIA10 $T=52780 106900 0 0 $X=52310 $Y=106670
X9099 2 digital_ldo_top_VIA10 $T=52780 110980 0 0 $X=52310 $Y=110750
X9100 2 digital_ldo_top_VIA10 $T=52780 115060 0 0 $X=52310 $Y=114830
X9101 2 digital_ldo_top_VIA10 $T=52780 119140 0 0 $X=52310 $Y=118910
X9102 2 digital_ldo_top_VIA10 $T=52780 123220 0 0 $X=52310 $Y=122990
X9103 2 digital_ldo_top_VIA10 $T=52780 127300 0 0 $X=52310 $Y=127070
X9104 3 digital_ldo_top_VIA10 $T=56460 11700 0 0 $X=55990 $Y=11470
X9105 3 digital_ldo_top_VIA10 $T=56460 15780 0 0 $X=55990 $Y=15550
X9106 3 digital_ldo_top_VIA10 $T=56460 19860 0 0 $X=55990 $Y=19630
X9107 3 digital_ldo_top_VIA10 $T=56460 23940 0 0 $X=55990 $Y=23710
X9108 3 digital_ldo_top_VIA10 $T=56460 28020 0 0 $X=55990 $Y=27790
X9109 3 digital_ldo_top_VIA10 $T=56460 32100 0 0 $X=55990 $Y=31870
X9110 3 digital_ldo_top_VIA10 $T=56460 36180 0 0 $X=55990 $Y=35950
X9111 3 digital_ldo_top_VIA10 $T=56460 40260 0 0 $X=55990 $Y=40030
X9112 3 digital_ldo_top_VIA10 $T=56460 44340 0 0 $X=55990 $Y=44110
X9113 3 digital_ldo_top_VIA10 $T=56460 48420 0 0 $X=55990 $Y=48190
X9114 3 digital_ldo_top_VIA10 $T=56460 52500 0 0 $X=55990 $Y=52270
X9115 3 digital_ldo_top_VIA10 $T=56460 56580 0 0 $X=55990 $Y=56350
X9116 3 digital_ldo_top_VIA10 $T=56460 60660 0 0 $X=55990 $Y=60430
X9117 3 digital_ldo_top_VIA10 $T=56460 64740 0 0 $X=55990 $Y=64510
X9118 3 digital_ldo_top_VIA10 $T=56460 68820 0 0 $X=55990 $Y=68590
X9119 3 digital_ldo_top_VIA10 $T=56460 72900 0 0 $X=55990 $Y=72670
X9120 3 digital_ldo_top_VIA10 $T=56460 76980 0 0 $X=55990 $Y=76750
X9121 3 digital_ldo_top_VIA10 $T=56460 81060 0 0 $X=55990 $Y=80830
X9122 3 digital_ldo_top_VIA10 $T=56460 85140 0 0 $X=55990 $Y=84910
X9123 3 digital_ldo_top_VIA10 $T=56460 89220 0 0 $X=55990 $Y=88990
X9124 3 digital_ldo_top_VIA10 $T=56460 93300 0 0 $X=55990 $Y=93070
X9125 3 digital_ldo_top_VIA10 $T=56460 97380 0 0 $X=55990 $Y=97150
X9126 3 digital_ldo_top_VIA10 $T=56460 101460 0 0 $X=55990 $Y=101230
X9127 3 digital_ldo_top_VIA10 $T=56460 105540 0 0 $X=55990 $Y=105310
X9128 3 digital_ldo_top_VIA10 $T=56460 109620 0 0 $X=55990 $Y=109390
X9129 3 digital_ldo_top_VIA10 $T=56460 113700 0 0 $X=55990 $Y=113470
X9130 3 digital_ldo_top_VIA10 $T=56460 117780 0 0 $X=55990 $Y=117550
X9131 3 digital_ldo_top_VIA10 $T=56460 121860 0 0 $X=55990 $Y=121630
X9132 3 digital_ldo_top_VIA10 $T=56460 125940 0 0 $X=55990 $Y=125710
X9133 2 digital_ldo_top_VIA10 $T=58300 13060 0 0 $X=57830 $Y=12830
X9134 2 digital_ldo_top_VIA10 $T=58300 17140 0 0 $X=57830 $Y=16910
X9135 2 digital_ldo_top_VIA10 $T=58300 21220 0 0 $X=57830 $Y=20990
X9136 2 digital_ldo_top_VIA10 $T=58300 25300 0 0 $X=57830 $Y=25070
X9137 2 digital_ldo_top_VIA10 $T=58300 29380 0 0 $X=57830 $Y=29150
X9138 2 digital_ldo_top_VIA10 $T=58300 33460 0 0 $X=57830 $Y=33230
X9139 2 digital_ldo_top_VIA10 $T=58300 37540 0 0 $X=57830 $Y=37310
X9140 2 digital_ldo_top_VIA10 $T=58300 41620 0 0 $X=57830 $Y=41390
X9141 2 digital_ldo_top_VIA10 $T=58300 45700 0 0 $X=57830 $Y=45470
X9142 2 digital_ldo_top_VIA10 $T=58300 49780 0 0 $X=57830 $Y=49550
X9143 2 digital_ldo_top_VIA10 $T=58300 53860 0 0 $X=57830 $Y=53630
X9144 2 digital_ldo_top_VIA10 $T=58300 57940 0 0 $X=57830 $Y=57710
X9145 2 digital_ldo_top_VIA10 $T=58300 62020 0 0 $X=57830 $Y=61790
X9146 2 digital_ldo_top_VIA10 $T=58300 66100 0 0 $X=57830 $Y=65870
X9147 2 digital_ldo_top_VIA10 $T=58300 70180 0 0 $X=57830 $Y=69950
X9148 2 digital_ldo_top_VIA10 $T=58300 74260 0 0 $X=57830 $Y=74030
X9149 2 digital_ldo_top_VIA10 $T=58300 78340 0 0 $X=57830 $Y=78110
X9150 2 digital_ldo_top_VIA10 $T=58300 82420 0 0 $X=57830 $Y=82190
X9151 2 digital_ldo_top_VIA10 $T=58300 86500 0 0 $X=57830 $Y=86270
X9152 2 digital_ldo_top_VIA10 $T=58300 90580 0 0 $X=57830 $Y=90350
X9153 2 digital_ldo_top_VIA10 $T=58300 94660 0 0 $X=57830 $Y=94430
X9154 2 digital_ldo_top_VIA10 $T=58300 98740 0 0 $X=57830 $Y=98510
X9155 2 digital_ldo_top_VIA10 $T=58300 102820 0 0 $X=57830 $Y=102590
X9156 2 digital_ldo_top_VIA10 $T=58300 106900 0 0 $X=57830 $Y=106670
X9157 2 digital_ldo_top_VIA10 $T=58300 110980 0 0 $X=57830 $Y=110750
X9158 2 digital_ldo_top_VIA10 $T=58300 115060 0 0 $X=57830 $Y=114830
X9159 2 digital_ldo_top_VIA10 $T=58300 119140 0 0 $X=57830 $Y=118910
X9160 2 digital_ldo_top_VIA10 $T=58300 123220 0 0 $X=57830 $Y=122990
X9161 2 digital_ldo_top_VIA10 $T=58300 127300 0 0 $X=57830 $Y=127070
X9162 3 digital_ldo_top_VIA10 $T=61980 11700 0 0 $X=61510 $Y=11470
X9163 3 digital_ldo_top_VIA10 $T=61980 15780 0 0 $X=61510 $Y=15550
X9164 3 digital_ldo_top_VIA10 $T=61980 19860 0 0 $X=61510 $Y=19630
X9165 3 digital_ldo_top_VIA10 $T=61980 23940 0 0 $X=61510 $Y=23710
X9166 3 digital_ldo_top_VIA10 $T=61980 28020 0 0 $X=61510 $Y=27790
X9167 3 digital_ldo_top_VIA10 $T=61980 32100 0 0 $X=61510 $Y=31870
X9168 3 digital_ldo_top_VIA10 $T=61980 36180 0 0 $X=61510 $Y=35950
X9169 3 digital_ldo_top_VIA10 $T=61980 40260 0 0 $X=61510 $Y=40030
X9170 3 digital_ldo_top_VIA10 $T=61980 44340 0 0 $X=61510 $Y=44110
X9171 3 digital_ldo_top_VIA10 $T=61980 48420 0 0 $X=61510 $Y=48190
X9172 3 digital_ldo_top_VIA10 $T=61980 52500 0 0 $X=61510 $Y=52270
X9173 3 digital_ldo_top_VIA10 $T=61980 56580 0 0 $X=61510 $Y=56350
X9174 3 digital_ldo_top_VIA10 $T=61980 60660 0 0 $X=61510 $Y=60430
X9175 3 digital_ldo_top_VIA10 $T=61980 64740 0 0 $X=61510 $Y=64510
X9176 3 digital_ldo_top_VIA10 $T=61980 68820 0 0 $X=61510 $Y=68590
X9177 3 digital_ldo_top_VIA10 $T=61980 72900 0 0 $X=61510 $Y=72670
X9178 3 digital_ldo_top_VIA10 $T=61980 76980 0 0 $X=61510 $Y=76750
X9179 3 digital_ldo_top_VIA10 $T=61980 81060 0 0 $X=61510 $Y=80830
X9180 3 digital_ldo_top_VIA10 $T=61980 85140 0 0 $X=61510 $Y=84910
X9181 3 digital_ldo_top_VIA10 $T=61980 89220 0 0 $X=61510 $Y=88990
X9182 3 digital_ldo_top_VIA10 $T=61980 93300 0 0 $X=61510 $Y=93070
X9183 3 digital_ldo_top_VIA10 $T=61980 97380 0 0 $X=61510 $Y=97150
X9184 3 digital_ldo_top_VIA10 $T=61980 101460 0 0 $X=61510 $Y=101230
X9185 3 digital_ldo_top_VIA10 $T=61980 105540 0 0 $X=61510 $Y=105310
X9186 3 digital_ldo_top_VIA10 $T=61980 109620 0 0 $X=61510 $Y=109390
X9187 3 digital_ldo_top_VIA10 $T=61980 113700 0 0 $X=61510 $Y=113470
X9188 3 digital_ldo_top_VIA10 $T=61980 117780 0 0 $X=61510 $Y=117550
X9189 3 digital_ldo_top_VIA10 $T=61980 121860 0 0 $X=61510 $Y=121630
X9190 3 digital_ldo_top_VIA10 $T=61980 125940 0 0 $X=61510 $Y=125710
X9191 2 digital_ldo_top_VIA10 $T=63820 13060 0 0 $X=63350 $Y=12830
X9192 2 digital_ldo_top_VIA10 $T=63820 17140 0 0 $X=63350 $Y=16910
X9193 2 digital_ldo_top_VIA10 $T=63820 21220 0 0 $X=63350 $Y=20990
X9194 2 digital_ldo_top_VIA10 $T=63820 25300 0 0 $X=63350 $Y=25070
X9195 2 digital_ldo_top_VIA10 $T=63820 29380 0 0 $X=63350 $Y=29150
X9196 2 digital_ldo_top_VIA10 $T=63820 33460 0 0 $X=63350 $Y=33230
X9197 2 digital_ldo_top_VIA10 $T=63820 37540 0 0 $X=63350 $Y=37310
X9198 2 digital_ldo_top_VIA10 $T=63820 41620 0 0 $X=63350 $Y=41390
X9199 2 digital_ldo_top_VIA10 $T=63820 45700 0 0 $X=63350 $Y=45470
X9200 2 digital_ldo_top_VIA10 $T=63820 49780 0 0 $X=63350 $Y=49550
X9201 2 digital_ldo_top_VIA10 $T=63820 53860 0 0 $X=63350 $Y=53630
X9202 2 digital_ldo_top_VIA10 $T=63820 57940 0 0 $X=63350 $Y=57710
X9203 2 digital_ldo_top_VIA10 $T=63820 62020 0 0 $X=63350 $Y=61790
X9204 2 digital_ldo_top_VIA10 $T=63820 66100 0 0 $X=63350 $Y=65870
X9205 2 digital_ldo_top_VIA10 $T=63820 70180 0 0 $X=63350 $Y=69950
X9206 2 digital_ldo_top_VIA10 $T=63820 74260 0 0 $X=63350 $Y=74030
X9207 2 digital_ldo_top_VIA10 $T=63820 78340 0 0 $X=63350 $Y=78110
X9208 2 digital_ldo_top_VIA10 $T=63820 82420 0 0 $X=63350 $Y=82190
X9209 2 digital_ldo_top_VIA10 $T=63820 86500 0 0 $X=63350 $Y=86270
X9210 2 digital_ldo_top_VIA10 $T=63820 90580 0 0 $X=63350 $Y=90350
X9211 2 digital_ldo_top_VIA10 $T=63820 94660 0 0 $X=63350 $Y=94430
X9212 2 digital_ldo_top_VIA10 $T=63820 98740 0 0 $X=63350 $Y=98510
X9213 2 digital_ldo_top_VIA10 $T=63820 102820 0 0 $X=63350 $Y=102590
X9214 2 digital_ldo_top_VIA10 $T=63820 106900 0 0 $X=63350 $Y=106670
X9215 2 digital_ldo_top_VIA10 $T=63820 110980 0 0 $X=63350 $Y=110750
X9216 2 digital_ldo_top_VIA10 $T=63820 115060 0 0 $X=63350 $Y=114830
X9217 2 digital_ldo_top_VIA10 $T=63820 119140 0 0 $X=63350 $Y=118910
X9218 2 digital_ldo_top_VIA10 $T=63820 123220 0 0 $X=63350 $Y=122990
X9219 2 digital_ldo_top_VIA10 $T=63820 127300 0 0 $X=63350 $Y=127070
X9220 3 digital_ldo_top_VIA10 $T=67500 11700 0 0 $X=67030 $Y=11470
X9221 3 digital_ldo_top_VIA10 $T=67500 15780 0 0 $X=67030 $Y=15550
X9222 3 digital_ldo_top_VIA10 $T=67500 19860 0 0 $X=67030 $Y=19630
X9223 3 digital_ldo_top_VIA10 $T=67500 23940 0 0 $X=67030 $Y=23710
X9224 3 digital_ldo_top_VIA10 $T=67500 28020 0 0 $X=67030 $Y=27790
X9225 3 digital_ldo_top_VIA10 $T=67500 32100 0 0 $X=67030 $Y=31870
X9226 3 digital_ldo_top_VIA10 $T=67500 36180 0 0 $X=67030 $Y=35950
X9227 3 digital_ldo_top_VIA10 $T=67500 40260 0 0 $X=67030 $Y=40030
X9228 3 digital_ldo_top_VIA10 $T=67500 44340 0 0 $X=67030 $Y=44110
X9229 3 digital_ldo_top_VIA10 $T=67500 48420 0 0 $X=67030 $Y=48190
X9230 3 digital_ldo_top_VIA10 $T=67500 52500 0 0 $X=67030 $Y=52270
X9231 3 digital_ldo_top_VIA10 $T=67500 56580 0 0 $X=67030 $Y=56350
X9232 3 digital_ldo_top_VIA10 $T=67500 60660 0 0 $X=67030 $Y=60430
X9233 3 digital_ldo_top_VIA10 $T=67500 64740 0 0 $X=67030 $Y=64510
X9234 3 digital_ldo_top_VIA10 $T=67500 68820 0 0 $X=67030 $Y=68590
X9235 3 digital_ldo_top_VIA10 $T=67500 72900 0 0 $X=67030 $Y=72670
X9236 3 digital_ldo_top_VIA10 $T=67500 76980 0 0 $X=67030 $Y=76750
X9237 3 digital_ldo_top_VIA10 $T=67500 81060 0 0 $X=67030 $Y=80830
X9238 3 digital_ldo_top_VIA10 $T=67500 85140 0 0 $X=67030 $Y=84910
X9239 3 digital_ldo_top_VIA10 $T=67500 89220 0 0 $X=67030 $Y=88990
X9240 3 digital_ldo_top_VIA10 $T=67500 93300 0 0 $X=67030 $Y=93070
X9241 3 digital_ldo_top_VIA10 $T=67500 97380 0 0 $X=67030 $Y=97150
X9242 3 digital_ldo_top_VIA10 $T=67500 101460 0 0 $X=67030 $Y=101230
X9243 3 digital_ldo_top_VIA10 $T=67500 105540 0 0 $X=67030 $Y=105310
X9244 3 digital_ldo_top_VIA10 $T=67500 109620 0 0 $X=67030 $Y=109390
X9245 3 digital_ldo_top_VIA10 $T=67500 113700 0 0 $X=67030 $Y=113470
X9246 3 digital_ldo_top_VIA10 $T=67500 117780 0 0 $X=67030 $Y=117550
X9247 3 digital_ldo_top_VIA10 $T=67500 121860 0 0 $X=67030 $Y=121630
X9248 3 digital_ldo_top_VIA10 $T=67500 125940 0 0 $X=67030 $Y=125710
X9249 2 digital_ldo_top_VIA10 $T=69340 13060 0 0 $X=68870 $Y=12830
X9250 2 digital_ldo_top_VIA10 $T=69340 17140 0 0 $X=68870 $Y=16910
X9251 2 digital_ldo_top_VIA10 $T=69340 21220 0 0 $X=68870 $Y=20990
X9252 2 digital_ldo_top_VIA10 $T=69340 25300 0 0 $X=68870 $Y=25070
X9253 2 digital_ldo_top_VIA10 $T=69340 29380 0 0 $X=68870 $Y=29150
X9254 2 digital_ldo_top_VIA10 $T=69340 33460 0 0 $X=68870 $Y=33230
X9255 2 digital_ldo_top_VIA10 $T=69340 37540 0 0 $X=68870 $Y=37310
X9256 2 digital_ldo_top_VIA10 $T=69340 41620 0 0 $X=68870 $Y=41390
X9257 2 digital_ldo_top_VIA10 $T=69340 45700 0 0 $X=68870 $Y=45470
X9258 2 digital_ldo_top_VIA10 $T=69340 49780 0 0 $X=68870 $Y=49550
X9259 2 digital_ldo_top_VIA10 $T=69340 53860 0 0 $X=68870 $Y=53630
X9260 2 digital_ldo_top_VIA10 $T=69340 57940 0 0 $X=68870 $Y=57710
X9261 2 digital_ldo_top_VIA10 $T=69340 62020 0 0 $X=68870 $Y=61790
X9262 2 digital_ldo_top_VIA10 $T=69340 66100 0 0 $X=68870 $Y=65870
X9263 2 digital_ldo_top_VIA10 $T=69340 70180 0 0 $X=68870 $Y=69950
X9264 2 digital_ldo_top_VIA10 $T=69340 74260 0 0 $X=68870 $Y=74030
X9265 2 digital_ldo_top_VIA10 $T=69340 78340 0 0 $X=68870 $Y=78110
X9266 2 digital_ldo_top_VIA10 $T=69340 82420 0 0 $X=68870 $Y=82190
X9267 2 digital_ldo_top_VIA10 $T=69340 86500 0 0 $X=68870 $Y=86270
X9268 2 digital_ldo_top_VIA10 $T=69340 90580 0 0 $X=68870 $Y=90350
X9269 2 digital_ldo_top_VIA10 $T=69340 94660 0 0 $X=68870 $Y=94430
X9270 2 digital_ldo_top_VIA10 $T=69340 98740 0 0 $X=68870 $Y=98510
X9271 2 digital_ldo_top_VIA10 $T=69340 102820 0 0 $X=68870 $Y=102590
X9272 2 digital_ldo_top_VIA10 $T=69340 106900 0 0 $X=68870 $Y=106670
X9273 2 digital_ldo_top_VIA10 $T=69340 110980 0 0 $X=68870 $Y=110750
X9274 2 digital_ldo_top_VIA10 $T=69340 115060 0 0 $X=68870 $Y=114830
X9275 2 digital_ldo_top_VIA10 $T=69340 119140 0 0 $X=68870 $Y=118910
X9276 2 digital_ldo_top_VIA10 $T=69340 123220 0 0 $X=68870 $Y=122990
X9277 2 digital_ldo_top_VIA10 $T=69340 127300 0 0 $X=68870 $Y=127070
X9278 3 digital_ldo_top_VIA10 $T=73020 11700 0 0 $X=72550 $Y=11470
X9279 3 digital_ldo_top_VIA10 $T=73020 15780 0 0 $X=72550 $Y=15550
X9280 3 digital_ldo_top_VIA10 $T=73020 19860 0 0 $X=72550 $Y=19630
X9281 3 digital_ldo_top_VIA10 $T=73020 23940 0 0 $X=72550 $Y=23710
X9282 3 digital_ldo_top_VIA10 $T=73020 28020 0 0 $X=72550 $Y=27790
X9283 3 digital_ldo_top_VIA10 $T=73020 32100 0 0 $X=72550 $Y=31870
X9284 3 digital_ldo_top_VIA10 $T=73020 36180 0 0 $X=72550 $Y=35950
X9285 3 digital_ldo_top_VIA10 $T=73020 40260 0 0 $X=72550 $Y=40030
X9286 3 digital_ldo_top_VIA10 $T=73020 44340 0 0 $X=72550 $Y=44110
X9287 3 digital_ldo_top_VIA10 $T=73020 48420 0 0 $X=72550 $Y=48190
X9288 3 digital_ldo_top_VIA10 $T=73020 52500 0 0 $X=72550 $Y=52270
X9289 3 digital_ldo_top_VIA10 $T=73020 56580 0 0 $X=72550 $Y=56350
X9290 3 digital_ldo_top_VIA10 $T=73020 60660 0 0 $X=72550 $Y=60430
X9291 3 digital_ldo_top_VIA10 $T=73020 64740 0 0 $X=72550 $Y=64510
X9292 3 digital_ldo_top_VIA10 $T=73020 68820 0 0 $X=72550 $Y=68590
X9293 3 digital_ldo_top_VIA10 $T=73020 72900 0 0 $X=72550 $Y=72670
X9294 3 digital_ldo_top_VIA10 $T=73020 76980 0 0 $X=72550 $Y=76750
X9295 3 digital_ldo_top_VIA10 $T=73020 81060 0 0 $X=72550 $Y=80830
X9296 3 digital_ldo_top_VIA10 $T=73020 85140 0 0 $X=72550 $Y=84910
X9297 3 digital_ldo_top_VIA10 $T=73020 89220 0 0 $X=72550 $Y=88990
X9298 3 digital_ldo_top_VIA10 $T=73020 93300 0 0 $X=72550 $Y=93070
X9299 3 digital_ldo_top_VIA10 $T=73020 97380 0 0 $X=72550 $Y=97150
X9300 3 digital_ldo_top_VIA10 $T=73020 101460 0 0 $X=72550 $Y=101230
X9301 3 digital_ldo_top_VIA10 $T=73020 105540 0 0 $X=72550 $Y=105310
X9302 3 digital_ldo_top_VIA10 $T=73020 109620 0 0 $X=72550 $Y=109390
X9303 3 digital_ldo_top_VIA10 $T=73020 113700 0 0 $X=72550 $Y=113470
X9304 3 digital_ldo_top_VIA10 $T=73020 117780 0 0 $X=72550 $Y=117550
X9305 3 digital_ldo_top_VIA10 $T=73020 121860 0 0 $X=72550 $Y=121630
X9306 3 digital_ldo_top_VIA10 $T=73020 125940 0 0 $X=72550 $Y=125710
X9307 2 digital_ldo_top_VIA10 $T=74860 13060 0 0 $X=74390 $Y=12830
X9308 2 digital_ldo_top_VIA10 $T=74860 17140 0 0 $X=74390 $Y=16910
X9309 2 digital_ldo_top_VIA10 $T=74860 21220 0 0 $X=74390 $Y=20990
X9310 2 digital_ldo_top_VIA10 $T=74860 25300 0 0 $X=74390 $Y=25070
X9311 2 digital_ldo_top_VIA10 $T=74860 29380 0 0 $X=74390 $Y=29150
X9312 2 digital_ldo_top_VIA10 $T=74860 33460 0 0 $X=74390 $Y=33230
X9313 2 digital_ldo_top_VIA10 $T=74860 37540 0 0 $X=74390 $Y=37310
X9314 2 digital_ldo_top_VIA10 $T=74860 41620 0 0 $X=74390 $Y=41390
X9315 2 digital_ldo_top_VIA10 $T=74860 45700 0 0 $X=74390 $Y=45470
X9316 2 digital_ldo_top_VIA10 $T=74860 49780 0 0 $X=74390 $Y=49550
X9317 2 digital_ldo_top_VIA10 $T=74860 53860 0 0 $X=74390 $Y=53630
X9318 2 digital_ldo_top_VIA10 $T=74860 57940 0 0 $X=74390 $Y=57710
X9319 2 digital_ldo_top_VIA10 $T=74860 62020 0 0 $X=74390 $Y=61790
X9320 2 digital_ldo_top_VIA10 $T=74860 66100 0 0 $X=74390 $Y=65870
X9321 2 digital_ldo_top_VIA10 $T=74860 70180 0 0 $X=74390 $Y=69950
X9322 2 digital_ldo_top_VIA10 $T=74860 74260 0 0 $X=74390 $Y=74030
X9323 2 digital_ldo_top_VIA10 $T=74860 78340 0 0 $X=74390 $Y=78110
X9324 2 digital_ldo_top_VIA10 $T=74860 82420 0 0 $X=74390 $Y=82190
X9325 2 digital_ldo_top_VIA10 $T=74860 86500 0 0 $X=74390 $Y=86270
X9326 2 digital_ldo_top_VIA10 $T=74860 90580 0 0 $X=74390 $Y=90350
X9327 2 digital_ldo_top_VIA10 $T=74860 94660 0 0 $X=74390 $Y=94430
X9328 2 digital_ldo_top_VIA10 $T=74860 98740 0 0 $X=74390 $Y=98510
X9329 2 digital_ldo_top_VIA10 $T=74860 102820 0 0 $X=74390 $Y=102590
X9330 2 digital_ldo_top_VIA10 $T=74860 106900 0 0 $X=74390 $Y=106670
X9331 2 digital_ldo_top_VIA10 $T=74860 110980 0 0 $X=74390 $Y=110750
X9332 2 digital_ldo_top_VIA10 $T=74860 115060 0 0 $X=74390 $Y=114830
X9333 2 digital_ldo_top_VIA10 $T=74860 119140 0 0 $X=74390 $Y=118910
X9334 2 digital_ldo_top_VIA10 $T=74860 123220 0 0 $X=74390 $Y=122990
X9335 2 digital_ldo_top_VIA10 $T=74860 127300 0 0 $X=74390 $Y=127070
X9336 3 digital_ldo_top_VIA10 $T=78540 11700 0 0 $X=78070 $Y=11470
X9337 3 digital_ldo_top_VIA10 $T=78540 15780 0 0 $X=78070 $Y=15550
X9338 3 digital_ldo_top_VIA10 $T=78540 19860 0 0 $X=78070 $Y=19630
X9339 3 digital_ldo_top_VIA10 $T=78540 23940 0 0 $X=78070 $Y=23710
X9340 3 digital_ldo_top_VIA10 $T=78540 28020 0 0 $X=78070 $Y=27790
X9341 3 digital_ldo_top_VIA10 $T=78540 32100 0 0 $X=78070 $Y=31870
X9342 3 digital_ldo_top_VIA10 $T=78540 36180 0 0 $X=78070 $Y=35950
X9343 3 digital_ldo_top_VIA10 $T=78540 40260 0 0 $X=78070 $Y=40030
X9344 3 digital_ldo_top_VIA10 $T=78540 44340 0 0 $X=78070 $Y=44110
X9345 3 digital_ldo_top_VIA10 $T=78540 48420 0 0 $X=78070 $Y=48190
X9346 3 digital_ldo_top_VIA10 $T=78540 52500 0 0 $X=78070 $Y=52270
X9347 3 digital_ldo_top_VIA10 $T=78540 56580 0 0 $X=78070 $Y=56350
X9348 3 digital_ldo_top_VIA10 $T=78540 60660 0 0 $X=78070 $Y=60430
X9349 3 digital_ldo_top_VIA10 $T=78540 64740 0 0 $X=78070 $Y=64510
X9350 3 digital_ldo_top_VIA10 $T=78540 68820 0 0 $X=78070 $Y=68590
X9351 3 digital_ldo_top_VIA10 $T=78540 72900 0 0 $X=78070 $Y=72670
X9352 3 digital_ldo_top_VIA10 $T=78540 76980 0 0 $X=78070 $Y=76750
X9353 3 digital_ldo_top_VIA10 $T=78540 81060 0 0 $X=78070 $Y=80830
X9354 3 digital_ldo_top_VIA10 $T=78540 85140 0 0 $X=78070 $Y=84910
X9355 3 digital_ldo_top_VIA10 $T=78540 89220 0 0 $X=78070 $Y=88990
X9356 3 digital_ldo_top_VIA10 $T=78540 93300 0 0 $X=78070 $Y=93070
X9357 3 digital_ldo_top_VIA10 $T=78540 97380 0 0 $X=78070 $Y=97150
X9358 3 digital_ldo_top_VIA10 $T=78540 101460 0 0 $X=78070 $Y=101230
X9359 3 digital_ldo_top_VIA10 $T=78540 105540 0 0 $X=78070 $Y=105310
X9360 3 digital_ldo_top_VIA10 $T=78540 109620 0 0 $X=78070 $Y=109390
X9361 3 digital_ldo_top_VIA10 $T=78540 113700 0 0 $X=78070 $Y=113470
X9362 3 digital_ldo_top_VIA10 $T=78540 117780 0 0 $X=78070 $Y=117550
X9363 3 digital_ldo_top_VIA10 $T=78540 121860 0 0 $X=78070 $Y=121630
X9364 3 digital_ldo_top_VIA10 $T=78540 125940 0 0 $X=78070 $Y=125710
X9365 2 digital_ldo_top_VIA10 $T=80380 13060 0 0 $X=79910 $Y=12830
X9366 2 digital_ldo_top_VIA10 $T=80380 17140 0 0 $X=79910 $Y=16910
X9367 2 digital_ldo_top_VIA10 $T=80380 21220 0 0 $X=79910 $Y=20990
X9368 2 digital_ldo_top_VIA10 $T=80380 25300 0 0 $X=79910 $Y=25070
X9369 2 digital_ldo_top_VIA10 $T=80380 29380 0 0 $X=79910 $Y=29150
X9370 2 digital_ldo_top_VIA10 $T=80380 33460 0 0 $X=79910 $Y=33230
X9371 2 digital_ldo_top_VIA10 $T=80380 37540 0 0 $X=79910 $Y=37310
X9372 2 digital_ldo_top_VIA10 $T=80380 41620 0 0 $X=79910 $Y=41390
X9373 2 digital_ldo_top_VIA10 $T=80380 45700 0 0 $X=79910 $Y=45470
X9374 2 digital_ldo_top_VIA10 $T=80380 49780 0 0 $X=79910 $Y=49550
X9375 2 digital_ldo_top_VIA10 $T=80380 53860 0 0 $X=79910 $Y=53630
X9376 2 digital_ldo_top_VIA10 $T=80380 57940 0 0 $X=79910 $Y=57710
X9377 2 digital_ldo_top_VIA10 $T=80380 62020 0 0 $X=79910 $Y=61790
X9378 2 digital_ldo_top_VIA10 $T=80380 66100 0 0 $X=79910 $Y=65870
X9379 2 digital_ldo_top_VIA10 $T=80380 70180 0 0 $X=79910 $Y=69950
X9380 2 digital_ldo_top_VIA10 $T=80380 74260 0 0 $X=79910 $Y=74030
X9381 2 digital_ldo_top_VIA10 $T=80380 78340 0 0 $X=79910 $Y=78110
X9382 2 digital_ldo_top_VIA10 $T=80380 82420 0 0 $X=79910 $Y=82190
X9383 2 digital_ldo_top_VIA10 $T=80380 86500 0 0 $X=79910 $Y=86270
X9384 2 digital_ldo_top_VIA10 $T=80380 90580 0 0 $X=79910 $Y=90350
X9385 2 digital_ldo_top_VIA10 $T=80380 94660 0 0 $X=79910 $Y=94430
X9386 2 digital_ldo_top_VIA10 $T=80380 98740 0 0 $X=79910 $Y=98510
X9387 2 digital_ldo_top_VIA10 $T=80380 102820 0 0 $X=79910 $Y=102590
X9388 2 digital_ldo_top_VIA10 $T=80380 106900 0 0 $X=79910 $Y=106670
X9389 2 digital_ldo_top_VIA10 $T=80380 110980 0 0 $X=79910 $Y=110750
X9390 2 digital_ldo_top_VIA10 $T=80380 115060 0 0 $X=79910 $Y=114830
X9391 2 digital_ldo_top_VIA10 $T=80380 119140 0 0 $X=79910 $Y=118910
X9392 2 digital_ldo_top_VIA10 $T=80380 123220 0 0 $X=79910 $Y=122990
X9393 2 digital_ldo_top_VIA10 $T=80380 127300 0 0 $X=79910 $Y=127070
X9394 3 digital_ldo_top_VIA10 $T=84060 11700 0 0 $X=83590 $Y=11470
X9395 3 digital_ldo_top_VIA10 $T=84060 15780 0 0 $X=83590 $Y=15550
X9396 3 digital_ldo_top_VIA10 $T=84060 19860 0 0 $X=83590 $Y=19630
X9397 3 digital_ldo_top_VIA10 $T=84060 23940 0 0 $X=83590 $Y=23710
X9398 3 digital_ldo_top_VIA10 $T=84060 28020 0 0 $X=83590 $Y=27790
X9399 3 digital_ldo_top_VIA10 $T=84060 32100 0 0 $X=83590 $Y=31870
X9400 3 digital_ldo_top_VIA10 $T=84060 36180 0 0 $X=83590 $Y=35950
X9401 3 digital_ldo_top_VIA10 $T=84060 40260 0 0 $X=83590 $Y=40030
X9402 3 digital_ldo_top_VIA10 $T=84060 44340 0 0 $X=83590 $Y=44110
X9403 3 digital_ldo_top_VIA10 $T=84060 48420 0 0 $X=83590 $Y=48190
X9404 3 digital_ldo_top_VIA10 $T=84060 52500 0 0 $X=83590 $Y=52270
X9405 3 digital_ldo_top_VIA10 $T=84060 56580 0 0 $X=83590 $Y=56350
X9406 3 digital_ldo_top_VIA10 $T=84060 60660 0 0 $X=83590 $Y=60430
X9407 3 digital_ldo_top_VIA10 $T=84060 64740 0 0 $X=83590 $Y=64510
X9408 3 digital_ldo_top_VIA10 $T=84060 68820 0 0 $X=83590 $Y=68590
X9409 3 digital_ldo_top_VIA10 $T=84060 72900 0 0 $X=83590 $Y=72670
X9410 3 digital_ldo_top_VIA10 $T=84060 76980 0 0 $X=83590 $Y=76750
X9411 3 digital_ldo_top_VIA10 $T=84060 81060 0 0 $X=83590 $Y=80830
X9412 3 digital_ldo_top_VIA10 $T=84060 85140 0 0 $X=83590 $Y=84910
X9413 3 digital_ldo_top_VIA10 $T=84060 89220 0 0 $X=83590 $Y=88990
X9414 3 digital_ldo_top_VIA10 $T=84060 93300 0 0 $X=83590 $Y=93070
X9415 3 digital_ldo_top_VIA10 $T=84060 97380 0 0 $X=83590 $Y=97150
X9416 3 digital_ldo_top_VIA10 $T=84060 101460 0 0 $X=83590 $Y=101230
X9417 3 digital_ldo_top_VIA10 $T=84060 105540 0 0 $X=83590 $Y=105310
X9418 3 digital_ldo_top_VIA10 $T=84060 109620 0 0 $X=83590 $Y=109390
X9419 3 digital_ldo_top_VIA10 $T=84060 113700 0 0 $X=83590 $Y=113470
X9420 3 digital_ldo_top_VIA10 $T=84060 117780 0 0 $X=83590 $Y=117550
X9421 3 digital_ldo_top_VIA10 $T=84060 121860 0 0 $X=83590 $Y=121630
X9422 3 digital_ldo_top_VIA10 $T=84060 125940 0 0 $X=83590 $Y=125710
X9423 2 digital_ldo_top_VIA10 $T=85900 13060 0 0 $X=85430 $Y=12830
X9424 2 digital_ldo_top_VIA10 $T=85900 17140 0 0 $X=85430 $Y=16910
X9425 2 digital_ldo_top_VIA10 $T=85900 21220 0 0 $X=85430 $Y=20990
X9426 2 digital_ldo_top_VIA10 $T=85900 25300 0 0 $X=85430 $Y=25070
X9427 2 digital_ldo_top_VIA10 $T=85900 29380 0 0 $X=85430 $Y=29150
X9428 2 digital_ldo_top_VIA10 $T=85900 33460 0 0 $X=85430 $Y=33230
X9429 2 digital_ldo_top_VIA10 $T=85900 37540 0 0 $X=85430 $Y=37310
X9430 2 digital_ldo_top_VIA10 $T=85900 41620 0 0 $X=85430 $Y=41390
X9431 2 digital_ldo_top_VIA10 $T=85900 45700 0 0 $X=85430 $Y=45470
X9432 2 digital_ldo_top_VIA10 $T=85900 49780 0 0 $X=85430 $Y=49550
X9433 2 digital_ldo_top_VIA10 $T=85900 53860 0 0 $X=85430 $Y=53630
X9434 2 digital_ldo_top_VIA10 $T=85900 57940 0 0 $X=85430 $Y=57710
X9435 2 digital_ldo_top_VIA10 $T=85900 62020 0 0 $X=85430 $Y=61790
X9436 2 digital_ldo_top_VIA10 $T=85900 66100 0 0 $X=85430 $Y=65870
X9437 2 digital_ldo_top_VIA10 $T=85900 70180 0 0 $X=85430 $Y=69950
X9438 2 digital_ldo_top_VIA10 $T=85900 74260 0 0 $X=85430 $Y=74030
X9439 2 digital_ldo_top_VIA10 $T=85900 78340 0 0 $X=85430 $Y=78110
X9440 2 digital_ldo_top_VIA10 $T=85900 82420 0 0 $X=85430 $Y=82190
X9441 2 digital_ldo_top_VIA10 $T=85900 86500 0 0 $X=85430 $Y=86270
X9442 2 digital_ldo_top_VIA10 $T=85900 90580 0 0 $X=85430 $Y=90350
X9443 2 digital_ldo_top_VIA10 $T=85900 94660 0 0 $X=85430 $Y=94430
X9444 2 digital_ldo_top_VIA10 $T=85900 98740 0 0 $X=85430 $Y=98510
X9445 2 digital_ldo_top_VIA10 $T=85900 102820 0 0 $X=85430 $Y=102590
X9446 2 digital_ldo_top_VIA10 $T=85900 106900 0 0 $X=85430 $Y=106670
X9447 2 digital_ldo_top_VIA10 $T=85900 110980 0 0 $X=85430 $Y=110750
X9448 2 digital_ldo_top_VIA10 $T=85900 115060 0 0 $X=85430 $Y=114830
X9449 2 digital_ldo_top_VIA10 $T=85900 119140 0 0 $X=85430 $Y=118910
X9450 2 digital_ldo_top_VIA10 $T=85900 123220 0 0 $X=85430 $Y=122990
X9451 2 digital_ldo_top_VIA10 $T=85900 127300 0 0 $X=85430 $Y=127070
X9452 3 digital_ldo_top_VIA10 $T=89580 11700 0 0 $X=89110 $Y=11470
X9453 3 digital_ldo_top_VIA10 $T=89580 15780 0 0 $X=89110 $Y=15550
X9454 3 digital_ldo_top_VIA10 $T=89580 19860 0 0 $X=89110 $Y=19630
X9455 3 digital_ldo_top_VIA10 $T=89580 23940 0 0 $X=89110 $Y=23710
X9456 3 digital_ldo_top_VIA10 $T=89580 28020 0 0 $X=89110 $Y=27790
X9457 3 digital_ldo_top_VIA10 $T=89580 32100 0 0 $X=89110 $Y=31870
X9458 3 digital_ldo_top_VIA10 $T=89580 36180 0 0 $X=89110 $Y=35950
X9459 3 digital_ldo_top_VIA10 $T=89580 40260 0 0 $X=89110 $Y=40030
X9460 3 digital_ldo_top_VIA10 $T=89580 44340 0 0 $X=89110 $Y=44110
X9461 3 digital_ldo_top_VIA10 $T=89580 48420 0 0 $X=89110 $Y=48190
X9462 3 digital_ldo_top_VIA10 $T=89580 52500 0 0 $X=89110 $Y=52270
X9463 3 digital_ldo_top_VIA10 $T=89580 56580 0 0 $X=89110 $Y=56350
X9464 3 digital_ldo_top_VIA10 $T=89580 60660 0 0 $X=89110 $Y=60430
X9465 3 digital_ldo_top_VIA10 $T=89580 64740 0 0 $X=89110 $Y=64510
X9466 3 digital_ldo_top_VIA10 $T=89580 68820 0 0 $X=89110 $Y=68590
X9467 3 digital_ldo_top_VIA10 $T=89580 72900 0 0 $X=89110 $Y=72670
X9468 3 digital_ldo_top_VIA10 $T=89580 76980 0 0 $X=89110 $Y=76750
X9469 3 digital_ldo_top_VIA10 $T=89580 81060 0 0 $X=89110 $Y=80830
X9470 3 digital_ldo_top_VIA10 $T=89580 85140 0 0 $X=89110 $Y=84910
X9471 3 digital_ldo_top_VIA10 $T=89580 89220 0 0 $X=89110 $Y=88990
X9472 3 digital_ldo_top_VIA10 $T=89580 93300 0 0 $X=89110 $Y=93070
X9473 3 digital_ldo_top_VIA10 $T=89580 97380 0 0 $X=89110 $Y=97150
X9474 3 digital_ldo_top_VIA10 $T=89580 101460 0 0 $X=89110 $Y=101230
X9475 3 digital_ldo_top_VIA10 $T=89580 105540 0 0 $X=89110 $Y=105310
X9476 3 digital_ldo_top_VIA10 $T=89580 109620 0 0 $X=89110 $Y=109390
X9477 3 digital_ldo_top_VIA10 $T=89580 113700 0 0 $X=89110 $Y=113470
X9478 3 digital_ldo_top_VIA10 $T=89580 117780 0 0 $X=89110 $Y=117550
X9479 3 digital_ldo_top_VIA10 $T=89580 121860 0 0 $X=89110 $Y=121630
X9480 3 digital_ldo_top_VIA10 $T=89580 125940 0 0 $X=89110 $Y=125710
X9481 2 digital_ldo_top_VIA10 $T=91420 13060 0 0 $X=90950 $Y=12830
X9482 2 digital_ldo_top_VIA10 $T=91420 17140 0 0 $X=90950 $Y=16910
X9483 2 digital_ldo_top_VIA10 $T=91420 21220 0 0 $X=90950 $Y=20990
X9484 2 digital_ldo_top_VIA10 $T=91420 25300 0 0 $X=90950 $Y=25070
X9485 2 digital_ldo_top_VIA10 $T=91420 29380 0 0 $X=90950 $Y=29150
X9486 2 digital_ldo_top_VIA10 $T=91420 33460 0 0 $X=90950 $Y=33230
X9487 2 digital_ldo_top_VIA10 $T=91420 37540 0 0 $X=90950 $Y=37310
X9488 2 digital_ldo_top_VIA10 $T=91420 41620 0 0 $X=90950 $Y=41390
X9489 2 digital_ldo_top_VIA10 $T=91420 45700 0 0 $X=90950 $Y=45470
X9490 2 digital_ldo_top_VIA10 $T=91420 49780 0 0 $X=90950 $Y=49550
X9491 2 digital_ldo_top_VIA10 $T=91420 53860 0 0 $X=90950 $Y=53630
X9492 2 digital_ldo_top_VIA10 $T=91420 57940 0 0 $X=90950 $Y=57710
X9493 2 digital_ldo_top_VIA10 $T=91420 62020 0 0 $X=90950 $Y=61790
X9494 2 digital_ldo_top_VIA10 $T=91420 66100 0 0 $X=90950 $Y=65870
X9495 2 digital_ldo_top_VIA10 $T=91420 70180 0 0 $X=90950 $Y=69950
X9496 2 digital_ldo_top_VIA10 $T=91420 74260 0 0 $X=90950 $Y=74030
X9497 2 digital_ldo_top_VIA10 $T=91420 78340 0 0 $X=90950 $Y=78110
X9498 2 digital_ldo_top_VIA10 $T=91420 82420 0 0 $X=90950 $Y=82190
X9499 2 digital_ldo_top_VIA10 $T=91420 86500 0 0 $X=90950 $Y=86270
X9500 2 digital_ldo_top_VIA10 $T=91420 90580 0 0 $X=90950 $Y=90350
X9501 2 digital_ldo_top_VIA10 $T=91420 94660 0 0 $X=90950 $Y=94430
X9502 2 digital_ldo_top_VIA10 $T=91420 98740 0 0 $X=90950 $Y=98510
X9503 2 digital_ldo_top_VIA10 $T=91420 102820 0 0 $X=90950 $Y=102590
X9504 2 digital_ldo_top_VIA10 $T=91420 106900 0 0 $X=90950 $Y=106670
X9505 2 digital_ldo_top_VIA10 $T=91420 110980 0 0 $X=90950 $Y=110750
X9506 2 digital_ldo_top_VIA10 $T=91420 115060 0 0 $X=90950 $Y=114830
X9507 2 digital_ldo_top_VIA10 $T=91420 119140 0 0 $X=90950 $Y=118910
X9508 2 digital_ldo_top_VIA10 $T=91420 123220 0 0 $X=90950 $Y=122990
X9509 2 digital_ldo_top_VIA10 $T=91420 127300 0 0 $X=90950 $Y=127070
X9510 3 digital_ldo_top_VIA10 $T=95100 11700 0 0 $X=94630 $Y=11470
X9511 3 digital_ldo_top_VIA10 $T=95100 15780 0 0 $X=94630 $Y=15550
X9512 3 digital_ldo_top_VIA10 $T=95100 19860 0 0 $X=94630 $Y=19630
X9513 3 digital_ldo_top_VIA10 $T=95100 23940 0 0 $X=94630 $Y=23710
X9514 3 digital_ldo_top_VIA10 $T=95100 28020 0 0 $X=94630 $Y=27790
X9515 3 digital_ldo_top_VIA10 $T=95100 32100 0 0 $X=94630 $Y=31870
X9516 3 digital_ldo_top_VIA10 $T=95100 36180 0 0 $X=94630 $Y=35950
X9517 3 digital_ldo_top_VIA10 $T=95100 40260 0 0 $X=94630 $Y=40030
X9518 3 digital_ldo_top_VIA10 $T=95100 44340 0 0 $X=94630 $Y=44110
X9519 3 digital_ldo_top_VIA10 $T=95100 48420 0 0 $X=94630 $Y=48190
X9520 3 digital_ldo_top_VIA10 $T=95100 52500 0 0 $X=94630 $Y=52270
X9521 3 digital_ldo_top_VIA10 $T=95100 56580 0 0 $X=94630 $Y=56350
X9522 3 digital_ldo_top_VIA10 $T=95100 60660 0 0 $X=94630 $Y=60430
X9523 3 digital_ldo_top_VIA10 $T=95100 64740 0 0 $X=94630 $Y=64510
X9524 3 digital_ldo_top_VIA10 $T=95100 68820 0 0 $X=94630 $Y=68590
X9525 3 digital_ldo_top_VIA10 $T=95100 72900 0 0 $X=94630 $Y=72670
X9526 3 digital_ldo_top_VIA10 $T=95100 76980 0 0 $X=94630 $Y=76750
X9527 3 digital_ldo_top_VIA10 $T=95100 81060 0 0 $X=94630 $Y=80830
X9528 3 digital_ldo_top_VIA10 $T=95100 85140 0 0 $X=94630 $Y=84910
X9529 3 digital_ldo_top_VIA10 $T=95100 89220 0 0 $X=94630 $Y=88990
X9530 3 digital_ldo_top_VIA10 $T=95100 93300 0 0 $X=94630 $Y=93070
X9531 3 digital_ldo_top_VIA10 $T=95100 97380 0 0 $X=94630 $Y=97150
X9532 3 digital_ldo_top_VIA10 $T=95100 101460 0 0 $X=94630 $Y=101230
X9533 3 digital_ldo_top_VIA10 $T=95100 105540 0 0 $X=94630 $Y=105310
X9534 3 digital_ldo_top_VIA10 $T=95100 109620 0 0 $X=94630 $Y=109390
X9535 3 digital_ldo_top_VIA10 $T=95100 113700 0 0 $X=94630 $Y=113470
X9536 3 digital_ldo_top_VIA10 $T=95100 117780 0 0 $X=94630 $Y=117550
X9537 3 digital_ldo_top_VIA10 $T=95100 121860 0 0 $X=94630 $Y=121630
X9538 3 digital_ldo_top_VIA10 $T=95100 125940 0 0 $X=94630 $Y=125710
X9539 2 digital_ldo_top_VIA10 $T=96940 13060 0 0 $X=96470 $Y=12830
X9540 2 digital_ldo_top_VIA10 $T=96940 17140 0 0 $X=96470 $Y=16910
X9541 2 digital_ldo_top_VIA10 $T=96940 21220 0 0 $X=96470 $Y=20990
X9542 2 digital_ldo_top_VIA10 $T=96940 25300 0 0 $X=96470 $Y=25070
X9543 2 digital_ldo_top_VIA10 $T=96940 29380 0 0 $X=96470 $Y=29150
X9544 2 digital_ldo_top_VIA10 $T=96940 33460 0 0 $X=96470 $Y=33230
X9545 2 digital_ldo_top_VIA10 $T=96940 37540 0 0 $X=96470 $Y=37310
X9546 2 digital_ldo_top_VIA10 $T=96940 41620 0 0 $X=96470 $Y=41390
X9547 2 digital_ldo_top_VIA10 $T=96940 45700 0 0 $X=96470 $Y=45470
X9548 2 digital_ldo_top_VIA10 $T=96940 49780 0 0 $X=96470 $Y=49550
X9549 2 digital_ldo_top_VIA10 $T=96940 53860 0 0 $X=96470 $Y=53630
X9550 2 digital_ldo_top_VIA10 $T=96940 57940 0 0 $X=96470 $Y=57710
X9551 2 digital_ldo_top_VIA10 $T=96940 62020 0 0 $X=96470 $Y=61790
X9552 2 digital_ldo_top_VIA10 $T=96940 66100 0 0 $X=96470 $Y=65870
X9553 2 digital_ldo_top_VIA10 $T=96940 70180 0 0 $X=96470 $Y=69950
X9554 2 digital_ldo_top_VIA10 $T=96940 74260 0 0 $X=96470 $Y=74030
X9555 2 digital_ldo_top_VIA10 $T=96940 78340 0 0 $X=96470 $Y=78110
X9556 2 digital_ldo_top_VIA10 $T=96940 82420 0 0 $X=96470 $Y=82190
X9557 2 digital_ldo_top_VIA10 $T=96940 86500 0 0 $X=96470 $Y=86270
X9558 2 digital_ldo_top_VIA10 $T=96940 90580 0 0 $X=96470 $Y=90350
X9559 2 digital_ldo_top_VIA10 $T=96940 94660 0 0 $X=96470 $Y=94430
X9560 2 digital_ldo_top_VIA10 $T=96940 98740 0 0 $X=96470 $Y=98510
X9561 2 digital_ldo_top_VIA10 $T=96940 102820 0 0 $X=96470 $Y=102590
X9562 2 digital_ldo_top_VIA10 $T=96940 106900 0 0 $X=96470 $Y=106670
X9563 2 digital_ldo_top_VIA10 $T=96940 110980 0 0 $X=96470 $Y=110750
X9564 2 digital_ldo_top_VIA10 $T=96940 115060 0 0 $X=96470 $Y=114830
X9565 2 digital_ldo_top_VIA10 $T=96940 119140 0 0 $X=96470 $Y=118910
X9566 2 digital_ldo_top_VIA10 $T=96940 123220 0 0 $X=96470 $Y=122990
X9567 2 digital_ldo_top_VIA10 $T=96940 127300 0 0 $X=96470 $Y=127070
X9568 3 digital_ldo_top_VIA10 $T=100620 11700 0 0 $X=100150 $Y=11470
X9569 3 digital_ldo_top_VIA10 $T=100620 15780 0 0 $X=100150 $Y=15550
X9570 3 digital_ldo_top_VIA10 $T=100620 19860 0 0 $X=100150 $Y=19630
X9571 3 digital_ldo_top_VIA10 $T=100620 23940 0 0 $X=100150 $Y=23710
X9572 3 digital_ldo_top_VIA10 $T=100620 28020 0 0 $X=100150 $Y=27790
X9573 3 digital_ldo_top_VIA10 $T=100620 32100 0 0 $X=100150 $Y=31870
X9574 3 digital_ldo_top_VIA10 $T=100620 36180 0 0 $X=100150 $Y=35950
X9575 3 digital_ldo_top_VIA10 $T=100620 40260 0 0 $X=100150 $Y=40030
X9576 3 digital_ldo_top_VIA10 $T=100620 44340 0 0 $X=100150 $Y=44110
X9577 3 digital_ldo_top_VIA10 $T=100620 48420 0 0 $X=100150 $Y=48190
X9578 3 digital_ldo_top_VIA10 $T=100620 52500 0 0 $X=100150 $Y=52270
X9579 3 digital_ldo_top_VIA10 $T=100620 56580 0 0 $X=100150 $Y=56350
X9580 3 digital_ldo_top_VIA10 $T=100620 60660 0 0 $X=100150 $Y=60430
X9581 3 digital_ldo_top_VIA10 $T=100620 64740 0 0 $X=100150 $Y=64510
X9582 3 digital_ldo_top_VIA10 $T=100620 68820 0 0 $X=100150 $Y=68590
X9583 3 digital_ldo_top_VIA10 $T=100620 72900 0 0 $X=100150 $Y=72670
X9584 3 digital_ldo_top_VIA10 $T=100620 76980 0 0 $X=100150 $Y=76750
X9585 3 digital_ldo_top_VIA10 $T=100620 81060 0 0 $X=100150 $Y=80830
X9586 3 digital_ldo_top_VIA10 $T=100620 85140 0 0 $X=100150 $Y=84910
X9587 3 digital_ldo_top_VIA10 $T=100620 89220 0 0 $X=100150 $Y=88990
X9588 3 digital_ldo_top_VIA10 $T=100620 93300 0 0 $X=100150 $Y=93070
X9589 3 digital_ldo_top_VIA10 $T=100620 97380 0 0 $X=100150 $Y=97150
X9590 3 digital_ldo_top_VIA10 $T=100620 101460 0 0 $X=100150 $Y=101230
X9591 3 digital_ldo_top_VIA10 $T=100620 105540 0 0 $X=100150 $Y=105310
X9592 3 digital_ldo_top_VIA10 $T=100620 109620 0 0 $X=100150 $Y=109390
X9593 3 digital_ldo_top_VIA10 $T=100620 113700 0 0 $X=100150 $Y=113470
X9594 3 digital_ldo_top_VIA10 $T=100620 117780 0 0 $X=100150 $Y=117550
X9595 3 digital_ldo_top_VIA10 $T=100620 121860 0 0 $X=100150 $Y=121630
X9596 3 digital_ldo_top_VIA10 $T=100620 125940 0 0 $X=100150 $Y=125710
X9597 2 digital_ldo_top_VIA10 $T=102460 13060 0 0 $X=101990 $Y=12830
X9598 2 digital_ldo_top_VIA10 $T=102460 17140 0 0 $X=101990 $Y=16910
X9599 2 digital_ldo_top_VIA10 $T=102460 21220 0 0 $X=101990 $Y=20990
X9600 2 digital_ldo_top_VIA10 $T=102460 25300 0 0 $X=101990 $Y=25070
X9601 2 digital_ldo_top_VIA10 $T=102460 29380 0 0 $X=101990 $Y=29150
X9602 2 digital_ldo_top_VIA10 $T=102460 33460 0 0 $X=101990 $Y=33230
X9603 2 digital_ldo_top_VIA10 $T=102460 37540 0 0 $X=101990 $Y=37310
X9604 2 digital_ldo_top_VIA10 $T=102460 41620 0 0 $X=101990 $Y=41390
X9605 2 digital_ldo_top_VIA10 $T=102460 45700 0 0 $X=101990 $Y=45470
X9606 2 digital_ldo_top_VIA10 $T=102460 49780 0 0 $X=101990 $Y=49550
X9607 2 digital_ldo_top_VIA10 $T=102460 53860 0 0 $X=101990 $Y=53630
X9608 2 digital_ldo_top_VIA10 $T=102460 57940 0 0 $X=101990 $Y=57710
X9609 2 digital_ldo_top_VIA10 $T=102460 62020 0 0 $X=101990 $Y=61790
X9610 2 digital_ldo_top_VIA10 $T=102460 66100 0 0 $X=101990 $Y=65870
X9611 2 digital_ldo_top_VIA10 $T=102460 70180 0 0 $X=101990 $Y=69950
X9612 2 digital_ldo_top_VIA10 $T=102460 74260 0 0 $X=101990 $Y=74030
X9613 2 digital_ldo_top_VIA10 $T=102460 78340 0 0 $X=101990 $Y=78110
X9614 2 digital_ldo_top_VIA10 $T=102460 82420 0 0 $X=101990 $Y=82190
X9615 2 digital_ldo_top_VIA10 $T=102460 86500 0 0 $X=101990 $Y=86270
X9616 2 digital_ldo_top_VIA10 $T=102460 90580 0 0 $X=101990 $Y=90350
X9617 2 digital_ldo_top_VIA10 $T=102460 94660 0 0 $X=101990 $Y=94430
X9618 2 digital_ldo_top_VIA10 $T=102460 98740 0 0 $X=101990 $Y=98510
X9619 2 digital_ldo_top_VIA10 $T=102460 102820 0 0 $X=101990 $Y=102590
X9620 2 digital_ldo_top_VIA10 $T=102460 106900 0 0 $X=101990 $Y=106670
X9621 2 digital_ldo_top_VIA10 $T=102460 110980 0 0 $X=101990 $Y=110750
X9622 2 digital_ldo_top_VIA10 $T=102460 115060 0 0 $X=101990 $Y=114830
X9623 2 digital_ldo_top_VIA10 $T=102460 119140 0 0 $X=101990 $Y=118910
X9624 2 digital_ldo_top_VIA10 $T=102460 123220 0 0 $X=101990 $Y=122990
X9625 2 digital_ldo_top_VIA10 $T=102460 127300 0 0 $X=101990 $Y=127070
X9626 3 digital_ldo_top_VIA10 $T=106140 11700 0 0 $X=105670 $Y=11470
X9627 3 digital_ldo_top_VIA10 $T=106140 15780 0 0 $X=105670 $Y=15550
X9628 3 digital_ldo_top_VIA10 $T=106140 19860 0 0 $X=105670 $Y=19630
X9629 3 digital_ldo_top_VIA10 $T=106140 23940 0 0 $X=105670 $Y=23710
X9630 3 digital_ldo_top_VIA10 $T=106140 32100 0 0 $X=105670 $Y=31870
X9631 3 digital_ldo_top_VIA10 $T=106140 85140 0 0 $X=105670 $Y=84910
X9632 3 digital_ldo_top_VIA10 $T=106140 89220 0 0 $X=105670 $Y=88990
X9633 3 digital_ldo_top_VIA10 $T=106140 93300 0 0 $X=105670 $Y=93070
X9634 3 digital_ldo_top_VIA10 $T=106140 97380 0 0 $X=105670 $Y=97150
X9635 3 digital_ldo_top_VIA10 $T=106140 101460 0 0 $X=105670 $Y=101230
X9636 3 digital_ldo_top_VIA10 $T=106140 105540 0 0 $X=105670 $Y=105310
X9637 3 digital_ldo_top_VIA10 $T=106140 109620 0 0 $X=105670 $Y=109390
X9638 3 digital_ldo_top_VIA10 $T=106140 113700 0 0 $X=105670 $Y=113470
X9639 3 digital_ldo_top_VIA10 $T=106140 117780 0 0 $X=105670 $Y=117550
X9640 3 digital_ldo_top_VIA10 $T=106140 121860 0 0 $X=105670 $Y=121630
X9641 3 digital_ldo_top_VIA10 $T=106140 125940 0 0 $X=105670 $Y=125710
X9642 2 digital_ldo_top_VIA10 $T=107980 13060 0 0 $X=107510 $Y=12830
X9643 2 digital_ldo_top_VIA10 $T=107980 17140 0 0 $X=107510 $Y=16910
X9644 2 digital_ldo_top_VIA10 $T=107980 21220 0 0 $X=107510 $Y=20990
X9645 2 digital_ldo_top_VIA10 $T=107980 25300 0 0 $X=107510 $Y=25070
X9646 2 digital_ldo_top_VIA10 $T=107980 86500 0 0 $X=107510 $Y=86270
X9647 2 digital_ldo_top_VIA10 $T=107980 90580 0 0 $X=107510 $Y=90350
X9648 2 digital_ldo_top_VIA10 $T=107980 94660 0 0 $X=107510 $Y=94430
X9649 2 digital_ldo_top_VIA10 $T=107980 98740 0 0 $X=107510 $Y=98510
X9650 2 digital_ldo_top_VIA10 $T=107980 102820 0 0 $X=107510 $Y=102590
X9651 2 digital_ldo_top_VIA10 $T=107980 106900 0 0 $X=107510 $Y=106670
X9652 2 digital_ldo_top_VIA10 $T=107980 110980 0 0 $X=107510 $Y=110750
X9653 2 digital_ldo_top_VIA10 $T=107980 115060 0 0 $X=107510 $Y=114830
X9654 2 digital_ldo_top_VIA10 $T=107980 119140 0 0 $X=107510 $Y=118910
X9655 2 digital_ldo_top_VIA10 $T=107980 123220 0 0 $X=107510 $Y=122990
X9656 2 digital_ldo_top_VIA10 $T=107980 127300 0 0 $X=107510 $Y=127070
X9657 3 digital_ldo_top_VIA10 $T=111660 11700 0 0 $X=111190 $Y=11470
X9658 3 digital_ldo_top_VIA10 $T=111660 15780 0 0 $X=111190 $Y=15550
X9659 3 digital_ldo_top_VIA10 $T=111660 19860 0 0 $X=111190 $Y=19630
X9660 3 digital_ldo_top_VIA10 $T=111660 23940 0 0 $X=111190 $Y=23710
X9661 3 digital_ldo_top_VIA10 $T=111660 32100 0 0 $X=111190 $Y=31870
X9662 3 digital_ldo_top_VIA10 $T=111660 85140 0 0 $X=111190 $Y=84910
X9663 3 digital_ldo_top_VIA10 $T=111660 89220 0 0 $X=111190 $Y=88990
X9664 3 digital_ldo_top_VIA10 $T=111660 93300 0 0 $X=111190 $Y=93070
X9665 3 digital_ldo_top_VIA10 $T=111660 97380 0 0 $X=111190 $Y=97150
X9666 3 digital_ldo_top_VIA10 $T=111660 101460 0 0 $X=111190 $Y=101230
X9667 3 digital_ldo_top_VIA10 $T=111660 105540 0 0 $X=111190 $Y=105310
X9668 3 digital_ldo_top_VIA10 $T=111660 109620 0 0 $X=111190 $Y=109390
X9669 3 digital_ldo_top_VIA10 $T=111660 113700 0 0 $X=111190 $Y=113470
X9670 3 digital_ldo_top_VIA10 $T=111660 117780 0 0 $X=111190 $Y=117550
X9671 3 digital_ldo_top_VIA10 $T=111660 121860 0 0 $X=111190 $Y=121630
X9672 3 digital_ldo_top_VIA10 $T=111660 125940 0 0 $X=111190 $Y=125710
X9673 2 digital_ldo_top_VIA10 $T=113500 13060 0 0 $X=113030 $Y=12830
X9674 2 digital_ldo_top_VIA10 $T=113500 17140 0 0 $X=113030 $Y=16910
X9675 2 digital_ldo_top_VIA10 $T=113500 21220 0 0 $X=113030 $Y=20990
X9676 2 digital_ldo_top_VIA10 $T=113500 25300 0 0 $X=113030 $Y=25070
X9677 2 digital_ldo_top_VIA10 $T=113500 86500 0 0 $X=113030 $Y=86270
X9678 2 digital_ldo_top_VIA10 $T=113500 90580 0 0 $X=113030 $Y=90350
X9679 2 digital_ldo_top_VIA10 $T=113500 94660 0 0 $X=113030 $Y=94430
X9680 2 digital_ldo_top_VIA10 $T=113500 98740 0 0 $X=113030 $Y=98510
X9681 2 digital_ldo_top_VIA10 $T=113500 102820 0 0 $X=113030 $Y=102590
X9682 2 digital_ldo_top_VIA10 $T=113500 106900 0 0 $X=113030 $Y=106670
X9683 2 digital_ldo_top_VIA10 $T=113500 110980 0 0 $X=113030 $Y=110750
X9684 2 digital_ldo_top_VIA10 $T=113500 115060 0 0 $X=113030 $Y=114830
X9685 2 digital_ldo_top_VIA10 $T=113500 119140 0 0 $X=113030 $Y=118910
X9686 2 digital_ldo_top_VIA10 $T=113500 123220 0 0 $X=113030 $Y=122990
X9687 2 digital_ldo_top_VIA10 $T=113500 127300 0 0 $X=113030 $Y=127070
X9688 3 digital_ldo_top_VIA10 $T=117180 11700 0 0 $X=116710 $Y=11470
X9689 3 digital_ldo_top_VIA10 $T=117180 15780 0 0 $X=116710 $Y=15550
X9690 3 digital_ldo_top_VIA10 $T=117180 19860 0 0 $X=116710 $Y=19630
X9691 3 digital_ldo_top_VIA10 $T=117180 23940 0 0 $X=116710 $Y=23710
X9692 3 digital_ldo_top_VIA10 $T=117180 32100 0 0 $X=116710 $Y=31870
X9693 3 digital_ldo_top_VIA10 $T=117180 85140 0 0 $X=116710 $Y=84910
X9694 3 digital_ldo_top_VIA10 $T=117180 89220 0 0 $X=116710 $Y=88990
X9695 3 digital_ldo_top_VIA10 $T=117180 93300 0 0 $X=116710 $Y=93070
X9696 3 digital_ldo_top_VIA10 $T=117180 97380 0 0 $X=116710 $Y=97150
X9697 3 digital_ldo_top_VIA10 $T=117180 101460 0 0 $X=116710 $Y=101230
X9698 3 digital_ldo_top_VIA10 $T=117180 105540 0 0 $X=116710 $Y=105310
X9699 3 digital_ldo_top_VIA10 $T=117180 109620 0 0 $X=116710 $Y=109390
X9700 3 digital_ldo_top_VIA10 $T=117180 113700 0 0 $X=116710 $Y=113470
X9701 3 digital_ldo_top_VIA10 $T=117180 117780 0 0 $X=116710 $Y=117550
X9702 3 digital_ldo_top_VIA10 $T=117180 121860 0 0 $X=116710 $Y=121630
X9703 3 digital_ldo_top_VIA10 $T=117180 125940 0 0 $X=116710 $Y=125710
X9704 2 digital_ldo_top_VIA10 $T=119020 13060 0 0 $X=118550 $Y=12830
X9705 2 digital_ldo_top_VIA10 $T=119020 17140 0 0 $X=118550 $Y=16910
X9706 2 digital_ldo_top_VIA10 $T=119020 21220 0 0 $X=118550 $Y=20990
X9707 2 digital_ldo_top_VIA10 $T=119020 25300 0 0 $X=118550 $Y=25070
X9708 2 digital_ldo_top_VIA10 $T=119020 86500 0 0 $X=118550 $Y=86270
X9709 2 digital_ldo_top_VIA10 $T=119020 90580 0 0 $X=118550 $Y=90350
X9710 2 digital_ldo_top_VIA10 $T=119020 94660 0 0 $X=118550 $Y=94430
X9711 2 digital_ldo_top_VIA10 $T=119020 98740 0 0 $X=118550 $Y=98510
X9712 2 digital_ldo_top_VIA10 $T=119020 102820 0 0 $X=118550 $Y=102590
X9713 2 digital_ldo_top_VIA10 $T=119020 106900 0 0 $X=118550 $Y=106670
X9714 2 digital_ldo_top_VIA10 $T=119020 110980 0 0 $X=118550 $Y=110750
X9715 2 digital_ldo_top_VIA10 $T=119020 115060 0 0 $X=118550 $Y=114830
X9716 2 digital_ldo_top_VIA10 $T=119020 119140 0 0 $X=118550 $Y=118910
X9717 2 digital_ldo_top_VIA10 $T=119020 123220 0 0 $X=118550 $Y=122990
X9718 2 digital_ldo_top_VIA10 $T=119020 127300 0 0 $X=118550 $Y=127070
X9719 3 digital_ldo_top_VIA10 $T=122700 11700 0 0 $X=122230 $Y=11470
X9720 3 digital_ldo_top_VIA10 $T=122700 15780 0 0 $X=122230 $Y=15550
X9721 3 digital_ldo_top_VIA10 $T=122700 19860 0 0 $X=122230 $Y=19630
X9722 3 digital_ldo_top_VIA10 $T=122700 23940 0 0 $X=122230 $Y=23710
X9723 3 digital_ldo_top_VIA10 $T=122700 32100 0 0 $X=122230 $Y=31870
X9724 3 digital_ldo_top_VIA10 $T=122700 85140 0 0 $X=122230 $Y=84910
X9725 3 digital_ldo_top_VIA10 $T=122700 89220 0 0 $X=122230 $Y=88990
X9726 3 digital_ldo_top_VIA10 $T=122700 93300 0 0 $X=122230 $Y=93070
X9727 3 digital_ldo_top_VIA10 $T=122700 97380 0 0 $X=122230 $Y=97150
X9728 3 digital_ldo_top_VIA10 $T=122700 101460 0 0 $X=122230 $Y=101230
X9729 3 digital_ldo_top_VIA10 $T=122700 105540 0 0 $X=122230 $Y=105310
X9730 3 digital_ldo_top_VIA10 $T=122700 109620 0 0 $X=122230 $Y=109390
X9731 3 digital_ldo_top_VIA10 $T=122700 113700 0 0 $X=122230 $Y=113470
X9732 3 digital_ldo_top_VIA10 $T=122700 117780 0 0 $X=122230 $Y=117550
X9733 3 digital_ldo_top_VIA10 $T=122700 121860 0 0 $X=122230 $Y=121630
X9734 3 digital_ldo_top_VIA10 $T=122700 125940 0 0 $X=122230 $Y=125710
X9735 2 digital_ldo_top_VIA10 $T=124540 13060 0 0 $X=124070 $Y=12830
X9736 2 digital_ldo_top_VIA10 $T=124540 17140 0 0 $X=124070 $Y=16910
X9737 2 digital_ldo_top_VIA10 $T=124540 21220 0 0 $X=124070 $Y=20990
X9738 2 digital_ldo_top_VIA10 $T=124540 25300 0 0 $X=124070 $Y=25070
X9739 2 digital_ldo_top_VIA10 $T=124540 86500 0 0 $X=124070 $Y=86270
X9740 2 digital_ldo_top_VIA10 $T=124540 90580 0 0 $X=124070 $Y=90350
X9741 2 digital_ldo_top_VIA10 $T=124540 94660 0 0 $X=124070 $Y=94430
X9742 2 digital_ldo_top_VIA10 $T=124540 98740 0 0 $X=124070 $Y=98510
X9743 2 digital_ldo_top_VIA10 $T=124540 102820 0 0 $X=124070 $Y=102590
X9744 2 digital_ldo_top_VIA10 $T=124540 106900 0 0 $X=124070 $Y=106670
X9745 2 digital_ldo_top_VIA10 $T=124540 110980 0 0 $X=124070 $Y=110750
X9746 2 digital_ldo_top_VIA10 $T=124540 115060 0 0 $X=124070 $Y=114830
X9747 2 digital_ldo_top_VIA10 $T=124540 119140 0 0 $X=124070 $Y=118910
X9748 2 digital_ldo_top_VIA10 $T=124540 123220 0 0 $X=124070 $Y=122990
X9749 2 digital_ldo_top_VIA10 $T=124540 127300 0 0 $X=124070 $Y=127070
X9750 3 digital_ldo_top_VIA10 $T=128220 11700 0 0 $X=127750 $Y=11470
X9751 3 digital_ldo_top_VIA10 $T=128220 15780 0 0 $X=127750 $Y=15550
X9752 3 digital_ldo_top_VIA10 $T=128220 19860 0 0 $X=127750 $Y=19630
X9753 3 digital_ldo_top_VIA10 $T=128220 32100 0 0 $X=127750 $Y=31870
X9754 3 digital_ldo_top_VIA10 $T=128220 85140 0 0 $X=127750 $Y=84910
X9755 3 digital_ldo_top_VIA10 $T=128220 89220 0 0 $X=127750 $Y=88990
X9756 3 digital_ldo_top_VIA10 $T=128220 93300 0 0 $X=127750 $Y=93070
X9757 3 digital_ldo_top_VIA10 $T=128220 97380 0 0 $X=127750 $Y=97150
X9758 3 digital_ldo_top_VIA10 $T=128220 101460 0 0 $X=127750 $Y=101230
X9759 3 digital_ldo_top_VIA10 $T=128220 105540 0 0 $X=127750 $Y=105310
X9760 3 digital_ldo_top_VIA10 $T=128220 109620 0 0 $X=127750 $Y=109390
X9761 3 digital_ldo_top_VIA10 $T=128220 113700 0 0 $X=127750 $Y=113470
X9762 3 digital_ldo_top_VIA10 $T=128220 117780 0 0 $X=127750 $Y=117550
X9763 3 digital_ldo_top_VIA10 $T=128220 121860 0 0 $X=127750 $Y=121630
X9764 3 digital_ldo_top_VIA10 $T=128220 125940 0 0 $X=127750 $Y=125710
X9765 2 digital_ldo_top_VIA10 $T=130060 13060 0 0 $X=129590 $Y=12830
X9766 2 digital_ldo_top_VIA10 $T=130060 17140 0 0 $X=129590 $Y=16910
X9767 2 digital_ldo_top_VIA10 $T=130060 21220 0 0 $X=129590 $Y=20990
X9768 2 digital_ldo_top_VIA10 $T=130060 25300 0 0 $X=129590 $Y=25070
X9769 2 digital_ldo_top_VIA10 $T=130060 86500 0 0 $X=129590 $Y=86270
X9770 2 digital_ldo_top_VIA10 $T=130060 90580 0 0 $X=129590 $Y=90350
X9771 2 digital_ldo_top_VIA10 $T=130060 94660 0 0 $X=129590 $Y=94430
X9772 2 digital_ldo_top_VIA10 $T=130060 98740 0 0 $X=129590 $Y=98510
X9773 2 digital_ldo_top_VIA10 $T=130060 102820 0 0 $X=129590 $Y=102590
X9774 2 digital_ldo_top_VIA10 $T=130060 106900 0 0 $X=129590 $Y=106670
X9775 2 digital_ldo_top_VIA10 $T=130060 110980 0 0 $X=129590 $Y=110750
X9776 2 digital_ldo_top_VIA10 $T=130060 115060 0 0 $X=129590 $Y=114830
X9777 2 digital_ldo_top_VIA10 $T=130060 119140 0 0 $X=129590 $Y=118910
X9778 2 digital_ldo_top_VIA10 $T=130060 123220 0 0 $X=129590 $Y=122990
X9779 2 digital_ldo_top_VIA10 $T=130060 127300 0 0 $X=129590 $Y=127070
X9780 3 digital_ldo_top_VIA10 $T=133740 11700 0 0 $X=133270 $Y=11470
X9781 3 digital_ldo_top_VIA10 $T=133740 15780 0 0 $X=133270 $Y=15550
X9782 3 digital_ldo_top_VIA10 $T=133740 19860 0 0 $X=133270 $Y=19630
X9783 3 digital_ldo_top_VIA10 $T=133740 23940 0 0 $X=133270 $Y=23710
X9784 3 digital_ldo_top_VIA10 $T=133740 32100 0 0 $X=133270 $Y=31870
X9785 3 digital_ldo_top_VIA10 $T=133740 85140 0 0 $X=133270 $Y=84910
X9786 3 digital_ldo_top_VIA10 $T=133740 89220 0 0 $X=133270 $Y=88990
X9787 3 digital_ldo_top_VIA10 $T=133740 93300 0 0 $X=133270 $Y=93070
X9788 3 digital_ldo_top_VIA10 $T=133740 97380 0 0 $X=133270 $Y=97150
X9789 3 digital_ldo_top_VIA10 $T=133740 101460 0 0 $X=133270 $Y=101230
X9790 3 digital_ldo_top_VIA10 $T=133740 105540 0 0 $X=133270 $Y=105310
X9791 3 digital_ldo_top_VIA10 $T=133740 109620 0 0 $X=133270 $Y=109390
X9792 3 digital_ldo_top_VIA10 $T=133740 113700 0 0 $X=133270 $Y=113470
X9793 3 digital_ldo_top_VIA10 $T=133740 117780 0 0 $X=133270 $Y=117550
X9794 3 digital_ldo_top_VIA10 $T=133740 121860 0 0 $X=133270 $Y=121630
X9795 3 digital_ldo_top_VIA10 $T=133740 125940 0 0 $X=133270 $Y=125710
X9796 2 digital_ldo_top_VIA10 $T=135580 13060 0 0 $X=135110 $Y=12830
X9797 2 digital_ldo_top_VIA10 $T=135580 17140 0 0 $X=135110 $Y=16910
X9798 2 digital_ldo_top_VIA10 $T=135580 21220 0 0 $X=135110 $Y=20990
X9799 2 digital_ldo_top_VIA10 $T=135580 25300 0 0 $X=135110 $Y=25070
X9800 2 digital_ldo_top_VIA10 $T=135580 86500 0 0 $X=135110 $Y=86270
X9801 2 digital_ldo_top_VIA10 $T=135580 90580 0 0 $X=135110 $Y=90350
X9802 2 digital_ldo_top_VIA10 $T=135580 94660 0 0 $X=135110 $Y=94430
X9803 2 digital_ldo_top_VIA10 $T=135580 98740 0 0 $X=135110 $Y=98510
X9804 2 digital_ldo_top_VIA10 $T=135580 102820 0 0 $X=135110 $Y=102590
X9805 2 digital_ldo_top_VIA10 $T=135580 106900 0 0 $X=135110 $Y=106670
X9806 2 digital_ldo_top_VIA10 $T=135580 110980 0 0 $X=135110 $Y=110750
X9807 2 digital_ldo_top_VIA10 $T=135580 115060 0 0 $X=135110 $Y=114830
X9808 2 digital_ldo_top_VIA10 $T=135580 119140 0 0 $X=135110 $Y=118910
X9809 2 digital_ldo_top_VIA10 $T=135580 123220 0 0 $X=135110 $Y=122990
X9810 2 digital_ldo_top_VIA10 $T=135580 127300 0 0 $X=135110 $Y=127070
X9811 3 digital_ldo_top_VIA10 $T=139260 11700 0 0 $X=138790 $Y=11470
X9812 3 digital_ldo_top_VIA10 $T=139260 15780 0 0 $X=138790 $Y=15550
X9813 3 digital_ldo_top_VIA10 $T=139260 19860 0 0 $X=138790 $Y=19630
X9814 3 digital_ldo_top_VIA10 $T=139260 23940 0 0 $X=138790 $Y=23710
X9815 3 digital_ldo_top_VIA10 $T=139260 32100 0 0 $X=138790 $Y=31870
X9816 3 digital_ldo_top_VIA10 $T=139260 85140 0 0 $X=138790 $Y=84910
X9817 3 digital_ldo_top_VIA10 $T=139260 89220 0 0 $X=138790 $Y=88990
X9818 3 digital_ldo_top_VIA10 $T=139260 93300 0 0 $X=138790 $Y=93070
X9819 3 digital_ldo_top_VIA10 $T=139260 97380 0 0 $X=138790 $Y=97150
X9820 3 digital_ldo_top_VIA10 $T=139260 101460 0 0 $X=138790 $Y=101230
X9821 3 digital_ldo_top_VIA10 $T=139260 105540 0 0 $X=138790 $Y=105310
X9822 3 digital_ldo_top_VIA10 $T=139260 109620 0 0 $X=138790 $Y=109390
X9823 3 digital_ldo_top_VIA10 $T=139260 113700 0 0 $X=138790 $Y=113470
X9824 3 digital_ldo_top_VIA10 $T=139260 117780 0 0 $X=138790 $Y=117550
X9825 3 digital_ldo_top_VIA10 $T=139260 121860 0 0 $X=138790 $Y=121630
X9826 3 digital_ldo_top_VIA10 $T=139260 125940 0 0 $X=138790 $Y=125710
X9827 2 digital_ldo_top_VIA10 $T=141100 13060 0 0 $X=140630 $Y=12830
X9828 2 digital_ldo_top_VIA10 $T=141100 17140 0 0 $X=140630 $Y=16910
X9829 2 digital_ldo_top_VIA10 $T=141100 21220 0 0 $X=140630 $Y=20990
X9830 2 digital_ldo_top_VIA10 $T=141100 86500 0 0 $X=140630 $Y=86270
X9831 2 digital_ldo_top_VIA10 $T=141100 90580 0 0 $X=140630 $Y=90350
X9832 2 digital_ldo_top_VIA10 $T=141100 94660 0 0 $X=140630 $Y=94430
X9833 2 digital_ldo_top_VIA10 $T=141100 98740 0 0 $X=140630 $Y=98510
X9834 2 digital_ldo_top_VIA10 $T=141100 102820 0 0 $X=140630 $Y=102590
X9835 2 digital_ldo_top_VIA10 $T=141100 106900 0 0 $X=140630 $Y=106670
X9836 2 digital_ldo_top_VIA10 $T=141100 110980 0 0 $X=140630 $Y=110750
X9837 2 digital_ldo_top_VIA10 $T=141100 115060 0 0 $X=140630 $Y=114830
X9838 2 digital_ldo_top_VIA10 $T=141100 119140 0 0 $X=140630 $Y=118910
X9839 2 digital_ldo_top_VIA10 $T=141100 123220 0 0 $X=140630 $Y=122990
X9840 2 digital_ldo_top_VIA10 $T=141100 127300 0 0 $X=140630 $Y=127070
X9841 3 digital_ldo_top_VIA10 $T=144780 11700 0 0 $X=144310 $Y=11470
X9842 3 digital_ldo_top_VIA10 $T=144780 15780 0 0 $X=144310 $Y=15550
X9843 3 digital_ldo_top_VIA10 $T=144780 19860 0 0 $X=144310 $Y=19630
X9844 3 digital_ldo_top_VIA10 $T=144780 23940 0 0 $X=144310 $Y=23710
X9845 3 digital_ldo_top_VIA10 $T=144780 32100 0 0 $X=144310 $Y=31870
X9846 3 digital_ldo_top_VIA10 $T=144780 85140 0 0 $X=144310 $Y=84910
X9847 3 digital_ldo_top_VIA10 $T=144780 89220 0 0 $X=144310 $Y=88990
X9848 3 digital_ldo_top_VIA10 $T=144780 93300 0 0 $X=144310 $Y=93070
X9849 3 digital_ldo_top_VIA10 $T=144780 97380 0 0 $X=144310 $Y=97150
X9850 3 digital_ldo_top_VIA10 $T=144780 101460 0 0 $X=144310 $Y=101230
X9851 3 digital_ldo_top_VIA10 $T=144780 105540 0 0 $X=144310 $Y=105310
X9852 3 digital_ldo_top_VIA10 $T=144780 109620 0 0 $X=144310 $Y=109390
X9853 3 digital_ldo_top_VIA10 $T=144780 113700 0 0 $X=144310 $Y=113470
X9854 3 digital_ldo_top_VIA10 $T=144780 117780 0 0 $X=144310 $Y=117550
X9855 3 digital_ldo_top_VIA10 $T=144780 121860 0 0 $X=144310 $Y=121630
X9856 3 digital_ldo_top_VIA10 $T=144780 125940 0 0 $X=144310 $Y=125710
X9857 2 digital_ldo_top_VIA10 $T=146620 13060 0 0 $X=146150 $Y=12830
X9858 2 digital_ldo_top_VIA10 $T=146620 17140 0 0 $X=146150 $Y=16910
X9859 2 digital_ldo_top_VIA10 $T=146620 21220 0 0 $X=146150 $Y=20990
X9860 2 digital_ldo_top_VIA10 $T=146620 25300 0 0 $X=146150 $Y=25070
X9861 2 digital_ldo_top_VIA10 $T=146620 86500 0 0 $X=146150 $Y=86270
X9862 2 digital_ldo_top_VIA10 $T=146620 90580 0 0 $X=146150 $Y=90350
X9863 2 digital_ldo_top_VIA10 $T=146620 94660 0 0 $X=146150 $Y=94430
X9864 2 digital_ldo_top_VIA10 $T=146620 98740 0 0 $X=146150 $Y=98510
X9865 2 digital_ldo_top_VIA10 $T=146620 102820 0 0 $X=146150 $Y=102590
X9866 2 digital_ldo_top_VIA10 $T=146620 106900 0 0 $X=146150 $Y=106670
X9867 2 digital_ldo_top_VIA10 $T=146620 110980 0 0 $X=146150 $Y=110750
X9868 2 digital_ldo_top_VIA10 $T=146620 115060 0 0 $X=146150 $Y=114830
X9869 2 digital_ldo_top_VIA10 $T=146620 119140 0 0 $X=146150 $Y=118910
X9870 2 digital_ldo_top_VIA10 $T=146620 123220 0 0 $X=146150 $Y=122990
X9871 2 digital_ldo_top_VIA10 $T=146620 127300 0 0 $X=146150 $Y=127070
X9872 3 digital_ldo_top_VIA10 $T=150300 11700 0 0 $X=149830 $Y=11470
X9873 3 digital_ldo_top_VIA10 $T=150300 15780 0 0 $X=149830 $Y=15550
X9874 3 digital_ldo_top_VIA10 $T=150300 19860 0 0 $X=149830 $Y=19630
X9875 3 digital_ldo_top_VIA10 $T=150300 23940 0 0 $X=149830 $Y=23710
X9876 3 digital_ldo_top_VIA10 $T=150300 32100 0 0 $X=149830 $Y=31870
X9877 3 digital_ldo_top_VIA10 $T=150300 85140 0 0 $X=149830 $Y=84910
X9878 3 digital_ldo_top_VIA10 $T=150300 89220 0 0 $X=149830 $Y=88990
X9879 3 digital_ldo_top_VIA10 $T=150300 93300 0 0 $X=149830 $Y=93070
X9880 3 digital_ldo_top_VIA10 $T=150300 97380 0 0 $X=149830 $Y=97150
X9881 3 digital_ldo_top_VIA10 $T=150300 101460 0 0 $X=149830 $Y=101230
X9882 3 digital_ldo_top_VIA10 $T=150300 105540 0 0 $X=149830 $Y=105310
X9883 3 digital_ldo_top_VIA10 $T=150300 109620 0 0 $X=149830 $Y=109390
X9884 3 digital_ldo_top_VIA10 $T=150300 113700 0 0 $X=149830 $Y=113470
X9885 3 digital_ldo_top_VIA10 $T=150300 117780 0 0 $X=149830 $Y=117550
X9886 3 digital_ldo_top_VIA10 $T=150300 121860 0 0 $X=149830 $Y=121630
X9887 3 digital_ldo_top_VIA10 $T=150300 125940 0 0 $X=149830 $Y=125710
X9888 2 digital_ldo_top_VIA10 $T=152140 13060 0 0 $X=151670 $Y=12830
X9889 2 digital_ldo_top_VIA10 $T=152140 17140 0 0 $X=151670 $Y=16910
X9890 2 digital_ldo_top_VIA10 $T=152140 21220 0 0 $X=151670 $Y=20990
X9891 2 digital_ldo_top_VIA10 $T=152140 25300 0 0 $X=151670 $Y=25070
X9892 2 digital_ldo_top_VIA10 $T=152140 86500 0 0 $X=151670 $Y=86270
X9893 2 digital_ldo_top_VIA10 $T=152140 90580 0 0 $X=151670 $Y=90350
X9894 2 digital_ldo_top_VIA10 $T=152140 94660 0 0 $X=151670 $Y=94430
X9895 2 digital_ldo_top_VIA10 $T=152140 98740 0 0 $X=151670 $Y=98510
X9896 2 digital_ldo_top_VIA10 $T=152140 102820 0 0 $X=151670 $Y=102590
X9897 2 digital_ldo_top_VIA10 $T=152140 106900 0 0 $X=151670 $Y=106670
X9898 2 digital_ldo_top_VIA10 $T=152140 110980 0 0 $X=151670 $Y=110750
X9899 2 digital_ldo_top_VIA10 $T=152140 115060 0 0 $X=151670 $Y=114830
X9900 2 digital_ldo_top_VIA10 $T=152140 119140 0 0 $X=151670 $Y=118910
X9901 2 digital_ldo_top_VIA10 $T=152140 123220 0 0 $X=151670 $Y=122990
X9902 2 digital_ldo_top_VIA10 $T=152140 127300 0 0 $X=151670 $Y=127070
X9903 3 digital_ldo_top_VIA10 $T=155820 11700 0 0 $X=155350 $Y=11470
X9904 3 digital_ldo_top_VIA10 $T=155820 15780 0 0 $X=155350 $Y=15550
X9905 3 digital_ldo_top_VIA10 $T=155820 19860 0 0 $X=155350 $Y=19630
X9906 3 digital_ldo_top_VIA10 $T=155820 23940 0 0 $X=155350 $Y=23710
X9907 3 digital_ldo_top_VIA10 $T=155820 32100 0 0 $X=155350 $Y=31870
X9908 3 digital_ldo_top_VIA10 $T=155820 85140 0 0 $X=155350 $Y=84910
X9909 3 digital_ldo_top_VIA10 $T=155820 89220 0 0 $X=155350 $Y=88990
X9910 3 digital_ldo_top_VIA10 $T=155820 93300 0 0 $X=155350 $Y=93070
X9911 3 digital_ldo_top_VIA10 $T=155820 97380 0 0 $X=155350 $Y=97150
X9912 3 digital_ldo_top_VIA10 $T=155820 101460 0 0 $X=155350 $Y=101230
X9913 3 digital_ldo_top_VIA10 $T=155820 105540 0 0 $X=155350 $Y=105310
X9914 3 digital_ldo_top_VIA10 $T=155820 109620 0 0 $X=155350 $Y=109390
X9915 3 digital_ldo_top_VIA10 $T=155820 113700 0 0 $X=155350 $Y=113470
X9916 3 digital_ldo_top_VIA10 $T=155820 117780 0 0 $X=155350 $Y=117550
X9917 3 digital_ldo_top_VIA10 $T=155820 121860 0 0 $X=155350 $Y=121630
X9918 3 digital_ldo_top_VIA10 $T=155820 125940 0 0 $X=155350 $Y=125710
X9919 2 digital_ldo_top_VIA10 $T=157660 13060 0 0 $X=157190 $Y=12830
X9920 2 digital_ldo_top_VIA10 $T=157660 17140 0 0 $X=157190 $Y=16910
X9921 2 digital_ldo_top_VIA10 $T=157660 21220 0 0 $X=157190 $Y=20990
X9922 2 digital_ldo_top_VIA10 $T=157660 25300 0 0 $X=157190 $Y=25070
X9923 2 digital_ldo_top_VIA10 $T=157660 86500 0 0 $X=157190 $Y=86270
X9924 2 digital_ldo_top_VIA10 $T=157660 90580 0 0 $X=157190 $Y=90350
X9925 2 digital_ldo_top_VIA10 $T=157660 94660 0 0 $X=157190 $Y=94430
X9926 2 digital_ldo_top_VIA10 $T=157660 98740 0 0 $X=157190 $Y=98510
X9927 2 digital_ldo_top_VIA10 $T=157660 102820 0 0 $X=157190 $Y=102590
X9928 2 digital_ldo_top_VIA10 $T=157660 106900 0 0 $X=157190 $Y=106670
X9929 2 digital_ldo_top_VIA10 $T=157660 110980 0 0 $X=157190 $Y=110750
X9930 2 digital_ldo_top_VIA10 $T=157660 115060 0 0 $X=157190 $Y=114830
X9931 2 digital_ldo_top_VIA10 $T=157660 119140 0 0 $X=157190 $Y=118910
X9932 2 digital_ldo_top_VIA10 $T=157660 123220 0 0 $X=157190 $Y=122990
X9933 2 digital_ldo_top_VIA10 $T=157660 127300 0 0 $X=157190 $Y=127070
X9934 3 digital_ldo_top_VIA10 $T=161340 11700 0 0 $X=160870 $Y=11470
X9935 3 digital_ldo_top_VIA10 $T=161340 15780 0 0 $X=160870 $Y=15550
X9936 3 digital_ldo_top_VIA10 $T=161340 19860 0 0 $X=160870 $Y=19630
X9937 3 digital_ldo_top_VIA10 $T=161340 23940 0 0 $X=160870 $Y=23710
X9938 3 digital_ldo_top_VIA10 $T=161340 32100 0 0 $X=160870 $Y=31870
X9939 3 digital_ldo_top_VIA10 $T=161340 85140 0 0 $X=160870 $Y=84910
X9940 3 digital_ldo_top_VIA10 $T=161340 89220 0 0 $X=160870 $Y=88990
X9941 3 digital_ldo_top_VIA10 $T=161340 93300 0 0 $X=160870 $Y=93070
X9942 3 digital_ldo_top_VIA10 $T=161340 97380 0 0 $X=160870 $Y=97150
X9943 3 digital_ldo_top_VIA10 $T=161340 101460 0 0 $X=160870 $Y=101230
X9944 3 digital_ldo_top_VIA10 $T=161340 105540 0 0 $X=160870 $Y=105310
X9945 3 digital_ldo_top_VIA10 $T=161340 109620 0 0 $X=160870 $Y=109390
X9946 3 digital_ldo_top_VIA10 $T=161340 113700 0 0 $X=160870 $Y=113470
X9947 3 digital_ldo_top_VIA10 $T=161340 117780 0 0 $X=160870 $Y=117550
X9948 3 digital_ldo_top_VIA10 $T=161340 121860 0 0 $X=160870 $Y=121630
X9949 3 digital_ldo_top_VIA10 $T=161340 125940 0 0 $X=160870 $Y=125710
X9950 2 digital_ldo_top_VIA10 $T=163180 13060 0 0 $X=162710 $Y=12830
X9951 2 digital_ldo_top_VIA10 $T=163180 17140 0 0 $X=162710 $Y=16910
X9952 2 digital_ldo_top_VIA10 $T=163180 21220 0 0 $X=162710 $Y=20990
X9953 2 digital_ldo_top_VIA10 $T=163180 25300 0 0 $X=162710 $Y=25070
X9954 2 digital_ldo_top_VIA10 $T=163180 86500 0 0 $X=162710 $Y=86270
X9955 2 digital_ldo_top_VIA10 $T=163180 90580 0 0 $X=162710 $Y=90350
X9956 2 digital_ldo_top_VIA10 $T=163180 94660 0 0 $X=162710 $Y=94430
X9957 2 digital_ldo_top_VIA10 $T=163180 98740 0 0 $X=162710 $Y=98510
X9958 2 digital_ldo_top_VIA10 $T=163180 102820 0 0 $X=162710 $Y=102590
X9959 2 digital_ldo_top_VIA10 $T=163180 106900 0 0 $X=162710 $Y=106670
X9960 2 digital_ldo_top_VIA10 $T=163180 110980 0 0 $X=162710 $Y=110750
X9961 2 digital_ldo_top_VIA10 $T=163180 115060 0 0 $X=162710 $Y=114830
X9962 2 digital_ldo_top_VIA10 $T=163180 119140 0 0 $X=162710 $Y=118910
X9963 2 digital_ldo_top_VIA10 $T=163180 123220 0 0 $X=162710 $Y=122990
X9964 2 digital_ldo_top_VIA10 $T=163180 127300 0 0 $X=162710 $Y=127070
X9965 3 digital_ldo_top_VIA10 $T=166860 11700 0 0 $X=166390 $Y=11470
X9966 3 digital_ldo_top_VIA10 $T=166860 15780 0 0 $X=166390 $Y=15550
X9967 3 digital_ldo_top_VIA10 $T=166860 19860 0 0 $X=166390 $Y=19630
X9968 3 digital_ldo_top_VIA10 $T=166860 32100 0 0 $X=166390 $Y=31870
X9969 3 digital_ldo_top_VIA10 $T=166860 85140 0 0 $X=166390 $Y=84910
X9970 3 digital_ldo_top_VIA10 $T=166860 89220 0 0 $X=166390 $Y=88990
X9971 3 digital_ldo_top_VIA10 $T=166860 93300 0 0 $X=166390 $Y=93070
X9972 3 digital_ldo_top_VIA10 $T=166860 97380 0 0 $X=166390 $Y=97150
X9973 3 digital_ldo_top_VIA10 $T=166860 101460 0 0 $X=166390 $Y=101230
X9974 3 digital_ldo_top_VIA10 $T=166860 105540 0 0 $X=166390 $Y=105310
X9975 3 digital_ldo_top_VIA10 $T=166860 109620 0 0 $X=166390 $Y=109390
X9976 3 digital_ldo_top_VIA10 $T=166860 113700 0 0 $X=166390 $Y=113470
X9977 3 digital_ldo_top_VIA10 $T=166860 117780 0 0 $X=166390 $Y=117550
X9978 3 digital_ldo_top_VIA10 $T=166860 121860 0 0 $X=166390 $Y=121630
X9979 3 digital_ldo_top_VIA10 $T=166860 125940 0 0 $X=166390 $Y=125710
X9980 2 digital_ldo_top_VIA10 $T=168700 13060 0 0 $X=168230 $Y=12830
X9981 2 digital_ldo_top_VIA10 $T=168700 17140 0 0 $X=168230 $Y=16910
X9982 2 digital_ldo_top_VIA10 $T=168700 21220 0 0 $X=168230 $Y=20990
X9983 2 digital_ldo_top_VIA10 $T=168700 25300 0 0 $X=168230 $Y=25070
X9984 2 digital_ldo_top_VIA10 $T=168700 86500 0 0 $X=168230 $Y=86270
X9985 2 digital_ldo_top_VIA10 $T=168700 90580 0 0 $X=168230 $Y=90350
X9986 2 digital_ldo_top_VIA10 $T=168700 94660 0 0 $X=168230 $Y=94430
X9987 2 digital_ldo_top_VIA10 $T=168700 98740 0 0 $X=168230 $Y=98510
X9988 2 digital_ldo_top_VIA10 $T=168700 102820 0 0 $X=168230 $Y=102590
X9989 2 digital_ldo_top_VIA10 $T=168700 106900 0 0 $X=168230 $Y=106670
X9990 2 digital_ldo_top_VIA10 $T=168700 110980 0 0 $X=168230 $Y=110750
X9991 2 digital_ldo_top_VIA10 $T=168700 115060 0 0 $X=168230 $Y=114830
X9992 2 digital_ldo_top_VIA10 $T=168700 119140 0 0 $X=168230 $Y=118910
X9993 2 digital_ldo_top_VIA10 $T=168700 123220 0 0 $X=168230 $Y=122990
X9994 2 digital_ldo_top_VIA10 $T=168700 127300 0 0 $X=168230 $Y=127070
X9995 3 digital_ldo_top_VIA10 $T=172380 11700 0 0 $X=171910 $Y=11470
X9996 3 digital_ldo_top_VIA10 $T=172380 15780 0 0 $X=171910 $Y=15550
X9997 3 digital_ldo_top_VIA10 $T=172380 19860 0 0 $X=171910 $Y=19630
X9998 3 digital_ldo_top_VIA10 $T=172380 23940 0 0 $X=171910 $Y=23710
X9999 3 digital_ldo_top_VIA10 $T=172380 32100 0 0 $X=171910 $Y=31870
X10000 3 digital_ldo_top_VIA10 $T=172380 85140 0 0 $X=171910 $Y=84910
X10001 3 digital_ldo_top_VIA10 $T=172380 89220 0 0 $X=171910 $Y=88990
X10002 3 digital_ldo_top_VIA10 $T=172380 93300 0 0 $X=171910 $Y=93070
X10003 3 digital_ldo_top_VIA10 $T=172380 97380 0 0 $X=171910 $Y=97150
X10004 3 digital_ldo_top_VIA10 $T=172380 101460 0 0 $X=171910 $Y=101230
X10005 3 digital_ldo_top_VIA10 $T=172380 105540 0 0 $X=171910 $Y=105310
X10006 3 digital_ldo_top_VIA10 $T=172380 109620 0 0 $X=171910 $Y=109390
X10007 3 digital_ldo_top_VIA10 $T=172380 113700 0 0 $X=171910 $Y=113470
X10008 3 digital_ldo_top_VIA10 $T=172380 117780 0 0 $X=171910 $Y=117550
X10009 3 digital_ldo_top_VIA10 $T=172380 121860 0 0 $X=171910 $Y=121630
X10010 3 digital_ldo_top_VIA10 $T=172380 125940 0 0 $X=171910 $Y=125710
X10011 2 digital_ldo_top_VIA10 $T=174220 13060 0 0 $X=173750 $Y=12830
X10012 2 digital_ldo_top_VIA10 $T=174220 17140 0 0 $X=173750 $Y=16910
X10013 2 digital_ldo_top_VIA10 $T=174220 21220 0 0 $X=173750 $Y=20990
X10014 2 digital_ldo_top_VIA10 $T=174220 25300 0 0 $X=173750 $Y=25070
X10015 2 digital_ldo_top_VIA10 $T=174220 86500 0 0 $X=173750 $Y=86270
X10016 2 digital_ldo_top_VIA10 $T=174220 90580 0 0 $X=173750 $Y=90350
X10017 2 digital_ldo_top_VIA10 $T=174220 94660 0 0 $X=173750 $Y=94430
X10018 2 digital_ldo_top_VIA10 $T=174220 98740 0 0 $X=173750 $Y=98510
X10019 2 digital_ldo_top_VIA10 $T=174220 102820 0 0 $X=173750 $Y=102590
X10020 2 digital_ldo_top_VIA10 $T=174220 106900 0 0 $X=173750 $Y=106670
X10021 2 digital_ldo_top_VIA10 $T=174220 110980 0 0 $X=173750 $Y=110750
X10022 2 digital_ldo_top_VIA10 $T=174220 115060 0 0 $X=173750 $Y=114830
X10023 2 digital_ldo_top_VIA10 $T=174220 119140 0 0 $X=173750 $Y=118910
X10024 2 digital_ldo_top_VIA10 $T=174220 123220 0 0 $X=173750 $Y=122990
X10025 2 digital_ldo_top_VIA10 $T=174220 127300 0 0 $X=173750 $Y=127070
X10026 3 digital_ldo_top_VIA10 $T=177900 11700 0 0 $X=177430 $Y=11470
X10027 3 digital_ldo_top_VIA10 $T=177900 15780 0 0 $X=177430 $Y=15550
X10028 3 digital_ldo_top_VIA10 $T=177900 19860 0 0 $X=177430 $Y=19630
X10029 3 digital_ldo_top_VIA10 $T=177900 23940 0 0 $X=177430 $Y=23710
X10030 3 digital_ldo_top_VIA10 $T=177900 32100 0 0 $X=177430 $Y=31870
X10031 3 digital_ldo_top_VIA10 $T=177900 85140 0 0 $X=177430 $Y=84910
X10032 3 digital_ldo_top_VIA10 $T=177900 89220 0 0 $X=177430 $Y=88990
X10033 3 digital_ldo_top_VIA10 $T=177900 93300 0 0 $X=177430 $Y=93070
X10034 3 digital_ldo_top_VIA10 $T=177900 97380 0 0 $X=177430 $Y=97150
X10035 3 digital_ldo_top_VIA10 $T=177900 101460 0 0 $X=177430 $Y=101230
X10036 3 digital_ldo_top_VIA10 $T=177900 105540 0 0 $X=177430 $Y=105310
X10037 3 digital_ldo_top_VIA10 $T=177900 109620 0 0 $X=177430 $Y=109390
X10038 3 digital_ldo_top_VIA10 $T=177900 113700 0 0 $X=177430 $Y=113470
X10039 3 digital_ldo_top_VIA10 $T=177900 117780 0 0 $X=177430 $Y=117550
X10040 3 digital_ldo_top_VIA10 $T=177900 121860 0 0 $X=177430 $Y=121630
X10041 3 digital_ldo_top_VIA10 $T=177900 125940 0 0 $X=177430 $Y=125710
X10042 2 digital_ldo_top_VIA10 $T=179740 13060 0 0 $X=179270 $Y=12830
X10043 2 digital_ldo_top_VIA10 $T=179740 17140 0 0 $X=179270 $Y=16910
X10044 2 digital_ldo_top_VIA10 $T=179740 21220 0 0 $X=179270 $Y=20990
X10045 2 digital_ldo_top_VIA10 $T=179740 86500 0 0 $X=179270 $Y=86270
X10046 2 digital_ldo_top_VIA10 $T=179740 90580 0 0 $X=179270 $Y=90350
X10047 2 digital_ldo_top_VIA10 $T=179740 94660 0 0 $X=179270 $Y=94430
X10048 2 digital_ldo_top_VIA10 $T=179740 98740 0 0 $X=179270 $Y=98510
X10049 2 digital_ldo_top_VIA10 $T=179740 102820 0 0 $X=179270 $Y=102590
X10050 2 digital_ldo_top_VIA10 $T=179740 106900 0 0 $X=179270 $Y=106670
X10051 2 digital_ldo_top_VIA10 $T=179740 110980 0 0 $X=179270 $Y=110750
X10052 2 digital_ldo_top_VIA10 $T=179740 115060 0 0 $X=179270 $Y=114830
X10053 2 digital_ldo_top_VIA10 $T=179740 119140 0 0 $X=179270 $Y=118910
X10054 2 digital_ldo_top_VIA10 $T=179740 123220 0 0 $X=179270 $Y=122990
X10055 2 digital_ldo_top_VIA10 $T=179740 127300 0 0 $X=179270 $Y=127070
X10056 3 digital_ldo_top_VIA10 $T=183420 11700 0 0 $X=182950 $Y=11470
X10057 3 digital_ldo_top_VIA10 $T=183420 15780 0 0 $X=182950 $Y=15550
X10058 3 digital_ldo_top_VIA10 $T=183420 19860 0 0 $X=182950 $Y=19630
X10059 3 digital_ldo_top_VIA10 $T=183420 23940 0 0 $X=182950 $Y=23710
X10060 3 digital_ldo_top_VIA10 $T=183420 32100 0 0 $X=182950 $Y=31870
X10061 3 digital_ldo_top_VIA10 $T=183420 85140 0 0 $X=182950 $Y=84910
X10062 3 digital_ldo_top_VIA10 $T=183420 89220 0 0 $X=182950 $Y=88990
X10063 3 digital_ldo_top_VIA10 $T=183420 93300 0 0 $X=182950 $Y=93070
X10064 3 digital_ldo_top_VIA10 $T=183420 97380 0 0 $X=182950 $Y=97150
X10065 3 digital_ldo_top_VIA10 $T=183420 101460 0 0 $X=182950 $Y=101230
X10066 3 digital_ldo_top_VIA10 $T=183420 105540 0 0 $X=182950 $Y=105310
X10067 3 digital_ldo_top_VIA10 $T=183420 109620 0 0 $X=182950 $Y=109390
X10068 3 digital_ldo_top_VIA10 $T=183420 113700 0 0 $X=182950 $Y=113470
X10069 3 digital_ldo_top_VIA10 $T=183420 117780 0 0 $X=182950 $Y=117550
X10070 3 digital_ldo_top_VIA10 $T=183420 121860 0 0 $X=182950 $Y=121630
X10071 3 digital_ldo_top_VIA10 $T=183420 125940 0 0 $X=182950 $Y=125710
X10072 2 digital_ldo_top_VIA10 $T=185260 13060 0 0 $X=184790 $Y=12830
X10073 2 digital_ldo_top_VIA10 $T=185260 17140 0 0 $X=184790 $Y=16910
X10074 2 digital_ldo_top_VIA10 $T=185260 21220 0 0 $X=184790 $Y=20990
X10075 2 digital_ldo_top_VIA10 $T=185260 25300 0 0 $X=184790 $Y=25070
X10076 2 digital_ldo_top_VIA10 $T=185260 86500 0 0 $X=184790 $Y=86270
X10077 2 digital_ldo_top_VIA10 $T=185260 90580 0 0 $X=184790 $Y=90350
X10078 2 digital_ldo_top_VIA10 $T=185260 94660 0 0 $X=184790 $Y=94430
X10079 2 digital_ldo_top_VIA10 $T=185260 98740 0 0 $X=184790 $Y=98510
X10080 2 digital_ldo_top_VIA10 $T=185260 102820 0 0 $X=184790 $Y=102590
X10081 2 digital_ldo_top_VIA10 $T=185260 106900 0 0 $X=184790 $Y=106670
X10082 2 digital_ldo_top_VIA10 $T=185260 110980 0 0 $X=184790 $Y=110750
X10083 2 digital_ldo_top_VIA10 $T=185260 115060 0 0 $X=184790 $Y=114830
X10084 2 digital_ldo_top_VIA10 $T=185260 119140 0 0 $X=184790 $Y=118910
X10085 2 digital_ldo_top_VIA10 $T=185260 123220 0 0 $X=184790 $Y=122990
X10086 2 digital_ldo_top_VIA10 $T=185260 127300 0 0 $X=184790 $Y=127070
X10087 3 digital_ldo_top_VIA10 $T=188940 11700 0 0 $X=188470 $Y=11470
X10088 3 digital_ldo_top_VIA10 $T=188940 15780 0 0 $X=188470 $Y=15550
X10089 3 digital_ldo_top_VIA10 $T=188940 19860 0 0 $X=188470 $Y=19630
X10090 3 digital_ldo_top_VIA10 $T=188940 23940 0 0 $X=188470 $Y=23710
X10091 3 digital_ldo_top_VIA10 $T=188940 32100 0 0 $X=188470 $Y=31870
X10092 3 digital_ldo_top_VIA10 $T=188940 85140 0 0 $X=188470 $Y=84910
X10093 3 digital_ldo_top_VIA10 $T=188940 89220 0 0 $X=188470 $Y=88990
X10094 3 digital_ldo_top_VIA10 $T=188940 93300 0 0 $X=188470 $Y=93070
X10095 3 digital_ldo_top_VIA10 $T=188940 97380 0 0 $X=188470 $Y=97150
X10096 3 digital_ldo_top_VIA10 $T=188940 101460 0 0 $X=188470 $Y=101230
X10097 3 digital_ldo_top_VIA10 $T=188940 105540 0 0 $X=188470 $Y=105310
X10098 3 digital_ldo_top_VIA10 $T=188940 109620 0 0 $X=188470 $Y=109390
X10099 3 digital_ldo_top_VIA10 $T=188940 113700 0 0 $X=188470 $Y=113470
X10100 3 digital_ldo_top_VIA10 $T=188940 117780 0 0 $X=188470 $Y=117550
X10101 3 digital_ldo_top_VIA10 $T=188940 121860 0 0 $X=188470 $Y=121630
X10102 3 digital_ldo_top_VIA10 $T=188940 125940 0 0 $X=188470 $Y=125710
X10103 2 digital_ldo_top_VIA10 $T=190780 13060 0 0 $X=190310 $Y=12830
X10104 2 digital_ldo_top_VIA10 $T=190780 17140 0 0 $X=190310 $Y=16910
X10105 2 digital_ldo_top_VIA10 $T=190780 21220 0 0 $X=190310 $Y=20990
X10106 2 digital_ldo_top_VIA10 $T=190780 25300 0 0 $X=190310 $Y=25070
X10107 2 digital_ldo_top_VIA10 $T=190780 86500 0 0 $X=190310 $Y=86270
X10108 2 digital_ldo_top_VIA10 $T=190780 90580 0 0 $X=190310 $Y=90350
X10109 2 digital_ldo_top_VIA10 $T=190780 94660 0 0 $X=190310 $Y=94430
X10110 2 digital_ldo_top_VIA10 $T=190780 98740 0 0 $X=190310 $Y=98510
X10111 2 digital_ldo_top_VIA10 $T=190780 102820 0 0 $X=190310 $Y=102590
X10112 2 digital_ldo_top_VIA10 $T=190780 106900 0 0 $X=190310 $Y=106670
X10113 2 digital_ldo_top_VIA10 $T=190780 110980 0 0 $X=190310 $Y=110750
X10114 2 digital_ldo_top_VIA10 $T=190780 115060 0 0 $X=190310 $Y=114830
X10115 2 digital_ldo_top_VIA10 $T=190780 119140 0 0 $X=190310 $Y=118910
X10116 2 digital_ldo_top_VIA10 $T=190780 123220 0 0 $X=190310 $Y=122990
X10117 2 digital_ldo_top_VIA10 $T=190780 127300 0 0 $X=190310 $Y=127070
X10118 3 digital_ldo_top_VIA10 $T=194460 11700 0 0 $X=193990 $Y=11470
X10119 3 digital_ldo_top_VIA10 $T=194460 15780 0 0 $X=193990 $Y=15550
X10120 3 digital_ldo_top_VIA10 $T=194460 19860 0 0 $X=193990 $Y=19630
X10121 3 digital_ldo_top_VIA10 $T=194460 23940 0 0 $X=193990 $Y=23710
X10122 3 digital_ldo_top_VIA10 $T=194460 32100 0 0 $X=193990 $Y=31870
X10123 3 digital_ldo_top_VIA10 $T=194460 85140 0 0 $X=193990 $Y=84910
X10124 3 digital_ldo_top_VIA10 $T=194460 89220 0 0 $X=193990 $Y=88990
X10125 3 digital_ldo_top_VIA10 $T=194460 93300 0 0 $X=193990 $Y=93070
X10126 3 digital_ldo_top_VIA10 $T=194460 97380 0 0 $X=193990 $Y=97150
X10127 3 digital_ldo_top_VIA10 $T=194460 101460 0 0 $X=193990 $Y=101230
X10128 3 digital_ldo_top_VIA10 $T=194460 105540 0 0 $X=193990 $Y=105310
X10129 3 digital_ldo_top_VIA10 $T=194460 109620 0 0 $X=193990 $Y=109390
X10130 3 digital_ldo_top_VIA10 $T=194460 113700 0 0 $X=193990 $Y=113470
X10131 3 digital_ldo_top_VIA10 $T=194460 117780 0 0 $X=193990 $Y=117550
X10132 3 digital_ldo_top_VIA10 $T=194460 121860 0 0 $X=193990 $Y=121630
X10133 3 digital_ldo_top_VIA10 $T=194460 125940 0 0 $X=193990 $Y=125710
X10134 2 digital_ldo_top_VIA10 $T=196300 13060 0 0 $X=195830 $Y=12830
X10135 2 digital_ldo_top_VIA10 $T=196300 17140 0 0 $X=195830 $Y=16910
X10136 2 digital_ldo_top_VIA10 $T=196300 21220 0 0 $X=195830 $Y=20990
X10137 2 digital_ldo_top_VIA10 $T=196300 25300 0 0 $X=195830 $Y=25070
X10138 2 digital_ldo_top_VIA10 $T=196300 86500 0 0 $X=195830 $Y=86270
X10139 2 digital_ldo_top_VIA10 $T=196300 90580 0 0 $X=195830 $Y=90350
X10140 2 digital_ldo_top_VIA10 $T=196300 94660 0 0 $X=195830 $Y=94430
X10141 2 digital_ldo_top_VIA10 $T=196300 98740 0 0 $X=195830 $Y=98510
X10142 2 digital_ldo_top_VIA10 $T=196300 102820 0 0 $X=195830 $Y=102590
X10143 2 digital_ldo_top_VIA10 $T=196300 106900 0 0 $X=195830 $Y=106670
X10144 2 digital_ldo_top_VIA10 $T=196300 110980 0 0 $X=195830 $Y=110750
X10145 2 digital_ldo_top_VIA10 $T=196300 115060 0 0 $X=195830 $Y=114830
X10146 2 digital_ldo_top_VIA10 $T=196300 119140 0 0 $X=195830 $Y=118910
X10147 2 digital_ldo_top_VIA10 $T=196300 123220 0 0 $X=195830 $Y=122990
X10148 2 digital_ldo_top_VIA10 $T=196300 127300 0 0 $X=195830 $Y=127070
X10149 3 digital_ldo_top_VIA10 $T=199980 11700 0 0 $X=199510 $Y=11470
X10150 3 digital_ldo_top_VIA10 $T=199980 15780 0 0 $X=199510 $Y=15550
X10151 3 digital_ldo_top_VIA10 $T=199980 19860 0 0 $X=199510 $Y=19630
X10152 3 digital_ldo_top_VIA10 $T=199980 23940 0 0 $X=199510 $Y=23710
X10153 3 digital_ldo_top_VIA10 $T=199980 32100 0 0 $X=199510 $Y=31870
X10154 3 digital_ldo_top_VIA10 $T=199980 85140 0 0 $X=199510 $Y=84910
X10155 3 digital_ldo_top_VIA10 $T=199980 89220 0 0 $X=199510 $Y=88990
X10156 3 digital_ldo_top_VIA10 $T=199980 93300 0 0 $X=199510 $Y=93070
X10157 3 digital_ldo_top_VIA10 $T=199980 97380 0 0 $X=199510 $Y=97150
X10158 3 digital_ldo_top_VIA10 $T=199980 101460 0 0 $X=199510 $Y=101230
X10159 3 digital_ldo_top_VIA10 $T=199980 105540 0 0 $X=199510 $Y=105310
X10160 3 digital_ldo_top_VIA10 $T=199980 109620 0 0 $X=199510 $Y=109390
X10161 3 digital_ldo_top_VIA10 $T=199980 113700 0 0 $X=199510 $Y=113470
X10162 3 digital_ldo_top_VIA10 $T=199980 117780 0 0 $X=199510 $Y=117550
X10163 3 digital_ldo_top_VIA10 $T=199980 121860 0 0 $X=199510 $Y=121630
X10164 3 digital_ldo_top_VIA10 $T=199980 125940 0 0 $X=199510 $Y=125710
X10165 2 digital_ldo_top_VIA10 $T=201820 13060 0 0 $X=201350 $Y=12830
X10166 2 digital_ldo_top_VIA10 $T=201820 17140 0 0 $X=201350 $Y=16910
X10167 2 digital_ldo_top_VIA10 $T=201820 21220 0 0 $X=201350 $Y=20990
X10168 2 digital_ldo_top_VIA10 $T=201820 25300 0 0 $X=201350 $Y=25070
X10169 2 digital_ldo_top_VIA10 $T=201820 86500 0 0 $X=201350 $Y=86270
X10170 2 digital_ldo_top_VIA10 $T=201820 90580 0 0 $X=201350 $Y=90350
X10171 2 digital_ldo_top_VIA10 $T=201820 94660 0 0 $X=201350 $Y=94430
X10172 2 digital_ldo_top_VIA10 $T=201820 98740 0 0 $X=201350 $Y=98510
X10173 2 digital_ldo_top_VIA10 $T=201820 102820 0 0 $X=201350 $Y=102590
X10174 2 digital_ldo_top_VIA10 $T=201820 106900 0 0 $X=201350 $Y=106670
X10175 2 digital_ldo_top_VIA10 $T=201820 110980 0 0 $X=201350 $Y=110750
X10176 2 digital_ldo_top_VIA10 $T=201820 115060 0 0 $X=201350 $Y=114830
X10177 2 digital_ldo_top_VIA10 $T=201820 119140 0 0 $X=201350 $Y=118910
X10178 2 digital_ldo_top_VIA10 $T=201820 123220 0 0 $X=201350 $Y=122990
X10179 2 digital_ldo_top_VIA10 $T=201820 127300 0 0 $X=201350 $Y=127070
X10180 3 digital_ldo_top_VIA10 $T=205500 11700 0 0 $X=205030 $Y=11470
X10181 3 digital_ldo_top_VIA10 $T=205500 15780 0 0 $X=205030 $Y=15550
X10182 3 digital_ldo_top_VIA10 $T=205500 19860 0 0 $X=205030 $Y=19630
X10183 3 digital_ldo_top_VIA10 $T=205500 32100 0 0 $X=205030 $Y=31870
X10184 3 digital_ldo_top_VIA10 $T=205500 85140 0 0 $X=205030 $Y=84910
X10185 3 digital_ldo_top_VIA10 $T=205500 89220 0 0 $X=205030 $Y=88990
X10186 3 digital_ldo_top_VIA10 $T=205500 93300 0 0 $X=205030 $Y=93070
X10187 3 digital_ldo_top_VIA10 $T=205500 97380 0 0 $X=205030 $Y=97150
X10188 3 digital_ldo_top_VIA10 $T=205500 101460 0 0 $X=205030 $Y=101230
X10189 3 digital_ldo_top_VIA10 $T=205500 105540 0 0 $X=205030 $Y=105310
X10190 3 digital_ldo_top_VIA10 $T=205500 109620 0 0 $X=205030 $Y=109390
X10191 3 digital_ldo_top_VIA10 $T=205500 113700 0 0 $X=205030 $Y=113470
X10192 3 digital_ldo_top_VIA10 $T=205500 117780 0 0 $X=205030 $Y=117550
X10193 3 digital_ldo_top_VIA10 $T=205500 121860 0 0 $X=205030 $Y=121630
X10194 3 digital_ldo_top_VIA10 $T=205500 125940 0 0 $X=205030 $Y=125710
X10195 2 digital_ldo_top_VIA10 $T=207340 13060 0 0 $X=206870 $Y=12830
X10196 2 digital_ldo_top_VIA10 $T=207340 17140 0 0 $X=206870 $Y=16910
X10197 2 digital_ldo_top_VIA10 $T=207340 21220 0 0 $X=206870 $Y=20990
X10198 2 digital_ldo_top_VIA10 $T=207340 25300 0 0 $X=206870 $Y=25070
X10199 2 digital_ldo_top_VIA10 $T=207340 86500 0 0 $X=206870 $Y=86270
X10200 2 digital_ldo_top_VIA10 $T=207340 90580 0 0 $X=206870 $Y=90350
X10201 2 digital_ldo_top_VIA10 $T=207340 94660 0 0 $X=206870 $Y=94430
X10202 2 digital_ldo_top_VIA10 $T=207340 98740 0 0 $X=206870 $Y=98510
X10203 2 digital_ldo_top_VIA10 $T=207340 102820 0 0 $X=206870 $Y=102590
X10204 2 digital_ldo_top_VIA10 $T=207340 106900 0 0 $X=206870 $Y=106670
X10205 2 digital_ldo_top_VIA10 $T=207340 110980 0 0 $X=206870 $Y=110750
X10206 2 digital_ldo_top_VIA10 $T=207340 115060 0 0 $X=206870 $Y=114830
X10207 2 digital_ldo_top_VIA10 $T=207340 119140 0 0 $X=206870 $Y=118910
X10208 2 digital_ldo_top_VIA10 $T=207340 123220 0 0 $X=206870 $Y=122990
X10209 2 digital_ldo_top_VIA10 $T=207340 127300 0 0 $X=206870 $Y=127070
X10210 3 digital_ldo_top_VIA10 $T=211020 11700 0 0 $X=210550 $Y=11470
X10211 3 digital_ldo_top_VIA10 $T=211020 15780 0 0 $X=210550 $Y=15550
X10212 3 digital_ldo_top_VIA10 $T=211020 19860 0 0 $X=210550 $Y=19630
X10213 3 digital_ldo_top_VIA10 $T=211020 23940 0 0 $X=210550 $Y=23710
X10214 3 digital_ldo_top_VIA10 $T=211020 32100 0 0 $X=210550 $Y=31870
X10215 3 digital_ldo_top_VIA10 $T=211020 85140 0 0 $X=210550 $Y=84910
X10216 3 digital_ldo_top_VIA10 $T=211020 89220 0 0 $X=210550 $Y=88990
X10217 3 digital_ldo_top_VIA10 $T=211020 93300 0 0 $X=210550 $Y=93070
X10218 3 digital_ldo_top_VIA10 $T=211020 97380 0 0 $X=210550 $Y=97150
X10219 3 digital_ldo_top_VIA10 $T=211020 101460 0 0 $X=210550 $Y=101230
X10220 3 digital_ldo_top_VIA10 $T=211020 105540 0 0 $X=210550 $Y=105310
X10221 3 digital_ldo_top_VIA10 $T=211020 109620 0 0 $X=210550 $Y=109390
X10222 3 digital_ldo_top_VIA10 $T=211020 113700 0 0 $X=210550 $Y=113470
X10223 3 digital_ldo_top_VIA10 $T=211020 117780 0 0 $X=210550 $Y=117550
X10224 3 digital_ldo_top_VIA10 $T=211020 121860 0 0 $X=210550 $Y=121630
X10225 3 digital_ldo_top_VIA10 $T=211020 125940 0 0 $X=210550 $Y=125710
X10226 2 digital_ldo_top_VIA10 $T=212860 13060 0 0 $X=212390 $Y=12830
X10227 2 digital_ldo_top_VIA10 $T=212860 17140 0 0 $X=212390 $Y=16910
X10228 2 digital_ldo_top_VIA10 $T=212860 21220 0 0 $X=212390 $Y=20990
X10229 2 digital_ldo_top_VIA10 $T=212860 25300 0 0 $X=212390 $Y=25070
X10230 2 digital_ldo_top_VIA10 $T=212860 86500 0 0 $X=212390 $Y=86270
X10231 2 digital_ldo_top_VIA10 $T=212860 90580 0 0 $X=212390 $Y=90350
X10232 2 digital_ldo_top_VIA10 $T=212860 94660 0 0 $X=212390 $Y=94430
X10233 2 digital_ldo_top_VIA10 $T=212860 98740 0 0 $X=212390 $Y=98510
X10234 2 digital_ldo_top_VIA10 $T=212860 102820 0 0 $X=212390 $Y=102590
X10235 2 digital_ldo_top_VIA10 $T=212860 106900 0 0 $X=212390 $Y=106670
X10236 2 digital_ldo_top_VIA10 $T=212860 110980 0 0 $X=212390 $Y=110750
X10237 2 digital_ldo_top_VIA10 $T=212860 115060 0 0 $X=212390 $Y=114830
X10238 2 digital_ldo_top_VIA10 $T=212860 119140 0 0 $X=212390 $Y=118910
X10239 2 digital_ldo_top_VIA10 $T=212860 123220 0 0 $X=212390 $Y=122990
X10240 2 digital_ldo_top_VIA10 $T=212860 127300 0 0 $X=212390 $Y=127070
X10241 3 digital_ldo_top_VIA10 $T=216540 11700 0 0 $X=216070 $Y=11470
X10242 3 digital_ldo_top_VIA10 $T=216540 15780 0 0 $X=216070 $Y=15550
X10243 3 digital_ldo_top_VIA10 $T=216540 19860 0 0 $X=216070 $Y=19630
X10244 3 digital_ldo_top_VIA10 $T=216540 23940 0 0 $X=216070 $Y=23710
X10245 3 digital_ldo_top_VIA10 $T=216540 32100 0 0 $X=216070 $Y=31870
X10246 3 digital_ldo_top_VIA10 $T=216540 85140 0 0 $X=216070 $Y=84910
X10247 3 digital_ldo_top_VIA10 $T=216540 89220 0 0 $X=216070 $Y=88990
X10248 3 digital_ldo_top_VIA10 $T=216540 93300 0 0 $X=216070 $Y=93070
X10249 3 digital_ldo_top_VIA10 $T=216540 97380 0 0 $X=216070 $Y=97150
X10250 3 digital_ldo_top_VIA10 $T=216540 101460 0 0 $X=216070 $Y=101230
X10251 3 digital_ldo_top_VIA10 $T=216540 105540 0 0 $X=216070 $Y=105310
X10252 3 digital_ldo_top_VIA10 $T=216540 109620 0 0 $X=216070 $Y=109390
X10253 3 digital_ldo_top_VIA10 $T=216540 113700 0 0 $X=216070 $Y=113470
X10254 3 digital_ldo_top_VIA10 $T=216540 117780 0 0 $X=216070 $Y=117550
X10255 3 digital_ldo_top_VIA10 $T=216540 121860 0 0 $X=216070 $Y=121630
X10256 3 digital_ldo_top_VIA10 $T=216540 125940 0 0 $X=216070 $Y=125710
X10257 2 digital_ldo_top_VIA10 $T=218380 13060 0 0 $X=217910 $Y=12830
X10258 2 digital_ldo_top_VIA10 $T=218380 17140 0 0 $X=217910 $Y=16910
X10259 2 digital_ldo_top_VIA10 $T=218380 21220 0 0 $X=217910 $Y=20990
X10260 2 digital_ldo_top_VIA10 $T=218380 86500 0 0 $X=217910 $Y=86270
X10261 2 digital_ldo_top_VIA10 $T=218380 90580 0 0 $X=217910 $Y=90350
X10262 2 digital_ldo_top_VIA10 $T=218380 94660 0 0 $X=217910 $Y=94430
X10263 2 digital_ldo_top_VIA10 $T=218380 98740 0 0 $X=217910 $Y=98510
X10264 2 digital_ldo_top_VIA10 $T=218380 102820 0 0 $X=217910 $Y=102590
X10265 2 digital_ldo_top_VIA10 $T=218380 106900 0 0 $X=217910 $Y=106670
X10266 2 digital_ldo_top_VIA10 $T=218380 110980 0 0 $X=217910 $Y=110750
X10267 2 digital_ldo_top_VIA10 $T=218380 115060 0 0 $X=217910 $Y=114830
X10268 2 digital_ldo_top_VIA10 $T=218380 119140 0 0 $X=217910 $Y=118910
X10269 2 digital_ldo_top_VIA10 $T=218380 123220 0 0 $X=217910 $Y=122990
X10270 2 digital_ldo_top_VIA10 $T=218380 127300 0 0 $X=217910 $Y=127070
X10271 3 digital_ldo_top_VIA10 $T=222060 11700 0 0 $X=221590 $Y=11470
X10272 3 digital_ldo_top_VIA10 $T=222060 15780 0 0 $X=221590 $Y=15550
X10273 3 digital_ldo_top_VIA10 $T=222060 19860 0 0 $X=221590 $Y=19630
X10274 3 digital_ldo_top_VIA10 $T=222060 23940 0 0 $X=221590 $Y=23710
X10275 3 digital_ldo_top_VIA10 $T=222060 32100 0 0 $X=221590 $Y=31870
X10276 3 digital_ldo_top_VIA10 $T=222060 85140 0 0 $X=221590 $Y=84910
X10277 3 digital_ldo_top_VIA10 $T=222060 89220 0 0 $X=221590 $Y=88990
X10278 3 digital_ldo_top_VIA10 $T=222060 93300 0 0 $X=221590 $Y=93070
X10279 3 digital_ldo_top_VIA10 $T=222060 97380 0 0 $X=221590 $Y=97150
X10280 3 digital_ldo_top_VIA10 $T=222060 101460 0 0 $X=221590 $Y=101230
X10281 3 digital_ldo_top_VIA10 $T=222060 105540 0 0 $X=221590 $Y=105310
X10282 3 digital_ldo_top_VIA10 $T=222060 109620 0 0 $X=221590 $Y=109390
X10283 3 digital_ldo_top_VIA10 $T=222060 113700 0 0 $X=221590 $Y=113470
X10284 3 digital_ldo_top_VIA10 $T=222060 117780 0 0 $X=221590 $Y=117550
X10285 3 digital_ldo_top_VIA10 $T=222060 121860 0 0 $X=221590 $Y=121630
X10286 3 digital_ldo_top_VIA10 $T=222060 125940 0 0 $X=221590 $Y=125710
X10287 2 digital_ldo_top_VIA10 $T=223900 13060 0 0 $X=223430 $Y=12830
X10288 2 digital_ldo_top_VIA10 $T=223900 17140 0 0 $X=223430 $Y=16910
X10289 2 digital_ldo_top_VIA10 $T=223900 21220 0 0 $X=223430 $Y=20990
X10290 2 digital_ldo_top_VIA10 $T=223900 25300 0 0 $X=223430 $Y=25070
X10291 2 digital_ldo_top_VIA10 $T=223900 86500 0 0 $X=223430 $Y=86270
X10292 2 digital_ldo_top_VIA10 $T=223900 90580 0 0 $X=223430 $Y=90350
X10293 2 digital_ldo_top_VIA10 $T=223900 94660 0 0 $X=223430 $Y=94430
X10294 2 digital_ldo_top_VIA10 $T=223900 98740 0 0 $X=223430 $Y=98510
X10295 2 digital_ldo_top_VIA10 $T=223900 102820 0 0 $X=223430 $Y=102590
X10296 2 digital_ldo_top_VIA10 $T=223900 106900 0 0 $X=223430 $Y=106670
X10297 2 digital_ldo_top_VIA10 $T=223900 110980 0 0 $X=223430 $Y=110750
X10298 2 digital_ldo_top_VIA10 $T=223900 115060 0 0 $X=223430 $Y=114830
X10299 2 digital_ldo_top_VIA10 $T=223900 119140 0 0 $X=223430 $Y=118910
X10300 2 digital_ldo_top_VIA10 $T=223900 123220 0 0 $X=223430 $Y=122990
X10301 2 digital_ldo_top_VIA10 $T=223900 127300 0 0 $X=223430 $Y=127070
X10302 3 digital_ldo_top_VIA10 $T=227580 11700 0 0 $X=227110 $Y=11470
X10303 3 digital_ldo_top_VIA10 $T=227580 15780 0 0 $X=227110 $Y=15550
X10304 3 digital_ldo_top_VIA10 $T=227580 19860 0 0 $X=227110 $Y=19630
X10305 3 digital_ldo_top_VIA10 $T=227580 23940 0 0 $X=227110 $Y=23710
X10306 3 digital_ldo_top_VIA10 $T=227580 32100 0 0 $X=227110 $Y=31870
X10307 3 digital_ldo_top_VIA10 $T=227580 85140 0 0 $X=227110 $Y=84910
X10308 3 digital_ldo_top_VIA10 $T=227580 89220 0 0 $X=227110 $Y=88990
X10309 3 digital_ldo_top_VIA10 $T=227580 93300 0 0 $X=227110 $Y=93070
X10310 3 digital_ldo_top_VIA10 $T=227580 97380 0 0 $X=227110 $Y=97150
X10311 3 digital_ldo_top_VIA10 $T=227580 101460 0 0 $X=227110 $Y=101230
X10312 3 digital_ldo_top_VIA10 $T=227580 105540 0 0 $X=227110 $Y=105310
X10313 3 digital_ldo_top_VIA10 $T=227580 109620 0 0 $X=227110 $Y=109390
X10314 3 digital_ldo_top_VIA10 $T=227580 113700 0 0 $X=227110 $Y=113470
X10315 3 digital_ldo_top_VIA10 $T=227580 117780 0 0 $X=227110 $Y=117550
X10316 3 digital_ldo_top_VIA10 $T=227580 121860 0 0 $X=227110 $Y=121630
X10317 3 digital_ldo_top_VIA10 $T=227580 125940 0 0 $X=227110 $Y=125710
X10318 2 digital_ldo_top_VIA10 $T=229420 13060 0 0 $X=228950 $Y=12830
X10319 2 digital_ldo_top_VIA10 $T=229420 17140 0 0 $X=228950 $Y=16910
X10320 2 digital_ldo_top_VIA10 $T=229420 21220 0 0 $X=228950 $Y=20990
X10321 2 digital_ldo_top_VIA10 $T=229420 25300 0 0 $X=228950 $Y=25070
X10322 2 digital_ldo_top_VIA10 $T=229420 86500 0 0 $X=228950 $Y=86270
X10323 2 digital_ldo_top_VIA10 $T=229420 90580 0 0 $X=228950 $Y=90350
X10324 2 digital_ldo_top_VIA10 $T=229420 94660 0 0 $X=228950 $Y=94430
X10325 2 digital_ldo_top_VIA10 $T=229420 98740 0 0 $X=228950 $Y=98510
X10326 2 digital_ldo_top_VIA10 $T=229420 102820 0 0 $X=228950 $Y=102590
X10327 2 digital_ldo_top_VIA10 $T=229420 106900 0 0 $X=228950 $Y=106670
X10328 2 digital_ldo_top_VIA10 $T=229420 110980 0 0 $X=228950 $Y=110750
X10329 2 digital_ldo_top_VIA10 $T=229420 115060 0 0 $X=228950 $Y=114830
X10330 2 digital_ldo_top_VIA10 $T=229420 119140 0 0 $X=228950 $Y=118910
X10331 2 digital_ldo_top_VIA10 $T=229420 123220 0 0 $X=228950 $Y=122990
X10332 2 digital_ldo_top_VIA10 $T=229420 127300 0 0 $X=228950 $Y=127070
X10333 3 digital_ldo_top_VIA10 $T=233100 11700 0 0 $X=232630 $Y=11470
X10334 3 digital_ldo_top_VIA10 $T=233100 15780 0 0 $X=232630 $Y=15550
X10335 3 digital_ldo_top_VIA10 $T=233100 19860 0 0 $X=232630 $Y=19630
X10336 3 digital_ldo_top_VIA10 $T=233100 23940 0 0 $X=232630 $Y=23710
X10337 3 digital_ldo_top_VIA10 $T=233100 32100 0 0 $X=232630 $Y=31870
X10338 3 digital_ldo_top_VIA10 $T=233100 85140 0 0 $X=232630 $Y=84910
X10339 3 digital_ldo_top_VIA10 $T=233100 89220 0 0 $X=232630 $Y=88990
X10340 3 digital_ldo_top_VIA10 $T=233100 93300 0 0 $X=232630 $Y=93070
X10341 3 digital_ldo_top_VIA10 $T=233100 97380 0 0 $X=232630 $Y=97150
X10342 3 digital_ldo_top_VIA10 $T=233100 101460 0 0 $X=232630 $Y=101230
X10343 3 digital_ldo_top_VIA10 $T=233100 105540 0 0 $X=232630 $Y=105310
X10344 3 digital_ldo_top_VIA10 $T=233100 109620 0 0 $X=232630 $Y=109390
X10345 3 digital_ldo_top_VIA10 $T=233100 113700 0 0 $X=232630 $Y=113470
X10346 3 digital_ldo_top_VIA10 $T=233100 117780 0 0 $X=232630 $Y=117550
X10347 3 digital_ldo_top_VIA10 $T=233100 121860 0 0 $X=232630 $Y=121630
X10348 3 digital_ldo_top_VIA10 $T=233100 125940 0 0 $X=232630 $Y=125710
X10349 2 digital_ldo_top_VIA10 $T=234940 13060 0 0 $X=234470 $Y=12830
X10350 2 digital_ldo_top_VIA10 $T=234940 17140 0 0 $X=234470 $Y=16910
X10351 2 digital_ldo_top_VIA10 $T=234940 21220 0 0 $X=234470 $Y=20990
X10352 2 digital_ldo_top_VIA10 $T=234940 25300 0 0 $X=234470 $Y=25070
X10353 2 digital_ldo_top_VIA10 $T=234940 86500 0 0 $X=234470 $Y=86270
X10354 2 digital_ldo_top_VIA10 $T=234940 90580 0 0 $X=234470 $Y=90350
X10355 2 digital_ldo_top_VIA10 $T=234940 94660 0 0 $X=234470 $Y=94430
X10356 2 digital_ldo_top_VIA10 $T=234940 98740 0 0 $X=234470 $Y=98510
X10357 2 digital_ldo_top_VIA10 $T=234940 102820 0 0 $X=234470 $Y=102590
X10358 2 digital_ldo_top_VIA10 $T=234940 106900 0 0 $X=234470 $Y=106670
X10359 2 digital_ldo_top_VIA10 $T=234940 110980 0 0 $X=234470 $Y=110750
X10360 2 digital_ldo_top_VIA10 $T=234940 115060 0 0 $X=234470 $Y=114830
X10361 2 digital_ldo_top_VIA10 $T=234940 119140 0 0 $X=234470 $Y=118910
X10362 2 digital_ldo_top_VIA10 $T=234940 123220 0 0 $X=234470 $Y=122990
X10363 2 digital_ldo_top_VIA10 $T=234940 127300 0 0 $X=234470 $Y=127070
X10364 3 digital_ldo_top_VIA10 $T=238620 11700 0 0 $X=238150 $Y=11470
X10365 3 digital_ldo_top_VIA10 $T=238620 15780 0 0 $X=238150 $Y=15550
X10366 3 digital_ldo_top_VIA10 $T=238620 19860 0 0 $X=238150 $Y=19630
X10367 3 digital_ldo_top_VIA10 $T=238620 23940 0 0 $X=238150 $Y=23710
X10368 3 digital_ldo_top_VIA10 $T=238620 32100 0 0 $X=238150 $Y=31870
X10369 3 digital_ldo_top_VIA10 $T=238620 85140 0 0 $X=238150 $Y=84910
X10370 3 digital_ldo_top_VIA10 $T=238620 89220 0 0 $X=238150 $Y=88990
X10371 3 digital_ldo_top_VIA10 $T=238620 93300 0 0 $X=238150 $Y=93070
X10372 3 digital_ldo_top_VIA10 $T=238620 97380 0 0 $X=238150 $Y=97150
X10373 3 digital_ldo_top_VIA10 $T=238620 101460 0 0 $X=238150 $Y=101230
X10374 3 digital_ldo_top_VIA10 $T=238620 105540 0 0 $X=238150 $Y=105310
X10375 3 digital_ldo_top_VIA10 $T=238620 109620 0 0 $X=238150 $Y=109390
X10376 3 digital_ldo_top_VIA10 $T=238620 113700 0 0 $X=238150 $Y=113470
X10377 3 digital_ldo_top_VIA10 $T=238620 117780 0 0 $X=238150 $Y=117550
X10378 3 digital_ldo_top_VIA10 $T=238620 121860 0 0 $X=238150 $Y=121630
X10379 3 digital_ldo_top_VIA10 $T=238620 125940 0 0 $X=238150 $Y=125710
X10380 2 digital_ldo_top_VIA10 $T=240460 13060 0 0 $X=239990 $Y=12830
X10381 2 digital_ldo_top_VIA10 $T=240460 17140 0 0 $X=239990 $Y=16910
X10382 2 digital_ldo_top_VIA10 $T=240460 21220 0 0 $X=239990 $Y=20990
X10383 2 digital_ldo_top_VIA10 $T=240460 25300 0 0 $X=239990 $Y=25070
X10384 2 digital_ldo_top_VIA10 $T=240460 86500 0 0 $X=239990 $Y=86270
X10385 2 digital_ldo_top_VIA10 $T=240460 90580 0 0 $X=239990 $Y=90350
X10386 2 digital_ldo_top_VIA10 $T=240460 94660 0 0 $X=239990 $Y=94430
X10387 2 digital_ldo_top_VIA10 $T=240460 98740 0 0 $X=239990 $Y=98510
X10388 2 digital_ldo_top_VIA10 $T=240460 102820 0 0 $X=239990 $Y=102590
X10389 2 digital_ldo_top_VIA10 $T=240460 106900 0 0 $X=239990 $Y=106670
X10390 2 digital_ldo_top_VIA10 $T=240460 110980 0 0 $X=239990 $Y=110750
X10391 2 digital_ldo_top_VIA10 $T=240460 115060 0 0 $X=239990 $Y=114830
X10392 2 digital_ldo_top_VIA10 $T=240460 119140 0 0 $X=239990 $Y=118910
X10393 2 digital_ldo_top_VIA10 $T=240460 123220 0 0 $X=239990 $Y=122990
X10394 2 digital_ldo_top_VIA10 $T=240460 127300 0 0 $X=239990 $Y=127070
X10395 3 digital_ldo_top_VIA10 $T=244140 11700 0 0 $X=243670 $Y=11470
X10396 3 digital_ldo_top_VIA10 $T=244140 15780 0 0 $X=243670 $Y=15550
X10397 3 digital_ldo_top_VIA10 $T=244140 19860 0 0 $X=243670 $Y=19630
X10398 3 digital_ldo_top_VIA10 $T=244140 32100 0 0 $X=243670 $Y=31870
X10399 3 digital_ldo_top_VIA10 $T=244140 85140 0 0 $X=243670 $Y=84910
X10400 3 digital_ldo_top_VIA10 $T=244140 89220 0 0 $X=243670 $Y=88990
X10401 3 digital_ldo_top_VIA10 $T=244140 93300 0 0 $X=243670 $Y=93070
X10402 3 digital_ldo_top_VIA10 $T=244140 97380 0 0 $X=243670 $Y=97150
X10403 3 digital_ldo_top_VIA10 $T=244140 101460 0 0 $X=243670 $Y=101230
X10404 3 digital_ldo_top_VIA10 $T=244140 105540 0 0 $X=243670 $Y=105310
X10405 3 digital_ldo_top_VIA10 $T=244140 109620 0 0 $X=243670 $Y=109390
X10406 3 digital_ldo_top_VIA10 $T=244140 113700 0 0 $X=243670 $Y=113470
X10407 3 digital_ldo_top_VIA10 $T=244140 117780 0 0 $X=243670 $Y=117550
X10408 3 digital_ldo_top_VIA10 $T=244140 121860 0 0 $X=243670 $Y=121630
X10409 3 digital_ldo_top_VIA10 $T=244140 125940 0 0 $X=243670 $Y=125710
X10410 2 digital_ldo_top_VIA10 $T=245980 13060 0 0 $X=245510 $Y=12830
X10411 2 digital_ldo_top_VIA10 $T=245980 17140 0 0 $X=245510 $Y=16910
X10412 2 digital_ldo_top_VIA10 $T=245980 21220 0 0 $X=245510 $Y=20990
X10413 2 digital_ldo_top_VIA10 $T=245980 25300 0 0 $X=245510 $Y=25070
X10414 2 digital_ldo_top_VIA10 $T=245980 86500 0 0 $X=245510 $Y=86270
X10415 2 digital_ldo_top_VIA10 $T=245980 90580 0 0 $X=245510 $Y=90350
X10416 2 digital_ldo_top_VIA10 $T=245980 94660 0 0 $X=245510 $Y=94430
X10417 2 digital_ldo_top_VIA10 $T=245980 98740 0 0 $X=245510 $Y=98510
X10418 2 digital_ldo_top_VIA10 $T=245980 102820 0 0 $X=245510 $Y=102590
X10419 2 digital_ldo_top_VIA10 $T=245980 106900 0 0 $X=245510 $Y=106670
X10420 2 digital_ldo_top_VIA10 $T=245980 110980 0 0 $X=245510 $Y=110750
X10421 2 digital_ldo_top_VIA10 $T=245980 115060 0 0 $X=245510 $Y=114830
X10422 2 digital_ldo_top_VIA10 $T=245980 119140 0 0 $X=245510 $Y=118910
X10423 2 digital_ldo_top_VIA10 $T=245980 123220 0 0 $X=245510 $Y=122990
X10424 2 digital_ldo_top_VIA10 $T=245980 127300 0 0 $X=245510 $Y=127070
X10425 3 digital_ldo_top_VIA10 $T=249660 11700 0 0 $X=249190 $Y=11470
X10426 3 digital_ldo_top_VIA10 $T=249660 15780 0 0 $X=249190 $Y=15550
X10427 3 digital_ldo_top_VIA10 $T=249660 19860 0 0 $X=249190 $Y=19630
X10428 3 digital_ldo_top_VIA10 $T=249660 23940 0 0 $X=249190 $Y=23710
X10429 3 digital_ldo_top_VIA10 $T=249660 32100 0 0 $X=249190 $Y=31870
X10430 3 digital_ldo_top_VIA10 $T=249660 85140 0 0 $X=249190 $Y=84910
X10431 3 digital_ldo_top_VIA10 $T=249660 89220 0 0 $X=249190 $Y=88990
X10432 3 digital_ldo_top_VIA10 $T=249660 93300 0 0 $X=249190 $Y=93070
X10433 3 digital_ldo_top_VIA10 $T=249660 97380 0 0 $X=249190 $Y=97150
X10434 3 digital_ldo_top_VIA10 $T=249660 101460 0 0 $X=249190 $Y=101230
X10435 3 digital_ldo_top_VIA10 $T=249660 105540 0 0 $X=249190 $Y=105310
X10436 3 digital_ldo_top_VIA10 $T=249660 109620 0 0 $X=249190 $Y=109390
X10437 3 digital_ldo_top_VIA10 $T=249660 113700 0 0 $X=249190 $Y=113470
X10438 3 digital_ldo_top_VIA10 $T=249660 117780 0 0 $X=249190 $Y=117550
X10439 3 digital_ldo_top_VIA10 $T=249660 121860 0 0 $X=249190 $Y=121630
X10440 3 digital_ldo_top_VIA10 $T=249660 125940 0 0 $X=249190 $Y=125710
X10441 2 digital_ldo_top_VIA10 $T=251500 13060 0 0 $X=251030 $Y=12830
X10442 2 digital_ldo_top_VIA10 $T=251500 17140 0 0 $X=251030 $Y=16910
X10443 2 digital_ldo_top_VIA10 $T=251500 21220 0 0 $X=251030 $Y=20990
X10444 2 digital_ldo_top_VIA10 $T=251500 25300 0 0 $X=251030 $Y=25070
X10445 2 digital_ldo_top_VIA10 $T=251500 86500 0 0 $X=251030 $Y=86270
X10446 2 digital_ldo_top_VIA10 $T=251500 90580 0 0 $X=251030 $Y=90350
X10447 2 digital_ldo_top_VIA10 $T=251500 94660 0 0 $X=251030 $Y=94430
X10448 2 digital_ldo_top_VIA10 $T=251500 98740 0 0 $X=251030 $Y=98510
X10449 2 digital_ldo_top_VIA10 $T=251500 102820 0 0 $X=251030 $Y=102590
X10450 2 digital_ldo_top_VIA10 $T=251500 106900 0 0 $X=251030 $Y=106670
X10451 2 digital_ldo_top_VIA10 $T=251500 110980 0 0 $X=251030 $Y=110750
X10452 2 digital_ldo_top_VIA10 $T=251500 115060 0 0 $X=251030 $Y=114830
X10453 2 digital_ldo_top_VIA10 $T=251500 119140 0 0 $X=251030 $Y=118910
X10454 2 digital_ldo_top_VIA10 $T=251500 123220 0 0 $X=251030 $Y=122990
X10455 2 digital_ldo_top_VIA10 $T=251500 127300 0 0 $X=251030 $Y=127070
X10456 3 digital_ldo_top_VIA10 $T=255180 11700 0 0 $X=254710 $Y=11470
X10457 3 digital_ldo_top_VIA10 $T=255180 15780 0 0 $X=254710 $Y=15550
X10458 3 digital_ldo_top_VIA10 $T=255180 19860 0 0 $X=254710 $Y=19630
X10459 3 digital_ldo_top_VIA10 $T=255180 23940 0 0 $X=254710 $Y=23710
X10460 3 digital_ldo_top_VIA10 $T=255180 32100 0 0 $X=254710 $Y=31870
X10461 3 digital_ldo_top_VIA10 $T=255180 85140 0 0 $X=254710 $Y=84910
X10462 3 digital_ldo_top_VIA10 $T=255180 89220 0 0 $X=254710 $Y=88990
X10463 3 digital_ldo_top_VIA10 $T=255180 93300 0 0 $X=254710 $Y=93070
X10464 3 digital_ldo_top_VIA10 $T=255180 97380 0 0 $X=254710 $Y=97150
X10465 3 digital_ldo_top_VIA10 $T=255180 101460 0 0 $X=254710 $Y=101230
X10466 3 digital_ldo_top_VIA10 $T=255180 105540 0 0 $X=254710 $Y=105310
X10467 3 digital_ldo_top_VIA10 $T=255180 109620 0 0 $X=254710 $Y=109390
X10468 3 digital_ldo_top_VIA10 $T=255180 113700 0 0 $X=254710 $Y=113470
X10469 3 digital_ldo_top_VIA10 $T=255180 117780 0 0 $X=254710 $Y=117550
X10470 3 digital_ldo_top_VIA10 $T=255180 121860 0 0 $X=254710 $Y=121630
X10471 3 digital_ldo_top_VIA10 $T=255180 125940 0 0 $X=254710 $Y=125710
X10472 2 digital_ldo_top_VIA10 $T=257020 13060 0 0 $X=256550 $Y=12830
X10473 2 digital_ldo_top_VIA10 $T=257020 17140 0 0 $X=256550 $Y=16910
X10474 2 digital_ldo_top_VIA10 $T=257020 21220 0 0 $X=256550 $Y=20990
X10475 2 digital_ldo_top_VIA10 $T=257020 86500 0 0 $X=256550 $Y=86270
X10476 2 digital_ldo_top_VIA10 $T=257020 90580 0 0 $X=256550 $Y=90350
X10477 2 digital_ldo_top_VIA10 $T=257020 94660 0 0 $X=256550 $Y=94430
X10478 2 digital_ldo_top_VIA10 $T=257020 98740 0 0 $X=256550 $Y=98510
X10479 2 digital_ldo_top_VIA10 $T=257020 102820 0 0 $X=256550 $Y=102590
X10480 2 digital_ldo_top_VIA10 $T=257020 106900 0 0 $X=256550 $Y=106670
X10481 2 digital_ldo_top_VIA10 $T=257020 110980 0 0 $X=256550 $Y=110750
X10482 2 digital_ldo_top_VIA10 $T=257020 115060 0 0 $X=256550 $Y=114830
X10483 2 digital_ldo_top_VIA10 $T=257020 119140 0 0 $X=256550 $Y=118910
X10484 2 digital_ldo_top_VIA10 $T=257020 123220 0 0 $X=256550 $Y=122990
X10485 2 digital_ldo_top_VIA10 $T=257020 127300 0 0 $X=256550 $Y=127070
X10486 3 digital_ldo_top_VIA10 $T=260700 11700 0 0 $X=260230 $Y=11470
X10487 3 digital_ldo_top_VIA10 $T=260700 15780 0 0 $X=260230 $Y=15550
X10488 3 digital_ldo_top_VIA10 $T=260700 19860 0 0 $X=260230 $Y=19630
X10489 3 digital_ldo_top_VIA10 $T=260700 23940 0 0 $X=260230 $Y=23710
X10490 3 digital_ldo_top_VIA10 $T=260700 32100 0 0 $X=260230 $Y=31870
X10491 3 digital_ldo_top_VIA10 $T=260700 85140 0 0 $X=260230 $Y=84910
X10492 3 digital_ldo_top_VIA10 $T=260700 89220 0 0 $X=260230 $Y=88990
X10493 3 digital_ldo_top_VIA10 $T=260700 93300 0 0 $X=260230 $Y=93070
X10494 3 digital_ldo_top_VIA10 $T=260700 97380 0 0 $X=260230 $Y=97150
X10495 3 digital_ldo_top_VIA10 $T=260700 101460 0 0 $X=260230 $Y=101230
X10496 3 digital_ldo_top_VIA10 $T=260700 105540 0 0 $X=260230 $Y=105310
X10497 3 digital_ldo_top_VIA10 $T=260700 109620 0 0 $X=260230 $Y=109390
X10498 3 digital_ldo_top_VIA10 $T=260700 113700 0 0 $X=260230 $Y=113470
X10499 3 digital_ldo_top_VIA10 $T=260700 117780 0 0 $X=260230 $Y=117550
X10500 3 digital_ldo_top_VIA10 $T=260700 121860 0 0 $X=260230 $Y=121630
X10501 3 digital_ldo_top_VIA10 $T=260700 125940 0 0 $X=260230 $Y=125710
X10502 2 digital_ldo_top_VIA10 $T=262540 13060 0 0 $X=262070 $Y=12830
X10503 2 digital_ldo_top_VIA10 $T=262540 17140 0 0 $X=262070 $Y=16910
X10504 2 digital_ldo_top_VIA10 $T=262540 21220 0 0 $X=262070 $Y=20990
X10505 2 digital_ldo_top_VIA10 $T=262540 25300 0 0 $X=262070 $Y=25070
X10506 2 digital_ldo_top_VIA10 $T=262540 86500 0 0 $X=262070 $Y=86270
X10507 2 digital_ldo_top_VIA10 $T=262540 90580 0 0 $X=262070 $Y=90350
X10508 2 digital_ldo_top_VIA10 $T=262540 94660 0 0 $X=262070 $Y=94430
X10509 2 digital_ldo_top_VIA10 $T=262540 98740 0 0 $X=262070 $Y=98510
X10510 2 digital_ldo_top_VIA10 $T=262540 102820 0 0 $X=262070 $Y=102590
X10511 2 digital_ldo_top_VIA10 $T=262540 106900 0 0 $X=262070 $Y=106670
X10512 2 digital_ldo_top_VIA10 $T=262540 110980 0 0 $X=262070 $Y=110750
X10513 2 digital_ldo_top_VIA10 $T=262540 115060 0 0 $X=262070 $Y=114830
X10514 2 digital_ldo_top_VIA10 $T=262540 119140 0 0 $X=262070 $Y=118910
X10515 2 digital_ldo_top_VIA10 $T=262540 123220 0 0 $X=262070 $Y=122990
X10516 2 digital_ldo_top_VIA10 $T=262540 127300 0 0 $X=262070 $Y=127070
X10517 3 digital_ldo_top_VIA10 $T=266220 11700 0 0 $X=265750 $Y=11470
X10518 3 digital_ldo_top_VIA10 $T=266220 15780 0 0 $X=265750 $Y=15550
X10519 3 digital_ldo_top_VIA10 $T=266220 19860 0 0 $X=265750 $Y=19630
X10520 3 digital_ldo_top_VIA10 $T=266220 23940 0 0 $X=265750 $Y=23710
X10521 3 digital_ldo_top_VIA10 $T=266220 32100 0 0 $X=265750 $Y=31870
X10522 3 digital_ldo_top_VIA10 $T=266220 85140 0 0 $X=265750 $Y=84910
X10523 3 digital_ldo_top_VIA10 $T=266220 89220 0 0 $X=265750 $Y=88990
X10524 3 digital_ldo_top_VIA10 $T=266220 93300 0 0 $X=265750 $Y=93070
X10525 3 digital_ldo_top_VIA10 $T=266220 97380 0 0 $X=265750 $Y=97150
X10526 3 digital_ldo_top_VIA10 $T=266220 101460 0 0 $X=265750 $Y=101230
X10527 3 digital_ldo_top_VIA10 $T=266220 105540 0 0 $X=265750 $Y=105310
X10528 3 digital_ldo_top_VIA10 $T=266220 109620 0 0 $X=265750 $Y=109390
X10529 3 digital_ldo_top_VIA10 $T=266220 113700 0 0 $X=265750 $Y=113470
X10530 3 digital_ldo_top_VIA10 $T=266220 117780 0 0 $X=265750 $Y=117550
X10531 3 digital_ldo_top_VIA10 $T=266220 121860 0 0 $X=265750 $Y=121630
X10532 3 digital_ldo_top_VIA10 $T=266220 125940 0 0 $X=265750 $Y=125710
X10533 2 digital_ldo_top_VIA10 $T=268060 13060 0 0 $X=267590 $Y=12830
X10534 2 digital_ldo_top_VIA10 $T=268060 17140 0 0 $X=267590 $Y=16910
X10535 2 digital_ldo_top_VIA10 $T=268060 21220 0 0 $X=267590 $Y=20990
X10536 2 digital_ldo_top_VIA10 $T=268060 25300 0 0 $X=267590 $Y=25070
X10537 2 digital_ldo_top_VIA10 $T=268060 86500 0 0 $X=267590 $Y=86270
X10538 2 digital_ldo_top_VIA10 $T=268060 90580 0 0 $X=267590 $Y=90350
X10539 2 digital_ldo_top_VIA10 $T=268060 94660 0 0 $X=267590 $Y=94430
X10540 2 digital_ldo_top_VIA10 $T=268060 98740 0 0 $X=267590 $Y=98510
X10541 2 digital_ldo_top_VIA10 $T=268060 102820 0 0 $X=267590 $Y=102590
X10542 2 digital_ldo_top_VIA10 $T=268060 106900 0 0 $X=267590 $Y=106670
X10543 2 digital_ldo_top_VIA10 $T=268060 110980 0 0 $X=267590 $Y=110750
X10544 2 digital_ldo_top_VIA10 $T=268060 115060 0 0 $X=267590 $Y=114830
X10545 2 digital_ldo_top_VIA10 $T=268060 119140 0 0 $X=267590 $Y=118910
X10546 2 digital_ldo_top_VIA10 $T=268060 123220 0 0 $X=267590 $Y=122990
X10547 2 digital_ldo_top_VIA10 $T=268060 127300 0 0 $X=267590 $Y=127070
X10548 3 digital_ldo_top_VIA10 $T=271740 11700 0 0 $X=271270 $Y=11470
X10549 3 digital_ldo_top_VIA10 $T=271740 15780 0 0 $X=271270 $Y=15550
X10550 3 digital_ldo_top_VIA10 $T=271740 19860 0 0 $X=271270 $Y=19630
X10551 3 digital_ldo_top_VIA10 $T=271740 23940 0 0 $X=271270 $Y=23710
X10552 3 digital_ldo_top_VIA10 $T=271740 32100 0 0 $X=271270 $Y=31870
X10553 3 digital_ldo_top_VIA10 $T=271740 85140 0 0 $X=271270 $Y=84910
X10554 3 digital_ldo_top_VIA10 $T=271740 89220 0 0 $X=271270 $Y=88990
X10555 3 digital_ldo_top_VIA10 $T=271740 93300 0 0 $X=271270 $Y=93070
X10556 3 digital_ldo_top_VIA10 $T=271740 97380 0 0 $X=271270 $Y=97150
X10557 3 digital_ldo_top_VIA10 $T=271740 101460 0 0 $X=271270 $Y=101230
X10558 3 digital_ldo_top_VIA10 $T=271740 105540 0 0 $X=271270 $Y=105310
X10559 3 digital_ldo_top_VIA10 $T=271740 109620 0 0 $X=271270 $Y=109390
X10560 3 digital_ldo_top_VIA10 $T=271740 113700 0 0 $X=271270 $Y=113470
X10561 3 digital_ldo_top_VIA10 $T=271740 117780 0 0 $X=271270 $Y=117550
X10562 3 digital_ldo_top_VIA10 $T=271740 121860 0 0 $X=271270 $Y=121630
X10563 3 digital_ldo_top_VIA10 $T=271740 125940 0 0 $X=271270 $Y=125710
X10564 2 digital_ldo_top_VIA10 $T=273580 13060 0 0 $X=273110 $Y=12830
X10565 2 digital_ldo_top_VIA10 $T=273580 17140 0 0 $X=273110 $Y=16910
X10566 2 digital_ldo_top_VIA10 $T=273580 21220 0 0 $X=273110 $Y=20990
X10567 2 digital_ldo_top_VIA10 $T=273580 25300 0 0 $X=273110 $Y=25070
X10568 2 digital_ldo_top_VIA10 $T=273580 86500 0 0 $X=273110 $Y=86270
X10569 2 digital_ldo_top_VIA10 $T=273580 90580 0 0 $X=273110 $Y=90350
X10570 2 digital_ldo_top_VIA10 $T=273580 94660 0 0 $X=273110 $Y=94430
X10571 2 digital_ldo_top_VIA10 $T=273580 98740 0 0 $X=273110 $Y=98510
X10572 2 digital_ldo_top_VIA10 $T=273580 102820 0 0 $X=273110 $Y=102590
X10573 2 digital_ldo_top_VIA10 $T=273580 106900 0 0 $X=273110 $Y=106670
X10574 2 digital_ldo_top_VIA10 $T=273580 110980 0 0 $X=273110 $Y=110750
X10575 2 digital_ldo_top_VIA10 $T=273580 115060 0 0 $X=273110 $Y=114830
X10576 2 digital_ldo_top_VIA10 $T=273580 119140 0 0 $X=273110 $Y=118910
X10577 2 digital_ldo_top_VIA10 $T=273580 123220 0 0 $X=273110 $Y=122990
X10578 2 digital_ldo_top_VIA10 $T=273580 127300 0 0 $X=273110 $Y=127070
X10579 3 digital_ldo_top_VIA10 $T=277260 11700 0 0 $X=276790 $Y=11470
X10580 3 digital_ldo_top_VIA10 $T=277260 15780 0 0 $X=276790 $Y=15550
X10581 3 digital_ldo_top_VIA10 $T=277260 19860 0 0 $X=276790 $Y=19630
X10582 3 digital_ldo_top_VIA10 $T=277260 23940 0 0 $X=276790 $Y=23710
X10583 3 digital_ldo_top_VIA10 $T=277260 32100 0 0 $X=276790 $Y=31870
X10584 3 digital_ldo_top_VIA10 $T=277260 85140 0 0 $X=276790 $Y=84910
X10585 3 digital_ldo_top_VIA10 $T=277260 89220 0 0 $X=276790 $Y=88990
X10586 3 digital_ldo_top_VIA10 $T=277260 93300 0 0 $X=276790 $Y=93070
X10587 3 digital_ldo_top_VIA10 $T=277260 97380 0 0 $X=276790 $Y=97150
X10588 3 digital_ldo_top_VIA10 $T=277260 101460 0 0 $X=276790 $Y=101230
X10589 3 digital_ldo_top_VIA10 $T=277260 105540 0 0 $X=276790 $Y=105310
X10590 3 digital_ldo_top_VIA10 $T=277260 109620 0 0 $X=276790 $Y=109390
X10591 3 digital_ldo_top_VIA10 $T=277260 113700 0 0 $X=276790 $Y=113470
X10592 3 digital_ldo_top_VIA10 $T=277260 117780 0 0 $X=276790 $Y=117550
X10593 3 digital_ldo_top_VIA10 $T=277260 121860 0 0 $X=276790 $Y=121630
X10594 3 digital_ldo_top_VIA10 $T=277260 125940 0 0 $X=276790 $Y=125710
X10595 2 digital_ldo_top_VIA10 $T=279100 13060 0 0 $X=278630 $Y=12830
X10596 2 digital_ldo_top_VIA10 $T=279100 17140 0 0 $X=278630 $Y=16910
X10597 2 digital_ldo_top_VIA10 $T=279100 21220 0 0 $X=278630 $Y=20990
X10598 2 digital_ldo_top_VIA10 $T=279100 25300 0 0 $X=278630 $Y=25070
X10599 2 digital_ldo_top_VIA10 $T=279100 86500 0 0 $X=278630 $Y=86270
X10600 2 digital_ldo_top_VIA10 $T=279100 90580 0 0 $X=278630 $Y=90350
X10601 2 digital_ldo_top_VIA10 $T=279100 94660 0 0 $X=278630 $Y=94430
X10602 2 digital_ldo_top_VIA10 $T=279100 98740 0 0 $X=278630 $Y=98510
X10603 2 digital_ldo_top_VIA10 $T=279100 102820 0 0 $X=278630 $Y=102590
X10604 2 digital_ldo_top_VIA10 $T=279100 106900 0 0 $X=278630 $Y=106670
X10605 2 digital_ldo_top_VIA10 $T=279100 110980 0 0 $X=278630 $Y=110750
X10606 2 digital_ldo_top_VIA10 $T=279100 115060 0 0 $X=278630 $Y=114830
X10607 2 digital_ldo_top_VIA10 $T=279100 119140 0 0 $X=278630 $Y=118910
X10608 2 digital_ldo_top_VIA10 $T=279100 123220 0 0 $X=278630 $Y=122990
X10609 2 digital_ldo_top_VIA10 $T=279100 127300 0 0 $X=278630 $Y=127070
X10610 3 digital_ldo_top_VIA10 $T=282780 11700 0 0 $X=282310 $Y=11470
X10611 3 digital_ldo_top_VIA10 $T=282780 15780 0 0 $X=282310 $Y=15550
X10612 3 digital_ldo_top_VIA10 $T=282780 19860 0 0 $X=282310 $Y=19630
X10613 3 digital_ldo_top_VIA10 $T=282780 32100 0 0 $X=282310 $Y=31870
X10614 3 digital_ldo_top_VIA10 $T=282780 85140 0 0 $X=282310 $Y=84910
X10615 3 digital_ldo_top_VIA10 $T=282780 89220 0 0 $X=282310 $Y=88990
X10616 3 digital_ldo_top_VIA10 $T=282780 93300 0 0 $X=282310 $Y=93070
X10617 3 digital_ldo_top_VIA10 $T=282780 97380 0 0 $X=282310 $Y=97150
X10618 3 digital_ldo_top_VIA10 $T=282780 101460 0 0 $X=282310 $Y=101230
X10619 3 digital_ldo_top_VIA10 $T=282780 105540 0 0 $X=282310 $Y=105310
X10620 3 digital_ldo_top_VIA10 $T=282780 109620 0 0 $X=282310 $Y=109390
X10621 3 digital_ldo_top_VIA10 $T=282780 113700 0 0 $X=282310 $Y=113470
X10622 3 digital_ldo_top_VIA10 $T=282780 117780 0 0 $X=282310 $Y=117550
X10623 3 digital_ldo_top_VIA10 $T=282780 121860 0 0 $X=282310 $Y=121630
X10624 3 digital_ldo_top_VIA10 $T=282780 125940 0 0 $X=282310 $Y=125710
X10625 2 digital_ldo_top_VIA10 $T=284620 13060 0 0 $X=284150 $Y=12830
X10626 2 digital_ldo_top_VIA10 $T=284620 17140 0 0 $X=284150 $Y=16910
X10627 2 digital_ldo_top_VIA10 $T=284620 21220 0 0 $X=284150 $Y=20990
X10628 2 digital_ldo_top_VIA10 $T=284620 25300 0 0 $X=284150 $Y=25070
X10629 2 digital_ldo_top_VIA10 $T=284620 86500 0 0 $X=284150 $Y=86270
X10630 2 digital_ldo_top_VIA10 $T=284620 90580 0 0 $X=284150 $Y=90350
X10631 2 digital_ldo_top_VIA10 $T=284620 94660 0 0 $X=284150 $Y=94430
X10632 2 digital_ldo_top_VIA10 $T=284620 98740 0 0 $X=284150 $Y=98510
X10633 2 digital_ldo_top_VIA10 $T=284620 102820 0 0 $X=284150 $Y=102590
X10634 2 digital_ldo_top_VIA10 $T=284620 106900 0 0 $X=284150 $Y=106670
X10635 2 digital_ldo_top_VIA10 $T=284620 110980 0 0 $X=284150 $Y=110750
X10636 2 digital_ldo_top_VIA10 $T=284620 115060 0 0 $X=284150 $Y=114830
X10637 2 digital_ldo_top_VIA10 $T=284620 119140 0 0 $X=284150 $Y=118910
X10638 2 digital_ldo_top_VIA10 $T=284620 123220 0 0 $X=284150 $Y=122990
X10639 2 digital_ldo_top_VIA10 $T=284620 127300 0 0 $X=284150 $Y=127070
X10640 3 digital_ldo_top_VIA10 $T=288300 11700 0 0 $X=287830 $Y=11470
X10641 3 digital_ldo_top_VIA10 $T=288300 15780 0 0 $X=287830 $Y=15550
X10642 3 digital_ldo_top_VIA10 $T=288300 19860 0 0 $X=287830 $Y=19630
X10643 3 digital_ldo_top_VIA10 $T=288300 23940 0 0 $X=287830 $Y=23710
X10644 3 digital_ldo_top_VIA10 $T=288300 32100 0 0 $X=287830 $Y=31870
X10645 3 digital_ldo_top_VIA10 $T=288300 85140 0 0 $X=287830 $Y=84910
X10646 3 digital_ldo_top_VIA10 $T=288300 89220 0 0 $X=287830 $Y=88990
X10647 3 digital_ldo_top_VIA10 $T=288300 93300 0 0 $X=287830 $Y=93070
X10648 3 digital_ldo_top_VIA10 $T=288300 97380 0 0 $X=287830 $Y=97150
X10649 3 digital_ldo_top_VIA10 $T=288300 101460 0 0 $X=287830 $Y=101230
X10650 3 digital_ldo_top_VIA10 $T=288300 105540 0 0 $X=287830 $Y=105310
X10651 3 digital_ldo_top_VIA10 $T=288300 109620 0 0 $X=287830 $Y=109390
X10652 3 digital_ldo_top_VIA10 $T=288300 113700 0 0 $X=287830 $Y=113470
X10653 3 digital_ldo_top_VIA10 $T=288300 117780 0 0 $X=287830 $Y=117550
X10654 3 digital_ldo_top_VIA10 $T=288300 121860 0 0 $X=287830 $Y=121630
X10655 3 digital_ldo_top_VIA10 $T=288300 125940 0 0 $X=287830 $Y=125710
X10656 2 digital_ldo_top_VIA10 $T=290140 13060 0 0 $X=289670 $Y=12830
X10657 2 digital_ldo_top_VIA10 $T=290140 17140 0 0 $X=289670 $Y=16910
X10658 2 digital_ldo_top_VIA10 $T=290140 21220 0 0 $X=289670 $Y=20990
X10659 2 digital_ldo_top_VIA10 $T=290140 25300 0 0 $X=289670 $Y=25070
X10660 2 digital_ldo_top_VIA10 $T=290140 86500 0 0 $X=289670 $Y=86270
X10661 2 digital_ldo_top_VIA10 $T=290140 90580 0 0 $X=289670 $Y=90350
X10662 2 digital_ldo_top_VIA10 $T=290140 94660 0 0 $X=289670 $Y=94430
X10663 2 digital_ldo_top_VIA10 $T=290140 98740 0 0 $X=289670 $Y=98510
X10664 2 digital_ldo_top_VIA10 $T=290140 102820 0 0 $X=289670 $Y=102590
X10665 2 digital_ldo_top_VIA10 $T=290140 106900 0 0 $X=289670 $Y=106670
X10666 2 digital_ldo_top_VIA10 $T=290140 110980 0 0 $X=289670 $Y=110750
X10667 2 digital_ldo_top_VIA10 $T=290140 115060 0 0 $X=289670 $Y=114830
X10668 2 digital_ldo_top_VIA10 $T=290140 119140 0 0 $X=289670 $Y=118910
X10669 2 digital_ldo_top_VIA10 $T=290140 123220 0 0 $X=289670 $Y=122990
X10670 2 digital_ldo_top_VIA10 $T=290140 127300 0 0 $X=289670 $Y=127070
X10671 3 digital_ldo_top_VIA10 $T=293820 11700 0 0 $X=293350 $Y=11470
X10672 3 digital_ldo_top_VIA10 $T=293820 15780 0 0 $X=293350 $Y=15550
X10673 3 digital_ldo_top_VIA10 $T=293820 19860 0 0 $X=293350 $Y=19630
X10674 3 digital_ldo_top_VIA10 $T=293820 85140 0 0 $X=293350 $Y=84910
X10675 3 digital_ldo_top_VIA10 $T=293820 89220 0 0 $X=293350 $Y=88990
X10676 3 digital_ldo_top_VIA10 $T=293820 93300 0 0 $X=293350 $Y=93070
X10677 3 digital_ldo_top_VIA10 $T=293820 97380 0 0 $X=293350 $Y=97150
X10678 3 digital_ldo_top_VIA10 $T=293820 101460 0 0 $X=293350 $Y=101230
X10679 3 digital_ldo_top_VIA10 $T=293820 105540 0 0 $X=293350 $Y=105310
X10680 3 digital_ldo_top_VIA10 $T=293820 109620 0 0 $X=293350 $Y=109390
X10681 3 digital_ldo_top_VIA10 $T=293820 113700 0 0 $X=293350 $Y=113470
X10682 3 digital_ldo_top_VIA10 $T=293820 117780 0 0 $X=293350 $Y=117550
X10683 3 digital_ldo_top_VIA10 $T=293820 121860 0 0 $X=293350 $Y=121630
X10684 3 digital_ldo_top_VIA10 $T=293820 125940 0 0 $X=293350 $Y=125710
X10685 2 digital_ldo_top_VIA10 $T=295660 13060 0 0 $X=295190 $Y=12830
X10686 2 digital_ldo_top_VIA10 $T=295660 17140 0 0 $X=295190 $Y=16910
X10687 2 digital_ldo_top_VIA10 $T=295660 21220 0 0 $X=295190 $Y=20990
X10688 2 digital_ldo_top_VIA10 $T=295660 25300 0 0 $X=295190 $Y=25070
X10689 2 digital_ldo_top_VIA10 $T=295660 86500 0 0 $X=295190 $Y=86270
X10690 2 digital_ldo_top_VIA10 $T=295660 90580 0 0 $X=295190 $Y=90350
X10691 2 digital_ldo_top_VIA10 $T=295660 94660 0 0 $X=295190 $Y=94430
X10692 2 digital_ldo_top_VIA10 $T=295660 98740 0 0 $X=295190 $Y=98510
X10693 2 digital_ldo_top_VIA10 $T=295660 102820 0 0 $X=295190 $Y=102590
X10694 2 digital_ldo_top_VIA10 $T=295660 106900 0 0 $X=295190 $Y=106670
X10695 2 digital_ldo_top_VIA10 $T=295660 110980 0 0 $X=295190 $Y=110750
X10696 2 digital_ldo_top_VIA10 $T=295660 115060 0 0 $X=295190 $Y=114830
X10697 2 digital_ldo_top_VIA10 $T=295660 119140 0 0 $X=295190 $Y=118910
X10698 2 digital_ldo_top_VIA10 $T=295660 123220 0 0 $X=295190 $Y=122990
X10699 2 digital_ldo_top_VIA10 $T=295660 127300 0 0 $X=295190 $Y=127070
X10700 3 digital_ldo_top_VIA10 $T=299340 11700 0 0 $X=298870 $Y=11470
X10701 3 digital_ldo_top_VIA10 $T=299340 15780 0 0 $X=298870 $Y=15550
X10702 3 digital_ldo_top_VIA10 $T=299340 19860 0 0 $X=298870 $Y=19630
X10703 3 digital_ldo_top_VIA10 $T=299340 23940 0 0 $X=298870 $Y=23710
X10704 3 digital_ldo_top_VIA10 $T=299340 32100 0 0 $X=298870 $Y=31870
X10705 3 digital_ldo_top_VIA10 $T=299340 85140 0 0 $X=298870 $Y=84910
X10706 3 digital_ldo_top_VIA10 $T=299340 89220 0 0 $X=298870 $Y=88990
X10707 3 digital_ldo_top_VIA10 $T=299340 93300 0 0 $X=298870 $Y=93070
X10708 3 digital_ldo_top_VIA10 $T=299340 97380 0 0 $X=298870 $Y=97150
X10709 3 digital_ldo_top_VIA10 $T=299340 101460 0 0 $X=298870 $Y=101230
X10710 3 digital_ldo_top_VIA10 $T=299340 105540 0 0 $X=298870 $Y=105310
X10711 3 digital_ldo_top_VIA10 $T=299340 109620 0 0 $X=298870 $Y=109390
X10712 3 digital_ldo_top_VIA10 $T=299340 113700 0 0 $X=298870 $Y=113470
X10713 3 digital_ldo_top_VIA10 $T=299340 117780 0 0 $X=298870 $Y=117550
X10714 3 digital_ldo_top_VIA10 $T=299340 121860 0 0 $X=298870 $Y=121630
X10715 3 digital_ldo_top_VIA10 $T=299340 125940 0 0 $X=298870 $Y=125710
X10716 2 digital_ldo_top_VIA10 $T=301180 13060 0 0 $X=300710 $Y=12830
X10717 2 digital_ldo_top_VIA10 $T=301180 17140 0 0 $X=300710 $Y=16910
X10718 2 digital_ldo_top_VIA10 $T=301180 21220 0 0 $X=300710 $Y=20990
X10719 2 digital_ldo_top_VIA10 $T=301180 25300 0 0 $X=300710 $Y=25070
X10720 2 digital_ldo_top_VIA10 $T=301180 86500 0 0 $X=300710 $Y=86270
X10721 2 digital_ldo_top_VIA10 $T=301180 90580 0 0 $X=300710 $Y=90350
X10722 2 digital_ldo_top_VIA10 $T=301180 94660 0 0 $X=300710 $Y=94430
X10723 2 digital_ldo_top_VIA10 $T=301180 98740 0 0 $X=300710 $Y=98510
X10724 2 digital_ldo_top_VIA10 $T=301180 102820 0 0 $X=300710 $Y=102590
X10725 2 digital_ldo_top_VIA10 $T=301180 106900 0 0 $X=300710 $Y=106670
X10726 2 digital_ldo_top_VIA10 $T=301180 110980 0 0 $X=300710 $Y=110750
X10727 2 digital_ldo_top_VIA10 $T=301180 115060 0 0 $X=300710 $Y=114830
X10728 2 digital_ldo_top_VIA10 $T=301180 119140 0 0 $X=300710 $Y=118910
X10729 2 digital_ldo_top_VIA10 $T=301180 123220 0 0 $X=300710 $Y=122990
X10730 2 digital_ldo_top_VIA10 $T=301180 127300 0 0 $X=300710 $Y=127070
X10731 3 digital_ldo_top_VIA10 $T=304860 11700 0 0 $X=304390 $Y=11470
X10732 3 digital_ldo_top_VIA10 $T=304860 15780 0 0 $X=304390 $Y=15550
X10733 3 digital_ldo_top_VIA10 $T=304860 19860 0 0 $X=304390 $Y=19630
X10734 3 digital_ldo_top_VIA10 $T=304860 23940 0 0 $X=304390 $Y=23710
X10735 3 digital_ldo_top_VIA10 $T=304860 32100 0 0 $X=304390 $Y=31870
X10736 3 digital_ldo_top_VIA10 $T=304860 85140 0 0 $X=304390 $Y=84910
X10737 3 digital_ldo_top_VIA10 $T=304860 89220 0 0 $X=304390 $Y=88990
X10738 3 digital_ldo_top_VIA10 $T=304860 93300 0 0 $X=304390 $Y=93070
X10739 3 digital_ldo_top_VIA10 $T=304860 97380 0 0 $X=304390 $Y=97150
X10740 3 digital_ldo_top_VIA10 $T=304860 101460 0 0 $X=304390 $Y=101230
X10741 3 digital_ldo_top_VIA10 $T=304860 105540 0 0 $X=304390 $Y=105310
X10742 3 digital_ldo_top_VIA10 $T=304860 109620 0 0 $X=304390 $Y=109390
X10743 3 digital_ldo_top_VIA10 $T=304860 113700 0 0 $X=304390 $Y=113470
X10744 3 digital_ldo_top_VIA10 $T=304860 117780 0 0 $X=304390 $Y=117550
X10745 3 digital_ldo_top_VIA10 $T=304860 121860 0 0 $X=304390 $Y=121630
X10746 3 digital_ldo_top_VIA10 $T=304860 125940 0 0 $X=304390 $Y=125710
X10747 2 digital_ldo_top_VIA10 $T=306700 13060 0 0 $X=306230 $Y=12830
X10748 2 digital_ldo_top_VIA10 $T=306700 17140 0 0 $X=306230 $Y=16910
X10749 2 digital_ldo_top_VIA10 $T=306700 21220 0 0 $X=306230 $Y=20990
X10750 2 digital_ldo_top_VIA10 $T=306700 25300 0 0 $X=306230 $Y=25070
X10751 2 digital_ldo_top_VIA10 $T=306700 86500 0 0 $X=306230 $Y=86270
X10752 2 digital_ldo_top_VIA10 $T=306700 90580 0 0 $X=306230 $Y=90350
X10753 2 digital_ldo_top_VIA10 $T=306700 94660 0 0 $X=306230 $Y=94430
X10754 2 digital_ldo_top_VIA10 $T=306700 98740 0 0 $X=306230 $Y=98510
X10755 2 digital_ldo_top_VIA10 $T=306700 102820 0 0 $X=306230 $Y=102590
X10756 2 digital_ldo_top_VIA10 $T=306700 106900 0 0 $X=306230 $Y=106670
X10757 2 digital_ldo_top_VIA10 $T=306700 110980 0 0 $X=306230 $Y=110750
X10758 2 digital_ldo_top_VIA10 $T=306700 115060 0 0 $X=306230 $Y=114830
X10759 2 digital_ldo_top_VIA10 $T=306700 119140 0 0 $X=306230 $Y=118910
X10760 2 digital_ldo_top_VIA10 $T=306700 123220 0 0 $X=306230 $Y=122990
X10761 2 digital_ldo_top_VIA10 $T=306700 127300 0 0 $X=306230 $Y=127070
X10762 3 digital_ldo_top_VIA10 $T=310380 11700 0 0 $X=309910 $Y=11470
X10763 3 digital_ldo_top_VIA10 $T=310380 15780 0 0 $X=309910 $Y=15550
X10764 3 digital_ldo_top_VIA10 $T=310380 19860 0 0 $X=309910 $Y=19630
X10765 3 digital_ldo_top_VIA10 $T=310380 23940 0 0 $X=309910 $Y=23710
X10766 3 digital_ldo_top_VIA10 $T=310380 28020 0 0 $X=309910 $Y=27790
X10767 3 digital_ldo_top_VIA10 $T=310380 32100 0 0 $X=309910 $Y=31870
X10768 3 digital_ldo_top_VIA10 $T=310380 36180 0 0 $X=309910 $Y=35950
X10769 3 digital_ldo_top_VIA10 $T=310380 40260 0 0 $X=309910 $Y=40030
X10770 3 digital_ldo_top_VIA10 $T=310380 44340 0 0 $X=309910 $Y=44110
X10771 3 digital_ldo_top_VIA10 $T=310380 48420 0 0 $X=309910 $Y=48190
X10772 3 digital_ldo_top_VIA10 $T=310380 52500 0 0 $X=309910 $Y=52270
X10773 3 digital_ldo_top_VIA10 $T=310380 56580 0 0 $X=309910 $Y=56350
X10774 3 digital_ldo_top_VIA10 $T=310380 60660 0 0 $X=309910 $Y=60430
X10775 3 digital_ldo_top_VIA10 $T=310380 64740 0 0 $X=309910 $Y=64510
X10776 3 digital_ldo_top_VIA10 $T=310380 68820 0 0 $X=309910 $Y=68590
X10777 3 digital_ldo_top_VIA10 $T=310380 72900 0 0 $X=309910 $Y=72670
X10778 3 digital_ldo_top_VIA10 $T=310380 76980 0 0 $X=309910 $Y=76750
X10779 3 digital_ldo_top_VIA10 $T=310380 81060 0 0 $X=309910 $Y=80830
X10780 3 digital_ldo_top_VIA10 $T=310380 85140 0 0 $X=309910 $Y=84910
X10781 3 digital_ldo_top_VIA10 $T=310380 89220 0 0 $X=309910 $Y=88990
X10782 3 digital_ldo_top_VIA10 $T=310380 93300 0 0 $X=309910 $Y=93070
X10783 3 digital_ldo_top_VIA10 $T=310380 97380 0 0 $X=309910 $Y=97150
X10784 3 digital_ldo_top_VIA10 $T=310380 101460 0 0 $X=309910 $Y=101230
X10785 3 digital_ldo_top_VIA10 $T=310380 105540 0 0 $X=309910 $Y=105310
X10786 3 digital_ldo_top_VIA10 $T=310380 109620 0 0 $X=309910 $Y=109390
X10787 3 digital_ldo_top_VIA10 $T=310380 113700 0 0 $X=309910 $Y=113470
X10788 3 digital_ldo_top_VIA10 $T=310380 117780 0 0 $X=309910 $Y=117550
X10789 3 digital_ldo_top_VIA10 $T=310380 121860 0 0 $X=309910 $Y=121630
X10790 3 digital_ldo_top_VIA10 $T=310380 125940 0 0 $X=309910 $Y=125710
X10791 2 digital_ldo_top_VIA10 $T=312220 13060 0 0 $X=311750 $Y=12830
X10792 2 digital_ldo_top_VIA10 $T=312220 17140 0 0 $X=311750 $Y=16910
X10793 2 digital_ldo_top_VIA10 $T=312220 21220 0 0 $X=311750 $Y=20990
X10794 2 digital_ldo_top_VIA10 $T=312220 25300 0 0 $X=311750 $Y=25070
X10795 2 digital_ldo_top_VIA10 $T=312220 29380 0 0 $X=311750 $Y=29150
X10796 2 digital_ldo_top_VIA10 $T=312220 33460 0 0 $X=311750 $Y=33230
X10797 2 digital_ldo_top_VIA10 $T=312220 37540 0 0 $X=311750 $Y=37310
X10798 2 digital_ldo_top_VIA10 $T=312220 41620 0 0 $X=311750 $Y=41390
X10799 2 digital_ldo_top_VIA10 $T=312220 45700 0 0 $X=311750 $Y=45470
X10800 2 digital_ldo_top_VIA10 $T=312220 49780 0 0 $X=311750 $Y=49550
X10801 2 digital_ldo_top_VIA10 $T=312220 53860 0 0 $X=311750 $Y=53630
X10802 2 digital_ldo_top_VIA10 $T=312220 57940 0 0 $X=311750 $Y=57710
X10803 2 digital_ldo_top_VIA10 $T=312220 62020 0 0 $X=311750 $Y=61790
X10804 2 digital_ldo_top_VIA10 $T=312220 66100 0 0 $X=311750 $Y=65870
X10805 2 digital_ldo_top_VIA10 $T=312220 70180 0 0 $X=311750 $Y=69950
X10806 2 digital_ldo_top_VIA10 $T=312220 74260 0 0 $X=311750 $Y=74030
X10807 2 digital_ldo_top_VIA10 $T=312220 78340 0 0 $X=311750 $Y=78110
X10808 2 digital_ldo_top_VIA10 $T=312220 82420 0 0 $X=311750 $Y=82190
X10809 2 digital_ldo_top_VIA10 $T=312220 86500 0 0 $X=311750 $Y=86270
X10810 2 digital_ldo_top_VIA10 $T=312220 90580 0 0 $X=311750 $Y=90350
X10811 2 digital_ldo_top_VIA10 $T=312220 94660 0 0 $X=311750 $Y=94430
X10812 2 digital_ldo_top_VIA10 $T=312220 98740 0 0 $X=311750 $Y=98510
X10813 2 digital_ldo_top_VIA10 $T=312220 102820 0 0 $X=311750 $Y=102590
X10814 2 digital_ldo_top_VIA10 $T=312220 106900 0 0 $X=311750 $Y=106670
X10815 2 digital_ldo_top_VIA10 $T=312220 110980 0 0 $X=311750 $Y=110750
X10816 2 digital_ldo_top_VIA10 $T=312220 115060 0 0 $X=311750 $Y=114830
X10817 2 digital_ldo_top_VIA10 $T=312220 119140 0 0 $X=311750 $Y=118910
X10818 2 digital_ldo_top_VIA10 $T=312220 123220 0 0 $X=311750 $Y=122990
X10819 2 digital_ldo_top_VIA10 $T=312220 127300 0 0 $X=311750 $Y=127070
X10820 3 digital_ldo_top_VIA10 $T=315900 11700 0 0 $X=315430 $Y=11470
X10821 3 digital_ldo_top_VIA10 $T=315900 15780 0 0 $X=315430 $Y=15550
X10822 3 digital_ldo_top_VIA10 $T=315900 19860 0 0 $X=315430 $Y=19630
X10823 3 digital_ldo_top_VIA10 $T=315900 23940 0 0 $X=315430 $Y=23710
X10824 3 digital_ldo_top_VIA10 $T=315900 28020 0 0 $X=315430 $Y=27790
X10825 3 digital_ldo_top_VIA10 $T=315900 32100 0 0 $X=315430 $Y=31870
X10826 3 digital_ldo_top_VIA10 $T=315900 36180 0 0 $X=315430 $Y=35950
X10827 3 digital_ldo_top_VIA10 $T=315900 40260 0 0 $X=315430 $Y=40030
X10828 3 digital_ldo_top_VIA10 $T=315900 44340 0 0 $X=315430 $Y=44110
X10829 3 digital_ldo_top_VIA10 $T=315900 48420 0 0 $X=315430 $Y=48190
X10830 3 digital_ldo_top_VIA10 $T=315900 52500 0 0 $X=315430 $Y=52270
X10831 3 digital_ldo_top_VIA10 $T=315900 56580 0 0 $X=315430 $Y=56350
X10832 3 digital_ldo_top_VIA10 $T=315900 60660 0 0 $X=315430 $Y=60430
X10833 3 digital_ldo_top_VIA10 $T=315900 64740 0 0 $X=315430 $Y=64510
X10834 3 digital_ldo_top_VIA10 $T=315900 68820 0 0 $X=315430 $Y=68590
X10835 3 digital_ldo_top_VIA10 $T=315900 72900 0 0 $X=315430 $Y=72670
X10836 3 digital_ldo_top_VIA10 $T=315900 76980 0 0 $X=315430 $Y=76750
X10837 3 digital_ldo_top_VIA10 $T=315900 81060 0 0 $X=315430 $Y=80830
X10838 3 digital_ldo_top_VIA10 $T=315900 85140 0 0 $X=315430 $Y=84910
X10839 3 digital_ldo_top_VIA10 $T=315900 89220 0 0 $X=315430 $Y=88990
X10840 3 digital_ldo_top_VIA10 $T=315900 93300 0 0 $X=315430 $Y=93070
X10841 3 digital_ldo_top_VIA10 $T=315900 97380 0 0 $X=315430 $Y=97150
X10842 3 digital_ldo_top_VIA10 $T=315900 101460 0 0 $X=315430 $Y=101230
X10843 3 digital_ldo_top_VIA10 $T=315900 105540 0 0 $X=315430 $Y=105310
X10844 3 digital_ldo_top_VIA10 $T=315900 109620 0 0 $X=315430 $Y=109390
X10845 3 digital_ldo_top_VIA10 $T=315900 113700 0 0 $X=315430 $Y=113470
X10846 3 digital_ldo_top_VIA10 $T=315900 117780 0 0 $X=315430 $Y=117550
X10847 3 digital_ldo_top_VIA10 $T=315900 121860 0 0 $X=315430 $Y=121630
X10848 3 digital_ldo_top_VIA10 $T=315900 125940 0 0 $X=315430 $Y=125710
X10849 2 digital_ldo_top_VIA10 $T=317740 13060 0 0 $X=317270 $Y=12830
X10850 2 digital_ldo_top_VIA10 $T=317740 17140 0 0 $X=317270 $Y=16910
X10851 2 digital_ldo_top_VIA10 $T=317740 21220 0 0 $X=317270 $Y=20990
X10852 2 digital_ldo_top_VIA10 $T=317740 25300 0 0 $X=317270 $Y=25070
X10853 2 digital_ldo_top_VIA10 $T=317740 29380 0 0 $X=317270 $Y=29150
X10854 2 digital_ldo_top_VIA10 $T=317740 33460 0 0 $X=317270 $Y=33230
X10855 2 digital_ldo_top_VIA10 $T=317740 37540 0 0 $X=317270 $Y=37310
X10856 2 digital_ldo_top_VIA10 $T=317740 41620 0 0 $X=317270 $Y=41390
X10857 2 digital_ldo_top_VIA10 $T=317740 45700 0 0 $X=317270 $Y=45470
X10858 2 digital_ldo_top_VIA10 $T=317740 49780 0 0 $X=317270 $Y=49550
X10859 2 digital_ldo_top_VIA10 $T=317740 53860 0 0 $X=317270 $Y=53630
X10860 2 digital_ldo_top_VIA10 $T=317740 57940 0 0 $X=317270 $Y=57710
X10861 2 digital_ldo_top_VIA10 $T=317740 62020 0 0 $X=317270 $Y=61790
X10862 2 digital_ldo_top_VIA10 $T=317740 66100 0 0 $X=317270 $Y=65870
X10863 2 digital_ldo_top_VIA10 $T=317740 70180 0 0 $X=317270 $Y=69950
X10864 2 digital_ldo_top_VIA10 $T=317740 74260 0 0 $X=317270 $Y=74030
X10865 2 digital_ldo_top_VIA10 $T=317740 78340 0 0 $X=317270 $Y=78110
X10866 2 digital_ldo_top_VIA10 $T=317740 82420 0 0 $X=317270 $Y=82190
X10867 2 digital_ldo_top_VIA10 $T=317740 86500 0 0 $X=317270 $Y=86270
X10868 2 digital_ldo_top_VIA10 $T=317740 90580 0 0 $X=317270 $Y=90350
X10869 2 digital_ldo_top_VIA10 $T=317740 94660 0 0 $X=317270 $Y=94430
X10870 2 digital_ldo_top_VIA10 $T=317740 98740 0 0 $X=317270 $Y=98510
X10871 2 digital_ldo_top_VIA10 $T=317740 102820 0 0 $X=317270 $Y=102590
X10872 2 digital_ldo_top_VIA10 $T=317740 106900 0 0 $X=317270 $Y=106670
X10873 2 digital_ldo_top_VIA10 $T=317740 110980 0 0 $X=317270 $Y=110750
X10874 2 digital_ldo_top_VIA10 $T=317740 115060 0 0 $X=317270 $Y=114830
X10875 2 digital_ldo_top_VIA10 $T=317740 119140 0 0 $X=317270 $Y=118910
X10876 2 digital_ldo_top_VIA10 $T=317740 123220 0 0 $X=317270 $Y=122990
X10877 2 digital_ldo_top_VIA10 $T=317740 127300 0 0 $X=317270 $Y=127070
X10878 3 digital_ldo_top_VIA10 $T=321420 11700 0 0 $X=320950 $Y=11470
X10879 3 digital_ldo_top_VIA10 $T=321420 15780 0 0 $X=320950 $Y=15550
X10880 3 digital_ldo_top_VIA10 $T=321420 19860 0 0 $X=320950 $Y=19630
X10881 3 digital_ldo_top_VIA10 $T=321420 23940 0 0 $X=320950 $Y=23710
X10882 3 digital_ldo_top_VIA10 $T=321420 28020 0 0 $X=320950 $Y=27790
X10883 3 digital_ldo_top_VIA10 $T=321420 32100 0 0 $X=320950 $Y=31870
X10884 3 digital_ldo_top_VIA10 $T=321420 36180 0 0 $X=320950 $Y=35950
X10885 3 digital_ldo_top_VIA10 $T=321420 40260 0 0 $X=320950 $Y=40030
X10886 3 digital_ldo_top_VIA10 $T=321420 44340 0 0 $X=320950 $Y=44110
X10887 3 digital_ldo_top_VIA10 $T=321420 48420 0 0 $X=320950 $Y=48190
X10888 3 digital_ldo_top_VIA10 $T=321420 52500 0 0 $X=320950 $Y=52270
X10889 3 digital_ldo_top_VIA10 $T=321420 56580 0 0 $X=320950 $Y=56350
X10890 3 digital_ldo_top_VIA10 $T=321420 60660 0 0 $X=320950 $Y=60430
X10891 3 digital_ldo_top_VIA10 $T=321420 64740 0 0 $X=320950 $Y=64510
X10892 3 digital_ldo_top_VIA10 $T=321420 68820 0 0 $X=320950 $Y=68590
X10893 3 digital_ldo_top_VIA10 $T=321420 72900 0 0 $X=320950 $Y=72670
X10894 3 digital_ldo_top_VIA10 $T=321420 76980 0 0 $X=320950 $Y=76750
X10895 3 digital_ldo_top_VIA10 $T=321420 81060 0 0 $X=320950 $Y=80830
X10896 3 digital_ldo_top_VIA10 $T=321420 85140 0 0 $X=320950 $Y=84910
X10897 3 digital_ldo_top_VIA10 $T=321420 89220 0 0 $X=320950 $Y=88990
X10898 3 digital_ldo_top_VIA10 $T=321420 93300 0 0 $X=320950 $Y=93070
X10899 3 digital_ldo_top_VIA10 $T=321420 97380 0 0 $X=320950 $Y=97150
X10900 3 digital_ldo_top_VIA10 $T=321420 101460 0 0 $X=320950 $Y=101230
X10901 3 digital_ldo_top_VIA10 $T=321420 105540 0 0 $X=320950 $Y=105310
X10902 3 digital_ldo_top_VIA10 $T=321420 109620 0 0 $X=320950 $Y=109390
X10903 3 digital_ldo_top_VIA10 $T=321420 113700 0 0 $X=320950 $Y=113470
X10904 3 digital_ldo_top_VIA10 $T=321420 117780 0 0 $X=320950 $Y=117550
X10905 3 digital_ldo_top_VIA10 $T=321420 121860 0 0 $X=320950 $Y=121630
X10906 3 digital_ldo_top_VIA10 $T=321420 125940 0 0 $X=320950 $Y=125710
X10907 2 digital_ldo_top_VIA10 $T=323260 13060 0 0 $X=322790 $Y=12830
X10908 2 digital_ldo_top_VIA10 $T=323260 17140 0 0 $X=322790 $Y=16910
X10909 2 digital_ldo_top_VIA10 $T=323260 21220 0 0 $X=322790 $Y=20990
X10910 2 digital_ldo_top_VIA10 $T=323260 25300 0 0 $X=322790 $Y=25070
X10911 2 digital_ldo_top_VIA10 $T=323260 29380 0 0 $X=322790 $Y=29150
X10912 2 digital_ldo_top_VIA10 $T=323260 33460 0 0 $X=322790 $Y=33230
X10913 2 digital_ldo_top_VIA10 $T=323260 37540 0 0 $X=322790 $Y=37310
X10914 2 digital_ldo_top_VIA10 $T=323260 41620 0 0 $X=322790 $Y=41390
X10915 2 digital_ldo_top_VIA10 $T=323260 45700 0 0 $X=322790 $Y=45470
X10916 2 digital_ldo_top_VIA10 $T=323260 49780 0 0 $X=322790 $Y=49550
X10917 2 digital_ldo_top_VIA10 $T=323260 53860 0 0 $X=322790 $Y=53630
X10918 2 digital_ldo_top_VIA10 $T=323260 57940 0 0 $X=322790 $Y=57710
X10919 2 digital_ldo_top_VIA10 $T=323260 62020 0 0 $X=322790 $Y=61790
X10920 2 digital_ldo_top_VIA10 $T=323260 66100 0 0 $X=322790 $Y=65870
X10921 2 digital_ldo_top_VIA10 $T=323260 70180 0 0 $X=322790 $Y=69950
X10922 2 digital_ldo_top_VIA10 $T=323260 74260 0 0 $X=322790 $Y=74030
X10923 2 digital_ldo_top_VIA10 $T=323260 78340 0 0 $X=322790 $Y=78110
X10924 2 digital_ldo_top_VIA10 $T=323260 82420 0 0 $X=322790 $Y=82190
X10925 2 digital_ldo_top_VIA10 $T=323260 86500 0 0 $X=322790 $Y=86270
X10926 2 digital_ldo_top_VIA10 $T=323260 90580 0 0 $X=322790 $Y=90350
X10927 2 digital_ldo_top_VIA10 $T=323260 94660 0 0 $X=322790 $Y=94430
X10928 2 digital_ldo_top_VIA10 $T=323260 98740 0 0 $X=322790 $Y=98510
X10929 2 digital_ldo_top_VIA10 $T=323260 102820 0 0 $X=322790 $Y=102590
X10930 2 digital_ldo_top_VIA10 $T=323260 106900 0 0 $X=322790 $Y=106670
X10931 2 digital_ldo_top_VIA10 $T=323260 110980 0 0 $X=322790 $Y=110750
X10932 2 digital_ldo_top_VIA10 $T=323260 115060 0 0 $X=322790 $Y=114830
X10933 2 digital_ldo_top_VIA10 $T=323260 119140 0 0 $X=322790 $Y=118910
X10934 2 digital_ldo_top_VIA10 $T=323260 123220 0 0 $X=322790 $Y=122990
X10935 2 digital_ldo_top_VIA10 $T=323260 127300 0 0 $X=322790 $Y=127070
X10936 3 digital_ldo_top_VIA10 $T=326940 11700 0 0 $X=326470 $Y=11470
X10937 3 digital_ldo_top_VIA10 $T=326940 15780 0 0 $X=326470 $Y=15550
X10938 3 digital_ldo_top_VIA10 $T=326940 19860 0 0 $X=326470 $Y=19630
X10939 3 digital_ldo_top_VIA10 $T=326940 23940 0 0 $X=326470 $Y=23710
X10940 3 digital_ldo_top_VIA10 $T=326940 28020 0 0 $X=326470 $Y=27790
X10941 3 digital_ldo_top_VIA10 $T=326940 32100 0 0 $X=326470 $Y=31870
X10942 3 digital_ldo_top_VIA10 $T=326940 36180 0 0 $X=326470 $Y=35950
X10943 3 digital_ldo_top_VIA10 $T=326940 40260 0 0 $X=326470 $Y=40030
X10944 3 digital_ldo_top_VIA10 $T=326940 44340 0 0 $X=326470 $Y=44110
X10945 3 digital_ldo_top_VIA10 $T=326940 48420 0 0 $X=326470 $Y=48190
X10946 3 digital_ldo_top_VIA10 $T=326940 52500 0 0 $X=326470 $Y=52270
X10947 3 digital_ldo_top_VIA10 $T=326940 56580 0 0 $X=326470 $Y=56350
X10948 3 digital_ldo_top_VIA10 $T=326940 60660 0 0 $X=326470 $Y=60430
X10949 3 digital_ldo_top_VIA10 $T=326940 64740 0 0 $X=326470 $Y=64510
X10950 3 digital_ldo_top_VIA10 $T=326940 68820 0 0 $X=326470 $Y=68590
X10951 3 digital_ldo_top_VIA10 $T=326940 72900 0 0 $X=326470 $Y=72670
X10952 3 digital_ldo_top_VIA10 $T=326940 76980 0 0 $X=326470 $Y=76750
X10953 3 digital_ldo_top_VIA10 $T=326940 81060 0 0 $X=326470 $Y=80830
X10954 3 digital_ldo_top_VIA10 $T=326940 85140 0 0 $X=326470 $Y=84910
X10955 3 digital_ldo_top_VIA10 $T=326940 89220 0 0 $X=326470 $Y=88990
X10956 3 digital_ldo_top_VIA10 $T=326940 93300 0 0 $X=326470 $Y=93070
X10957 3 digital_ldo_top_VIA10 $T=326940 97380 0 0 $X=326470 $Y=97150
X10958 3 digital_ldo_top_VIA10 $T=326940 101460 0 0 $X=326470 $Y=101230
X10959 3 digital_ldo_top_VIA10 $T=326940 105540 0 0 $X=326470 $Y=105310
X10960 3 digital_ldo_top_VIA10 $T=326940 109620 0 0 $X=326470 $Y=109390
X10961 3 digital_ldo_top_VIA10 $T=326940 113700 0 0 $X=326470 $Y=113470
X10962 3 digital_ldo_top_VIA10 $T=326940 117780 0 0 $X=326470 $Y=117550
X10963 3 digital_ldo_top_VIA10 $T=326940 121860 0 0 $X=326470 $Y=121630
X10964 3 digital_ldo_top_VIA10 $T=326940 125940 0 0 $X=326470 $Y=125710
X10965 2 digital_ldo_top_VIA10 $T=328780 13060 0 0 $X=328310 $Y=12830
X10966 2 digital_ldo_top_VIA10 $T=328780 17140 0 0 $X=328310 $Y=16910
X10967 2 digital_ldo_top_VIA10 $T=328780 21220 0 0 $X=328310 $Y=20990
X10968 2 digital_ldo_top_VIA10 $T=328780 25300 0 0 $X=328310 $Y=25070
X10969 2 digital_ldo_top_VIA10 $T=328780 29380 0 0 $X=328310 $Y=29150
X10970 2 digital_ldo_top_VIA10 $T=328780 33460 0 0 $X=328310 $Y=33230
X10971 2 digital_ldo_top_VIA10 $T=328780 37540 0 0 $X=328310 $Y=37310
X10972 2 digital_ldo_top_VIA10 $T=328780 41620 0 0 $X=328310 $Y=41390
X10973 2 digital_ldo_top_VIA10 $T=328780 45700 0 0 $X=328310 $Y=45470
X10974 2 digital_ldo_top_VIA10 $T=328780 49780 0 0 $X=328310 $Y=49550
X10975 2 digital_ldo_top_VIA10 $T=328780 53860 0 0 $X=328310 $Y=53630
X10976 2 digital_ldo_top_VIA10 $T=328780 57940 0 0 $X=328310 $Y=57710
X10977 2 digital_ldo_top_VIA10 $T=328780 62020 0 0 $X=328310 $Y=61790
X10978 2 digital_ldo_top_VIA10 $T=328780 66100 0 0 $X=328310 $Y=65870
X10979 2 digital_ldo_top_VIA10 $T=328780 70180 0 0 $X=328310 $Y=69950
X10980 2 digital_ldo_top_VIA10 $T=328780 74260 0 0 $X=328310 $Y=74030
X10981 2 digital_ldo_top_VIA10 $T=328780 78340 0 0 $X=328310 $Y=78110
X10982 2 digital_ldo_top_VIA10 $T=328780 82420 0 0 $X=328310 $Y=82190
X10983 2 digital_ldo_top_VIA10 $T=328780 86500 0 0 $X=328310 $Y=86270
X10984 2 digital_ldo_top_VIA10 $T=328780 90580 0 0 $X=328310 $Y=90350
X10985 2 digital_ldo_top_VIA10 $T=328780 94660 0 0 $X=328310 $Y=94430
X10986 2 digital_ldo_top_VIA10 $T=328780 98740 0 0 $X=328310 $Y=98510
X10987 2 digital_ldo_top_VIA10 $T=328780 102820 0 0 $X=328310 $Y=102590
X10988 2 digital_ldo_top_VIA10 $T=328780 106900 0 0 $X=328310 $Y=106670
X10989 2 digital_ldo_top_VIA10 $T=328780 110980 0 0 $X=328310 $Y=110750
X10990 2 digital_ldo_top_VIA10 $T=328780 115060 0 0 $X=328310 $Y=114830
X10991 2 digital_ldo_top_VIA10 $T=328780 119140 0 0 $X=328310 $Y=118910
X10992 2 digital_ldo_top_VIA10 $T=328780 123220 0 0 $X=328310 $Y=122990
X10993 2 digital_ldo_top_VIA10 $T=328780 127300 0 0 $X=328310 $Y=127070
X10994 3 digital_ldo_top_VIA10 $T=332460 11700 0 0 $X=331990 $Y=11470
X10995 3 digital_ldo_top_VIA10 $T=332460 15780 0 0 $X=331990 $Y=15550
X10996 3 digital_ldo_top_VIA10 $T=332460 19860 0 0 $X=331990 $Y=19630
X10997 3 digital_ldo_top_VIA10 $T=332460 23940 0 0 $X=331990 $Y=23710
X10998 3 digital_ldo_top_VIA10 $T=332460 28020 0 0 $X=331990 $Y=27790
X10999 3 digital_ldo_top_VIA10 $T=332460 32100 0 0 $X=331990 $Y=31870
X11000 3 digital_ldo_top_VIA10 $T=332460 36180 0 0 $X=331990 $Y=35950
X11001 3 digital_ldo_top_VIA10 $T=332460 40260 0 0 $X=331990 $Y=40030
X11002 3 digital_ldo_top_VIA10 $T=332460 44340 0 0 $X=331990 $Y=44110
X11003 3 digital_ldo_top_VIA10 $T=332460 48420 0 0 $X=331990 $Y=48190
X11004 3 digital_ldo_top_VIA10 $T=332460 52500 0 0 $X=331990 $Y=52270
X11005 3 digital_ldo_top_VIA10 $T=332460 56580 0 0 $X=331990 $Y=56350
X11006 3 digital_ldo_top_VIA10 $T=332460 60660 0 0 $X=331990 $Y=60430
X11007 3 digital_ldo_top_VIA10 $T=332460 64740 0 0 $X=331990 $Y=64510
X11008 3 digital_ldo_top_VIA10 $T=332460 68820 0 0 $X=331990 $Y=68590
X11009 3 digital_ldo_top_VIA10 $T=332460 72900 0 0 $X=331990 $Y=72670
X11010 3 digital_ldo_top_VIA10 $T=332460 76980 0 0 $X=331990 $Y=76750
X11011 3 digital_ldo_top_VIA10 $T=332460 81060 0 0 $X=331990 $Y=80830
X11012 3 digital_ldo_top_VIA10 $T=332460 85140 0 0 $X=331990 $Y=84910
X11013 3 digital_ldo_top_VIA10 $T=332460 89220 0 0 $X=331990 $Y=88990
X11014 3 digital_ldo_top_VIA10 $T=332460 93300 0 0 $X=331990 $Y=93070
X11015 3 digital_ldo_top_VIA10 $T=332460 97380 0 0 $X=331990 $Y=97150
X11016 3 digital_ldo_top_VIA10 $T=332460 101460 0 0 $X=331990 $Y=101230
X11017 3 digital_ldo_top_VIA10 $T=332460 105540 0 0 $X=331990 $Y=105310
X11018 3 digital_ldo_top_VIA10 $T=332460 109620 0 0 $X=331990 $Y=109390
X11019 3 digital_ldo_top_VIA10 $T=332460 113700 0 0 $X=331990 $Y=113470
X11020 3 digital_ldo_top_VIA10 $T=332460 117780 0 0 $X=331990 $Y=117550
X11021 3 digital_ldo_top_VIA10 $T=332460 121860 0 0 $X=331990 $Y=121630
X11022 3 digital_ldo_top_VIA10 $T=332460 125940 0 0 $X=331990 $Y=125710
X11023 2 digital_ldo_top_VIA10 $T=334300 13060 0 0 $X=333830 $Y=12830
X11024 2 digital_ldo_top_VIA10 $T=334300 17140 0 0 $X=333830 $Y=16910
X11025 2 digital_ldo_top_VIA10 $T=334300 21220 0 0 $X=333830 $Y=20990
X11026 2 digital_ldo_top_VIA10 $T=334300 25300 0 0 $X=333830 $Y=25070
X11027 2 digital_ldo_top_VIA10 $T=334300 29380 0 0 $X=333830 $Y=29150
X11028 2 digital_ldo_top_VIA10 $T=334300 33460 0 0 $X=333830 $Y=33230
X11029 2 digital_ldo_top_VIA10 $T=334300 37540 0 0 $X=333830 $Y=37310
X11030 2 digital_ldo_top_VIA10 $T=334300 41620 0 0 $X=333830 $Y=41390
X11031 2 digital_ldo_top_VIA10 $T=334300 45700 0 0 $X=333830 $Y=45470
X11032 2 digital_ldo_top_VIA10 $T=334300 49780 0 0 $X=333830 $Y=49550
X11033 2 digital_ldo_top_VIA10 $T=334300 53860 0 0 $X=333830 $Y=53630
X11034 2 digital_ldo_top_VIA10 $T=334300 57940 0 0 $X=333830 $Y=57710
X11035 2 digital_ldo_top_VIA10 $T=334300 62020 0 0 $X=333830 $Y=61790
X11036 2 digital_ldo_top_VIA10 $T=334300 66100 0 0 $X=333830 $Y=65870
X11037 2 digital_ldo_top_VIA10 $T=334300 70180 0 0 $X=333830 $Y=69950
X11038 2 digital_ldo_top_VIA10 $T=334300 74260 0 0 $X=333830 $Y=74030
X11039 2 digital_ldo_top_VIA10 $T=334300 78340 0 0 $X=333830 $Y=78110
X11040 2 digital_ldo_top_VIA10 $T=334300 82420 0 0 $X=333830 $Y=82190
X11041 2 digital_ldo_top_VIA10 $T=334300 86500 0 0 $X=333830 $Y=86270
X11042 2 digital_ldo_top_VIA10 $T=334300 90580 0 0 $X=333830 $Y=90350
X11043 2 digital_ldo_top_VIA10 $T=334300 94660 0 0 $X=333830 $Y=94430
X11044 2 digital_ldo_top_VIA10 $T=334300 98740 0 0 $X=333830 $Y=98510
X11045 2 digital_ldo_top_VIA10 $T=334300 102820 0 0 $X=333830 $Y=102590
X11046 2 digital_ldo_top_VIA10 $T=334300 106900 0 0 $X=333830 $Y=106670
X11047 2 digital_ldo_top_VIA10 $T=334300 110980 0 0 $X=333830 $Y=110750
X11048 2 digital_ldo_top_VIA10 $T=334300 115060 0 0 $X=333830 $Y=114830
X11049 2 digital_ldo_top_VIA10 $T=334300 119140 0 0 $X=333830 $Y=118910
X11050 2 digital_ldo_top_VIA10 $T=334300 123220 0 0 $X=333830 $Y=122990
X11051 2 digital_ldo_top_VIA10 $T=334300 127300 0 0 $X=333830 $Y=127070
X11052 3 digital_ldo_top_VIA10 $T=337980 11700 0 0 $X=337510 $Y=11470
X11053 3 digital_ldo_top_VIA10 $T=337980 15780 0 0 $X=337510 $Y=15550
X11054 3 digital_ldo_top_VIA10 $T=337980 19860 0 0 $X=337510 $Y=19630
X11055 3 digital_ldo_top_VIA10 $T=337980 23940 0 0 $X=337510 $Y=23710
X11056 3 digital_ldo_top_VIA10 $T=337980 28020 0 0 $X=337510 $Y=27790
X11057 3 digital_ldo_top_VIA10 $T=337980 32100 0 0 $X=337510 $Y=31870
X11058 3 digital_ldo_top_VIA10 $T=337980 36180 0 0 $X=337510 $Y=35950
X11059 3 digital_ldo_top_VIA10 $T=337980 40260 0 0 $X=337510 $Y=40030
X11060 3 digital_ldo_top_VIA10 $T=337980 44340 0 0 $X=337510 $Y=44110
X11061 3 digital_ldo_top_VIA10 $T=337980 48420 0 0 $X=337510 $Y=48190
X11062 3 digital_ldo_top_VIA10 $T=337980 52500 0 0 $X=337510 $Y=52270
X11063 3 digital_ldo_top_VIA10 $T=337980 56580 0 0 $X=337510 $Y=56350
X11064 3 digital_ldo_top_VIA10 $T=337980 60660 0 0 $X=337510 $Y=60430
X11065 3 digital_ldo_top_VIA10 $T=337980 64740 0 0 $X=337510 $Y=64510
X11066 3 digital_ldo_top_VIA10 $T=337980 68820 0 0 $X=337510 $Y=68590
X11067 3 digital_ldo_top_VIA10 $T=337980 72900 0 0 $X=337510 $Y=72670
X11068 3 digital_ldo_top_VIA10 $T=337980 76980 0 0 $X=337510 $Y=76750
X11069 3 digital_ldo_top_VIA10 $T=337980 81060 0 0 $X=337510 $Y=80830
X11070 3 digital_ldo_top_VIA10 $T=337980 85140 0 0 $X=337510 $Y=84910
X11071 3 digital_ldo_top_VIA10 $T=337980 89220 0 0 $X=337510 $Y=88990
X11072 3 digital_ldo_top_VIA10 $T=337980 93300 0 0 $X=337510 $Y=93070
X11073 3 digital_ldo_top_VIA10 $T=337980 97380 0 0 $X=337510 $Y=97150
X11074 3 digital_ldo_top_VIA10 $T=337980 101460 0 0 $X=337510 $Y=101230
X11075 3 digital_ldo_top_VIA10 $T=337980 105540 0 0 $X=337510 $Y=105310
X11076 3 digital_ldo_top_VIA10 $T=337980 109620 0 0 $X=337510 $Y=109390
X11077 3 digital_ldo_top_VIA10 $T=337980 113700 0 0 $X=337510 $Y=113470
X11078 3 digital_ldo_top_VIA10 $T=337980 117780 0 0 $X=337510 $Y=117550
X11079 3 digital_ldo_top_VIA10 $T=337980 121860 0 0 $X=337510 $Y=121630
X11080 3 digital_ldo_top_VIA10 $T=337980 125940 0 0 $X=337510 $Y=125710
X11081 2 digital_ldo_top_VIA10 $T=339820 13060 0 0 $X=339350 $Y=12830
X11082 2 digital_ldo_top_VIA10 $T=339820 17140 0 0 $X=339350 $Y=16910
X11083 2 digital_ldo_top_VIA10 $T=339820 21220 0 0 $X=339350 $Y=20990
X11084 2 digital_ldo_top_VIA10 $T=339820 25300 0 0 $X=339350 $Y=25070
X11085 2 digital_ldo_top_VIA10 $T=339820 29380 0 0 $X=339350 $Y=29150
X11086 2 digital_ldo_top_VIA10 $T=339820 33460 0 0 $X=339350 $Y=33230
X11087 2 digital_ldo_top_VIA10 $T=339820 37540 0 0 $X=339350 $Y=37310
X11088 2 digital_ldo_top_VIA10 $T=339820 41620 0 0 $X=339350 $Y=41390
X11089 2 digital_ldo_top_VIA10 $T=339820 45700 0 0 $X=339350 $Y=45470
X11090 2 digital_ldo_top_VIA10 $T=339820 49780 0 0 $X=339350 $Y=49550
X11091 2 digital_ldo_top_VIA10 $T=339820 53860 0 0 $X=339350 $Y=53630
X11092 2 digital_ldo_top_VIA10 $T=339820 57940 0 0 $X=339350 $Y=57710
X11093 2 digital_ldo_top_VIA10 $T=339820 62020 0 0 $X=339350 $Y=61790
X11094 2 digital_ldo_top_VIA10 $T=339820 66100 0 0 $X=339350 $Y=65870
X11095 2 digital_ldo_top_VIA10 $T=339820 70180 0 0 $X=339350 $Y=69950
X11096 2 digital_ldo_top_VIA10 $T=339820 74260 0 0 $X=339350 $Y=74030
X11097 2 digital_ldo_top_VIA10 $T=339820 78340 0 0 $X=339350 $Y=78110
X11098 2 digital_ldo_top_VIA10 $T=339820 82420 0 0 $X=339350 $Y=82190
X11099 2 digital_ldo_top_VIA10 $T=339820 86500 0 0 $X=339350 $Y=86270
X11100 2 digital_ldo_top_VIA10 $T=339820 90580 0 0 $X=339350 $Y=90350
X11101 2 digital_ldo_top_VIA10 $T=339820 94660 0 0 $X=339350 $Y=94430
X11102 2 digital_ldo_top_VIA10 $T=339820 98740 0 0 $X=339350 $Y=98510
X11103 2 digital_ldo_top_VIA10 $T=339820 102820 0 0 $X=339350 $Y=102590
X11104 2 digital_ldo_top_VIA10 $T=339820 106900 0 0 $X=339350 $Y=106670
X11105 2 digital_ldo_top_VIA10 $T=339820 110980 0 0 $X=339350 $Y=110750
X11106 2 digital_ldo_top_VIA10 $T=339820 115060 0 0 $X=339350 $Y=114830
X11107 2 digital_ldo_top_VIA10 $T=339820 119140 0 0 $X=339350 $Y=118910
X11108 2 digital_ldo_top_VIA10 $T=339820 123220 0 0 $X=339350 $Y=122990
X11109 2 digital_ldo_top_VIA10 $T=339820 127300 0 0 $X=339350 $Y=127070
X11110 3 digital_ldo_top_VIA10 $T=343500 11700 0 0 $X=343030 $Y=11470
X11111 3 digital_ldo_top_VIA10 $T=343500 15780 0 0 $X=343030 $Y=15550
X11112 3 digital_ldo_top_VIA10 $T=343500 19860 0 0 $X=343030 $Y=19630
X11113 3 digital_ldo_top_VIA10 $T=343500 23940 0 0 $X=343030 $Y=23710
X11114 3 digital_ldo_top_VIA10 $T=343500 28020 0 0 $X=343030 $Y=27790
X11115 3 digital_ldo_top_VIA10 $T=343500 32100 0 0 $X=343030 $Y=31870
X11116 3 digital_ldo_top_VIA10 $T=343500 36180 0 0 $X=343030 $Y=35950
X11117 3 digital_ldo_top_VIA10 $T=343500 40260 0 0 $X=343030 $Y=40030
X11118 3 digital_ldo_top_VIA10 $T=343500 44340 0 0 $X=343030 $Y=44110
X11119 3 digital_ldo_top_VIA10 $T=343500 48420 0 0 $X=343030 $Y=48190
X11120 3 digital_ldo_top_VIA10 $T=343500 52500 0 0 $X=343030 $Y=52270
X11121 3 digital_ldo_top_VIA10 $T=343500 56580 0 0 $X=343030 $Y=56350
X11122 3 digital_ldo_top_VIA10 $T=343500 60660 0 0 $X=343030 $Y=60430
X11123 3 digital_ldo_top_VIA10 $T=343500 64740 0 0 $X=343030 $Y=64510
X11124 3 digital_ldo_top_VIA10 $T=343500 68820 0 0 $X=343030 $Y=68590
X11125 3 digital_ldo_top_VIA10 $T=343500 72900 0 0 $X=343030 $Y=72670
X11126 3 digital_ldo_top_VIA10 $T=343500 76980 0 0 $X=343030 $Y=76750
X11127 3 digital_ldo_top_VIA10 $T=343500 81060 0 0 $X=343030 $Y=80830
X11128 3 digital_ldo_top_VIA10 $T=343500 85140 0 0 $X=343030 $Y=84910
X11129 3 digital_ldo_top_VIA10 $T=343500 89220 0 0 $X=343030 $Y=88990
X11130 3 digital_ldo_top_VIA10 $T=343500 93300 0 0 $X=343030 $Y=93070
X11131 3 digital_ldo_top_VIA10 $T=343500 97380 0 0 $X=343030 $Y=97150
X11132 3 digital_ldo_top_VIA10 $T=343500 101460 0 0 $X=343030 $Y=101230
X11133 3 digital_ldo_top_VIA10 $T=343500 105540 0 0 $X=343030 $Y=105310
X11134 3 digital_ldo_top_VIA10 $T=343500 109620 0 0 $X=343030 $Y=109390
X11135 3 digital_ldo_top_VIA10 $T=343500 113700 0 0 $X=343030 $Y=113470
X11136 3 digital_ldo_top_VIA10 $T=343500 117780 0 0 $X=343030 $Y=117550
X11137 3 digital_ldo_top_VIA10 $T=343500 121860 0 0 $X=343030 $Y=121630
X11138 3 digital_ldo_top_VIA10 $T=343500 125940 0 0 $X=343030 $Y=125710
X11139 2 digital_ldo_top_VIA10 $T=345340 13060 0 0 $X=344870 $Y=12830
X11140 2 digital_ldo_top_VIA10 $T=345340 17140 0 0 $X=344870 $Y=16910
X11141 2 digital_ldo_top_VIA10 $T=345340 21220 0 0 $X=344870 $Y=20990
X11142 2 digital_ldo_top_VIA10 $T=345340 25300 0 0 $X=344870 $Y=25070
X11143 2 digital_ldo_top_VIA10 $T=345340 29380 0 0 $X=344870 $Y=29150
X11144 2 digital_ldo_top_VIA10 $T=345340 33460 0 0 $X=344870 $Y=33230
X11145 2 digital_ldo_top_VIA10 $T=345340 37540 0 0 $X=344870 $Y=37310
X11146 2 digital_ldo_top_VIA10 $T=345340 41620 0 0 $X=344870 $Y=41390
X11147 2 digital_ldo_top_VIA10 $T=345340 45700 0 0 $X=344870 $Y=45470
X11148 2 digital_ldo_top_VIA10 $T=345340 49780 0 0 $X=344870 $Y=49550
X11149 2 digital_ldo_top_VIA10 $T=345340 53860 0 0 $X=344870 $Y=53630
X11150 2 digital_ldo_top_VIA10 $T=345340 57940 0 0 $X=344870 $Y=57710
X11151 2 digital_ldo_top_VIA10 $T=345340 62020 0 0 $X=344870 $Y=61790
X11152 2 digital_ldo_top_VIA10 $T=345340 66100 0 0 $X=344870 $Y=65870
X11153 2 digital_ldo_top_VIA10 $T=345340 70180 0 0 $X=344870 $Y=69950
X11154 2 digital_ldo_top_VIA10 $T=345340 74260 0 0 $X=344870 $Y=74030
X11155 2 digital_ldo_top_VIA10 $T=345340 78340 0 0 $X=344870 $Y=78110
X11156 2 digital_ldo_top_VIA10 $T=345340 82420 0 0 $X=344870 $Y=82190
X11157 2 digital_ldo_top_VIA10 $T=345340 86500 0 0 $X=344870 $Y=86270
X11158 2 digital_ldo_top_VIA10 $T=345340 90580 0 0 $X=344870 $Y=90350
X11159 2 digital_ldo_top_VIA10 $T=345340 94660 0 0 $X=344870 $Y=94430
X11160 2 digital_ldo_top_VIA10 $T=345340 98740 0 0 $X=344870 $Y=98510
X11161 2 digital_ldo_top_VIA10 $T=345340 102820 0 0 $X=344870 $Y=102590
X11162 2 digital_ldo_top_VIA10 $T=345340 106900 0 0 $X=344870 $Y=106670
X11163 2 digital_ldo_top_VIA10 $T=345340 110980 0 0 $X=344870 $Y=110750
X11164 2 digital_ldo_top_VIA10 $T=345340 115060 0 0 $X=344870 $Y=114830
X11165 2 digital_ldo_top_VIA10 $T=345340 119140 0 0 $X=344870 $Y=118910
X11166 2 digital_ldo_top_VIA10 $T=345340 123220 0 0 $X=344870 $Y=122990
X11167 2 digital_ldo_top_VIA10 $T=345340 127300 0 0 $X=344870 $Y=127070
X11168 3 digital_ldo_top_VIA10 $T=349020 11700 0 0 $X=348550 $Y=11470
X11169 3 digital_ldo_top_VIA10 $T=349020 15780 0 0 $X=348550 $Y=15550
X11170 3 digital_ldo_top_VIA10 $T=349020 19860 0 0 $X=348550 $Y=19630
X11171 3 digital_ldo_top_VIA10 $T=349020 23940 0 0 $X=348550 $Y=23710
X11172 3 digital_ldo_top_VIA10 $T=349020 28020 0 0 $X=348550 $Y=27790
X11173 3 digital_ldo_top_VIA10 $T=349020 32100 0 0 $X=348550 $Y=31870
X11174 3 digital_ldo_top_VIA10 $T=349020 36180 0 0 $X=348550 $Y=35950
X11175 3 digital_ldo_top_VIA10 $T=349020 40260 0 0 $X=348550 $Y=40030
X11176 3 digital_ldo_top_VIA10 $T=349020 44340 0 0 $X=348550 $Y=44110
X11177 3 digital_ldo_top_VIA10 $T=349020 48420 0 0 $X=348550 $Y=48190
X11178 3 digital_ldo_top_VIA10 $T=349020 52500 0 0 $X=348550 $Y=52270
X11179 3 digital_ldo_top_VIA10 $T=349020 56580 0 0 $X=348550 $Y=56350
X11180 3 digital_ldo_top_VIA10 $T=349020 60660 0 0 $X=348550 $Y=60430
X11181 3 digital_ldo_top_VIA10 $T=349020 64740 0 0 $X=348550 $Y=64510
X11182 3 digital_ldo_top_VIA10 $T=349020 68820 0 0 $X=348550 $Y=68590
X11183 3 digital_ldo_top_VIA10 $T=349020 72900 0 0 $X=348550 $Y=72670
X11184 3 digital_ldo_top_VIA10 $T=349020 76980 0 0 $X=348550 $Y=76750
X11185 3 digital_ldo_top_VIA10 $T=349020 81060 0 0 $X=348550 $Y=80830
X11186 3 digital_ldo_top_VIA10 $T=349020 85140 0 0 $X=348550 $Y=84910
X11187 3 digital_ldo_top_VIA10 $T=349020 89220 0 0 $X=348550 $Y=88990
X11188 3 digital_ldo_top_VIA10 $T=349020 93300 0 0 $X=348550 $Y=93070
X11189 3 digital_ldo_top_VIA10 $T=349020 97380 0 0 $X=348550 $Y=97150
X11190 3 digital_ldo_top_VIA10 $T=349020 101460 0 0 $X=348550 $Y=101230
X11191 3 digital_ldo_top_VIA10 $T=349020 105540 0 0 $X=348550 $Y=105310
X11192 3 digital_ldo_top_VIA10 $T=349020 109620 0 0 $X=348550 $Y=109390
X11193 3 digital_ldo_top_VIA10 $T=349020 113700 0 0 $X=348550 $Y=113470
X11194 3 digital_ldo_top_VIA10 $T=349020 117780 0 0 $X=348550 $Y=117550
X11195 3 digital_ldo_top_VIA10 $T=349020 121860 0 0 $X=348550 $Y=121630
X11196 3 digital_ldo_top_VIA10 $T=349020 125940 0 0 $X=348550 $Y=125710
X11197 2 digital_ldo_top_VIA10 $T=350860 13060 0 0 $X=350390 $Y=12830
X11198 2 digital_ldo_top_VIA10 $T=350860 17140 0 0 $X=350390 $Y=16910
X11199 2 digital_ldo_top_VIA10 $T=350860 21220 0 0 $X=350390 $Y=20990
X11200 2 digital_ldo_top_VIA10 $T=350860 25300 0 0 $X=350390 $Y=25070
X11201 2 digital_ldo_top_VIA10 $T=350860 29380 0 0 $X=350390 $Y=29150
X11202 2 digital_ldo_top_VIA10 $T=350860 33460 0 0 $X=350390 $Y=33230
X11203 2 digital_ldo_top_VIA10 $T=350860 37540 0 0 $X=350390 $Y=37310
X11204 2 digital_ldo_top_VIA10 $T=350860 41620 0 0 $X=350390 $Y=41390
X11205 2 digital_ldo_top_VIA10 $T=350860 45700 0 0 $X=350390 $Y=45470
X11206 2 digital_ldo_top_VIA10 $T=350860 49780 0 0 $X=350390 $Y=49550
X11207 2 digital_ldo_top_VIA10 $T=350860 53860 0 0 $X=350390 $Y=53630
X11208 2 digital_ldo_top_VIA10 $T=350860 57940 0 0 $X=350390 $Y=57710
X11209 2 digital_ldo_top_VIA10 $T=350860 62020 0 0 $X=350390 $Y=61790
X11210 2 digital_ldo_top_VIA10 $T=350860 66100 0 0 $X=350390 $Y=65870
X11211 2 digital_ldo_top_VIA10 $T=350860 70180 0 0 $X=350390 $Y=69950
X11212 2 digital_ldo_top_VIA10 $T=350860 74260 0 0 $X=350390 $Y=74030
X11213 2 digital_ldo_top_VIA10 $T=350860 78340 0 0 $X=350390 $Y=78110
X11214 2 digital_ldo_top_VIA10 $T=350860 82420 0 0 $X=350390 $Y=82190
X11215 2 digital_ldo_top_VIA10 $T=350860 86500 0 0 $X=350390 $Y=86270
X11216 2 digital_ldo_top_VIA10 $T=350860 90580 0 0 $X=350390 $Y=90350
X11217 2 digital_ldo_top_VIA10 $T=350860 94660 0 0 $X=350390 $Y=94430
X11218 2 digital_ldo_top_VIA10 $T=350860 98740 0 0 $X=350390 $Y=98510
X11219 2 digital_ldo_top_VIA10 $T=350860 102820 0 0 $X=350390 $Y=102590
X11220 2 digital_ldo_top_VIA10 $T=350860 106900 0 0 $X=350390 $Y=106670
X11221 2 digital_ldo_top_VIA10 $T=350860 110980 0 0 $X=350390 $Y=110750
X11222 2 digital_ldo_top_VIA10 $T=350860 115060 0 0 $X=350390 $Y=114830
X11223 2 digital_ldo_top_VIA10 $T=350860 119140 0 0 $X=350390 $Y=118910
X11224 2 digital_ldo_top_VIA10 $T=350860 123220 0 0 $X=350390 $Y=122990
X11225 2 digital_ldo_top_VIA10 $T=350860 127300 0 0 $X=350390 $Y=127070
X11226 3 digital_ldo_top_VIA10 $T=354540 11700 0 0 $X=354070 $Y=11470
X11227 3 digital_ldo_top_VIA10 $T=354540 15780 0 0 $X=354070 $Y=15550
X11228 3 digital_ldo_top_VIA10 $T=354540 19860 0 0 $X=354070 $Y=19630
X11229 3 digital_ldo_top_VIA10 $T=354540 23940 0 0 $X=354070 $Y=23710
X11230 3 digital_ldo_top_VIA10 $T=354540 28020 0 0 $X=354070 $Y=27790
X11231 3 digital_ldo_top_VIA10 $T=354540 32100 0 0 $X=354070 $Y=31870
X11232 3 digital_ldo_top_VIA10 $T=354540 36180 0 0 $X=354070 $Y=35950
X11233 3 digital_ldo_top_VIA10 $T=354540 40260 0 0 $X=354070 $Y=40030
X11234 3 digital_ldo_top_VIA10 $T=354540 44340 0 0 $X=354070 $Y=44110
X11235 3 digital_ldo_top_VIA10 $T=354540 48420 0 0 $X=354070 $Y=48190
X11236 3 digital_ldo_top_VIA10 $T=354540 52500 0 0 $X=354070 $Y=52270
X11237 3 digital_ldo_top_VIA10 $T=354540 56580 0 0 $X=354070 $Y=56350
X11238 3 digital_ldo_top_VIA10 $T=354540 60660 0 0 $X=354070 $Y=60430
X11239 3 digital_ldo_top_VIA10 $T=354540 64740 0 0 $X=354070 $Y=64510
X11240 3 digital_ldo_top_VIA10 $T=354540 68820 0 0 $X=354070 $Y=68590
X11241 3 digital_ldo_top_VIA10 $T=354540 72900 0 0 $X=354070 $Y=72670
X11242 3 digital_ldo_top_VIA10 $T=354540 76980 0 0 $X=354070 $Y=76750
X11243 3 digital_ldo_top_VIA10 $T=354540 81060 0 0 $X=354070 $Y=80830
X11244 3 digital_ldo_top_VIA10 $T=354540 85140 0 0 $X=354070 $Y=84910
X11245 3 digital_ldo_top_VIA10 $T=354540 89220 0 0 $X=354070 $Y=88990
X11246 3 digital_ldo_top_VIA10 $T=354540 93300 0 0 $X=354070 $Y=93070
X11247 3 digital_ldo_top_VIA10 $T=354540 97380 0 0 $X=354070 $Y=97150
X11248 3 digital_ldo_top_VIA10 $T=354540 101460 0 0 $X=354070 $Y=101230
X11249 3 digital_ldo_top_VIA10 $T=354540 105540 0 0 $X=354070 $Y=105310
X11250 3 digital_ldo_top_VIA10 $T=354540 109620 0 0 $X=354070 $Y=109390
X11251 3 digital_ldo_top_VIA10 $T=354540 113700 0 0 $X=354070 $Y=113470
X11252 3 digital_ldo_top_VIA10 $T=354540 117780 0 0 $X=354070 $Y=117550
X11253 3 digital_ldo_top_VIA10 $T=354540 121860 0 0 $X=354070 $Y=121630
X11254 3 digital_ldo_top_VIA10 $T=354540 125940 0 0 $X=354070 $Y=125710
X11255 2 digital_ldo_top_VIA10 $T=356380 13060 0 0 $X=355910 $Y=12830
X11256 2 digital_ldo_top_VIA10 $T=356380 17140 0 0 $X=355910 $Y=16910
X11257 2 digital_ldo_top_VIA10 $T=356380 21220 0 0 $X=355910 $Y=20990
X11258 2 digital_ldo_top_VIA10 $T=356380 25300 0 0 $X=355910 $Y=25070
X11259 2 digital_ldo_top_VIA10 $T=356380 29380 0 0 $X=355910 $Y=29150
X11260 2 digital_ldo_top_VIA10 $T=356380 33460 0 0 $X=355910 $Y=33230
X11261 2 digital_ldo_top_VIA10 $T=356380 37540 0 0 $X=355910 $Y=37310
X11262 2 digital_ldo_top_VIA10 $T=356380 41620 0 0 $X=355910 $Y=41390
X11263 2 digital_ldo_top_VIA10 $T=356380 45700 0 0 $X=355910 $Y=45470
X11264 2 digital_ldo_top_VIA10 $T=356380 49780 0 0 $X=355910 $Y=49550
X11265 2 digital_ldo_top_VIA10 $T=356380 53860 0 0 $X=355910 $Y=53630
X11266 2 digital_ldo_top_VIA10 $T=356380 57940 0 0 $X=355910 $Y=57710
X11267 2 digital_ldo_top_VIA10 $T=356380 62020 0 0 $X=355910 $Y=61790
X11268 2 digital_ldo_top_VIA10 $T=356380 66100 0 0 $X=355910 $Y=65870
X11269 2 digital_ldo_top_VIA10 $T=356380 70180 0 0 $X=355910 $Y=69950
X11270 2 digital_ldo_top_VIA10 $T=356380 74260 0 0 $X=355910 $Y=74030
X11271 2 digital_ldo_top_VIA10 $T=356380 78340 0 0 $X=355910 $Y=78110
X11272 2 digital_ldo_top_VIA10 $T=356380 82420 0 0 $X=355910 $Y=82190
X11273 2 digital_ldo_top_VIA10 $T=356380 86500 0 0 $X=355910 $Y=86270
X11274 2 digital_ldo_top_VIA10 $T=356380 90580 0 0 $X=355910 $Y=90350
X11275 2 digital_ldo_top_VIA10 $T=356380 94660 0 0 $X=355910 $Y=94430
X11276 2 digital_ldo_top_VIA10 $T=356380 98740 0 0 $X=355910 $Y=98510
X11277 2 digital_ldo_top_VIA10 $T=356380 102820 0 0 $X=355910 $Y=102590
X11278 2 digital_ldo_top_VIA10 $T=356380 106900 0 0 $X=355910 $Y=106670
X11279 2 digital_ldo_top_VIA10 $T=356380 110980 0 0 $X=355910 $Y=110750
X11280 2 digital_ldo_top_VIA10 $T=356380 115060 0 0 $X=355910 $Y=114830
X11281 2 digital_ldo_top_VIA10 $T=356380 119140 0 0 $X=355910 $Y=118910
X11282 2 digital_ldo_top_VIA10 $T=356380 123220 0 0 $X=355910 $Y=122990
X11283 2 digital_ldo_top_VIA10 $T=356380 127300 0 0 $X=355910 $Y=127070
X11284 3 digital_ldo_top_VIA10 $T=360060 11700 0 0 $X=359590 $Y=11470
X11285 3 digital_ldo_top_VIA10 $T=360060 15780 0 0 $X=359590 $Y=15550
X11286 3 digital_ldo_top_VIA10 $T=360060 19860 0 0 $X=359590 $Y=19630
X11287 3 digital_ldo_top_VIA10 $T=360060 23940 0 0 $X=359590 $Y=23710
X11288 3 digital_ldo_top_VIA10 $T=360060 28020 0 0 $X=359590 $Y=27790
X11289 3 digital_ldo_top_VIA10 $T=360060 32100 0 0 $X=359590 $Y=31870
X11290 3 digital_ldo_top_VIA10 $T=360060 36180 0 0 $X=359590 $Y=35950
X11291 3 digital_ldo_top_VIA10 $T=360060 40260 0 0 $X=359590 $Y=40030
X11292 3 digital_ldo_top_VIA10 $T=360060 44340 0 0 $X=359590 $Y=44110
X11293 3 digital_ldo_top_VIA10 $T=360060 48420 0 0 $X=359590 $Y=48190
X11294 3 digital_ldo_top_VIA10 $T=360060 52500 0 0 $X=359590 $Y=52270
X11295 3 digital_ldo_top_VIA10 $T=360060 56580 0 0 $X=359590 $Y=56350
X11296 3 digital_ldo_top_VIA10 $T=360060 60660 0 0 $X=359590 $Y=60430
X11297 3 digital_ldo_top_VIA10 $T=360060 64740 0 0 $X=359590 $Y=64510
X11298 3 digital_ldo_top_VIA10 $T=360060 68820 0 0 $X=359590 $Y=68590
X11299 3 digital_ldo_top_VIA10 $T=360060 72900 0 0 $X=359590 $Y=72670
X11300 3 digital_ldo_top_VIA10 $T=360060 76980 0 0 $X=359590 $Y=76750
X11301 3 digital_ldo_top_VIA10 $T=360060 81060 0 0 $X=359590 $Y=80830
X11302 3 digital_ldo_top_VIA10 $T=360060 85140 0 0 $X=359590 $Y=84910
X11303 3 digital_ldo_top_VIA10 $T=360060 89220 0 0 $X=359590 $Y=88990
X11304 3 digital_ldo_top_VIA10 $T=360060 93300 0 0 $X=359590 $Y=93070
X11305 3 digital_ldo_top_VIA10 $T=360060 97380 0 0 $X=359590 $Y=97150
X11306 3 digital_ldo_top_VIA10 $T=360060 101460 0 0 $X=359590 $Y=101230
X11307 3 digital_ldo_top_VIA10 $T=360060 105540 0 0 $X=359590 $Y=105310
X11308 3 digital_ldo_top_VIA10 $T=360060 109620 0 0 $X=359590 $Y=109390
X11309 3 digital_ldo_top_VIA10 $T=360060 113700 0 0 $X=359590 $Y=113470
X11310 3 digital_ldo_top_VIA10 $T=360060 117780 0 0 $X=359590 $Y=117550
X11311 3 digital_ldo_top_VIA10 $T=360060 121860 0 0 $X=359590 $Y=121630
X11312 3 digital_ldo_top_VIA10 $T=360060 125940 0 0 $X=359590 $Y=125710
X11313 2 digital_ldo_top_VIA10 $T=361900 13060 0 0 $X=361430 $Y=12830
X11314 2 digital_ldo_top_VIA10 $T=361900 17140 0 0 $X=361430 $Y=16910
X11315 2 digital_ldo_top_VIA10 $T=361900 21220 0 0 $X=361430 $Y=20990
X11316 2 digital_ldo_top_VIA10 $T=361900 25300 0 0 $X=361430 $Y=25070
X11317 2 digital_ldo_top_VIA10 $T=361900 29380 0 0 $X=361430 $Y=29150
X11318 2 digital_ldo_top_VIA10 $T=361900 33460 0 0 $X=361430 $Y=33230
X11319 2 digital_ldo_top_VIA10 $T=361900 37540 0 0 $X=361430 $Y=37310
X11320 2 digital_ldo_top_VIA10 $T=361900 41620 0 0 $X=361430 $Y=41390
X11321 2 digital_ldo_top_VIA10 $T=361900 45700 0 0 $X=361430 $Y=45470
X11322 2 digital_ldo_top_VIA10 $T=361900 49780 0 0 $X=361430 $Y=49550
X11323 2 digital_ldo_top_VIA10 $T=361900 53860 0 0 $X=361430 $Y=53630
X11324 2 digital_ldo_top_VIA10 $T=361900 57940 0 0 $X=361430 $Y=57710
X11325 2 digital_ldo_top_VIA10 $T=361900 62020 0 0 $X=361430 $Y=61790
X11326 2 digital_ldo_top_VIA10 $T=361900 66100 0 0 $X=361430 $Y=65870
X11327 2 digital_ldo_top_VIA10 $T=361900 70180 0 0 $X=361430 $Y=69950
X11328 2 digital_ldo_top_VIA10 $T=361900 74260 0 0 $X=361430 $Y=74030
X11329 2 digital_ldo_top_VIA10 $T=361900 78340 0 0 $X=361430 $Y=78110
X11330 2 digital_ldo_top_VIA10 $T=361900 82420 0 0 $X=361430 $Y=82190
X11331 2 digital_ldo_top_VIA10 $T=361900 86500 0 0 $X=361430 $Y=86270
X11332 2 digital_ldo_top_VIA10 $T=361900 90580 0 0 $X=361430 $Y=90350
X11333 2 digital_ldo_top_VIA10 $T=361900 94660 0 0 $X=361430 $Y=94430
X11334 2 digital_ldo_top_VIA10 $T=361900 98740 0 0 $X=361430 $Y=98510
X11335 2 digital_ldo_top_VIA10 $T=361900 102820 0 0 $X=361430 $Y=102590
X11336 2 digital_ldo_top_VIA10 $T=361900 106900 0 0 $X=361430 $Y=106670
X11337 2 digital_ldo_top_VIA10 $T=361900 110980 0 0 $X=361430 $Y=110750
X11338 2 digital_ldo_top_VIA10 $T=361900 115060 0 0 $X=361430 $Y=114830
X11339 2 digital_ldo_top_VIA10 $T=361900 119140 0 0 $X=361430 $Y=118910
X11340 2 digital_ldo_top_VIA10 $T=361900 123220 0 0 $X=361430 $Y=122990
X11341 2 digital_ldo_top_VIA10 $T=361900 127300 0 0 $X=361430 $Y=127070
X11342 3 digital_ldo_top_VIA10 $T=365580 11700 0 0 $X=365110 $Y=11470
X11343 3 digital_ldo_top_VIA10 $T=365580 15780 0 0 $X=365110 $Y=15550
X11344 3 digital_ldo_top_VIA10 $T=365580 19860 0 0 $X=365110 $Y=19630
X11345 3 digital_ldo_top_VIA10 $T=365580 23940 0 0 $X=365110 $Y=23710
X11346 3 digital_ldo_top_VIA10 $T=365580 28020 0 0 $X=365110 $Y=27790
X11347 3 digital_ldo_top_VIA10 $T=365580 32100 0 0 $X=365110 $Y=31870
X11348 3 digital_ldo_top_VIA10 $T=365580 36180 0 0 $X=365110 $Y=35950
X11349 3 digital_ldo_top_VIA10 $T=365580 40260 0 0 $X=365110 $Y=40030
X11350 3 digital_ldo_top_VIA10 $T=365580 44340 0 0 $X=365110 $Y=44110
X11351 3 digital_ldo_top_VIA10 $T=365580 48420 0 0 $X=365110 $Y=48190
X11352 3 digital_ldo_top_VIA10 $T=365580 52500 0 0 $X=365110 $Y=52270
X11353 3 digital_ldo_top_VIA10 $T=365580 56580 0 0 $X=365110 $Y=56350
X11354 3 digital_ldo_top_VIA10 $T=365580 60660 0 0 $X=365110 $Y=60430
X11355 3 digital_ldo_top_VIA10 $T=365580 64740 0 0 $X=365110 $Y=64510
X11356 3 digital_ldo_top_VIA10 $T=365580 68820 0 0 $X=365110 $Y=68590
X11357 3 digital_ldo_top_VIA10 $T=365580 72900 0 0 $X=365110 $Y=72670
X11358 3 digital_ldo_top_VIA10 $T=365580 76980 0 0 $X=365110 $Y=76750
X11359 3 digital_ldo_top_VIA10 $T=365580 81060 0 0 $X=365110 $Y=80830
X11360 3 digital_ldo_top_VIA10 $T=365580 85140 0 0 $X=365110 $Y=84910
X11361 3 digital_ldo_top_VIA10 $T=365580 89220 0 0 $X=365110 $Y=88990
X11362 3 digital_ldo_top_VIA10 $T=365580 93300 0 0 $X=365110 $Y=93070
X11363 3 digital_ldo_top_VIA10 $T=365580 97380 0 0 $X=365110 $Y=97150
X11364 3 digital_ldo_top_VIA10 $T=365580 101460 0 0 $X=365110 $Y=101230
X11365 3 digital_ldo_top_VIA10 $T=365580 105540 0 0 $X=365110 $Y=105310
X11366 3 digital_ldo_top_VIA10 $T=365580 109620 0 0 $X=365110 $Y=109390
X11367 3 digital_ldo_top_VIA10 $T=365580 113700 0 0 $X=365110 $Y=113470
X11368 3 digital_ldo_top_VIA10 $T=365580 117780 0 0 $X=365110 $Y=117550
X11369 3 digital_ldo_top_VIA10 $T=365580 121860 0 0 $X=365110 $Y=121630
X11370 3 digital_ldo_top_VIA10 $T=365580 125940 0 0 $X=365110 $Y=125710
X11371 2 digital_ldo_top_VIA10 $T=367420 13060 0 0 $X=366950 $Y=12830
X11372 2 digital_ldo_top_VIA10 $T=367420 17140 0 0 $X=366950 $Y=16910
X11373 2 digital_ldo_top_VIA10 $T=367420 21220 0 0 $X=366950 $Y=20990
X11374 2 digital_ldo_top_VIA10 $T=367420 25300 0 0 $X=366950 $Y=25070
X11375 2 digital_ldo_top_VIA10 $T=367420 29380 0 0 $X=366950 $Y=29150
X11376 2 digital_ldo_top_VIA10 $T=367420 33460 0 0 $X=366950 $Y=33230
X11377 2 digital_ldo_top_VIA10 $T=367420 37540 0 0 $X=366950 $Y=37310
X11378 2 digital_ldo_top_VIA10 $T=367420 41620 0 0 $X=366950 $Y=41390
X11379 2 digital_ldo_top_VIA10 $T=367420 45700 0 0 $X=366950 $Y=45470
X11380 2 digital_ldo_top_VIA10 $T=367420 49780 0 0 $X=366950 $Y=49550
X11381 2 digital_ldo_top_VIA10 $T=367420 53860 0 0 $X=366950 $Y=53630
X11382 2 digital_ldo_top_VIA10 $T=367420 57940 0 0 $X=366950 $Y=57710
X11383 2 digital_ldo_top_VIA10 $T=367420 62020 0 0 $X=366950 $Y=61790
X11384 2 digital_ldo_top_VIA10 $T=367420 66100 0 0 $X=366950 $Y=65870
X11385 2 digital_ldo_top_VIA10 $T=367420 70180 0 0 $X=366950 $Y=69950
X11386 2 digital_ldo_top_VIA10 $T=367420 74260 0 0 $X=366950 $Y=74030
X11387 2 digital_ldo_top_VIA10 $T=367420 78340 0 0 $X=366950 $Y=78110
X11388 2 digital_ldo_top_VIA10 $T=367420 82420 0 0 $X=366950 $Y=82190
X11389 2 digital_ldo_top_VIA10 $T=367420 86500 0 0 $X=366950 $Y=86270
X11390 2 digital_ldo_top_VIA10 $T=367420 90580 0 0 $X=366950 $Y=90350
X11391 2 digital_ldo_top_VIA10 $T=367420 94660 0 0 $X=366950 $Y=94430
X11392 2 digital_ldo_top_VIA10 $T=367420 98740 0 0 $X=366950 $Y=98510
X11393 2 digital_ldo_top_VIA10 $T=367420 102820 0 0 $X=366950 $Y=102590
X11394 2 digital_ldo_top_VIA10 $T=367420 106900 0 0 $X=366950 $Y=106670
X11395 2 digital_ldo_top_VIA10 $T=367420 110980 0 0 $X=366950 $Y=110750
X11396 2 digital_ldo_top_VIA10 $T=367420 115060 0 0 $X=366950 $Y=114830
X11397 2 digital_ldo_top_VIA10 $T=367420 119140 0 0 $X=366950 $Y=118910
X11398 2 digital_ldo_top_VIA10 $T=367420 123220 0 0 $X=366950 $Y=122990
X11399 2 digital_ldo_top_VIA10 $T=367420 127300 0 0 $X=366950 $Y=127070
X11400 3 digital_ldo_top_VIA10 $T=371100 11700 0 0 $X=370630 $Y=11470
X11401 3 digital_ldo_top_VIA10 $T=371100 15780 0 0 $X=370630 $Y=15550
X11402 3 digital_ldo_top_VIA10 $T=371100 19860 0 0 $X=370630 $Y=19630
X11403 3 digital_ldo_top_VIA10 $T=371100 23940 0 0 $X=370630 $Y=23710
X11404 3 digital_ldo_top_VIA10 $T=371100 28020 0 0 $X=370630 $Y=27790
X11405 3 digital_ldo_top_VIA10 $T=371100 32100 0 0 $X=370630 $Y=31870
X11406 3 digital_ldo_top_VIA10 $T=371100 36180 0 0 $X=370630 $Y=35950
X11407 3 digital_ldo_top_VIA10 $T=371100 40260 0 0 $X=370630 $Y=40030
X11408 3 digital_ldo_top_VIA10 $T=371100 44340 0 0 $X=370630 $Y=44110
X11409 3 digital_ldo_top_VIA10 $T=371100 48420 0 0 $X=370630 $Y=48190
X11410 3 digital_ldo_top_VIA10 $T=371100 52500 0 0 $X=370630 $Y=52270
X11411 3 digital_ldo_top_VIA10 $T=371100 56580 0 0 $X=370630 $Y=56350
X11412 3 digital_ldo_top_VIA10 $T=371100 60660 0 0 $X=370630 $Y=60430
X11413 3 digital_ldo_top_VIA10 $T=371100 64740 0 0 $X=370630 $Y=64510
X11414 3 digital_ldo_top_VIA10 $T=371100 68820 0 0 $X=370630 $Y=68590
X11415 3 digital_ldo_top_VIA10 $T=371100 72900 0 0 $X=370630 $Y=72670
X11416 3 digital_ldo_top_VIA10 $T=371100 76980 0 0 $X=370630 $Y=76750
X11417 3 digital_ldo_top_VIA10 $T=371100 81060 0 0 $X=370630 $Y=80830
X11418 3 digital_ldo_top_VIA10 $T=371100 85140 0 0 $X=370630 $Y=84910
X11419 3 digital_ldo_top_VIA10 $T=371100 89220 0 0 $X=370630 $Y=88990
X11420 3 digital_ldo_top_VIA10 $T=371100 93300 0 0 $X=370630 $Y=93070
X11421 3 digital_ldo_top_VIA10 $T=371100 97380 0 0 $X=370630 $Y=97150
X11422 3 digital_ldo_top_VIA10 $T=371100 101460 0 0 $X=370630 $Y=101230
X11423 3 digital_ldo_top_VIA10 $T=371100 105540 0 0 $X=370630 $Y=105310
X11424 3 digital_ldo_top_VIA10 $T=371100 109620 0 0 $X=370630 $Y=109390
X11425 3 digital_ldo_top_VIA10 $T=371100 113700 0 0 $X=370630 $Y=113470
X11426 3 digital_ldo_top_VIA10 $T=371100 117780 0 0 $X=370630 $Y=117550
X11427 3 digital_ldo_top_VIA10 $T=371100 121860 0 0 $X=370630 $Y=121630
X11428 3 digital_ldo_top_VIA10 $T=371100 125940 0 0 $X=370630 $Y=125710
X11429 2 digital_ldo_top_VIA10 $T=372940 13060 0 0 $X=372470 $Y=12830
X11430 2 digital_ldo_top_VIA10 $T=372940 17140 0 0 $X=372470 $Y=16910
X11431 2 digital_ldo_top_VIA10 $T=372940 21220 0 0 $X=372470 $Y=20990
X11432 2 digital_ldo_top_VIA10 $T=372940 25300 0 0 $X=372470 $Y=25070
X11433 2 digital_ldo_top_VIA10 $T=372940 29380 0 0 $X=372470 $Y=29150
X11434 2 digital_ldo_top_VIA10 $T=372940 33460 0 0 $X=372470 $Y=33230
X11435 2 digital_ldo_top_VIA10 $T=372940 37540 0 0 $X=372470 $Y=37310
X11436 2 digital_ldo_top_VIA10 $T=372940 41620 0 0 $X=372470 $Y=41390
X11437 2 digital_ldo_top_VIA10 $T=372940 45700 0 0 $X=372470 $Y=45470
X11438 2 digital_ldo_top_VIA10 $T=372940 49780 0 0 $X=372470 $Y=49550
X11439 2 digital_ldo_top_VIA10 $T=372940 53860 0 0 $X=372470 $Y=53630
X11440 2 digital_ldo_top_VIA10 $T=372940 57940 0 0 $X=372470 $Y=57710
X11441 2 digital_ldo_top_VIA10 $T=372940 62020 0 0 $X=372470 $Y=61790
X11442 2 digital_ldo_top_VIA10 $T=372940 66100 0 0 $X=372470 $Y=65870
X11443 2 digital_ldo_top_VIA10 $T=372940 70180 0 0 $X=372470 $Y=69950
X11444 2 digital_ldo_top_VIA10 $T=372940 74260 0 0 $X=372470 $Y=74030
X11445 2 digital_ldo_top_VIA10 $T=372940 78340 0 0 $X=372470 $Y=78110
X11446 2 digital_ldo_top_VIA10 $T=372940 82420 0 0 $X=372470 $Y=82190
X11447 2 digital_ldo_top_VIA10 $T=372940 86500 0 0 $X=372470 $Y=86270
X11448 2 digital_ldo_top_VIA10 $T=372940 90580 0 0 $X=372470 $Y=90350
X11449 2 digital_ldo_top_VIA10 $T=372940 94660 0 0 $X=372470 $Y=94430
X11450 2 digital_ldo_top_VIA10 $T=372940 98740 0 0 $X=372470 $Y=98510
X11451 2 digital_ldo_top_VIA10 $T=372940 102820 0 0 $X=372470 $Y=102590
X11452 2 digital_ldo_top_VIA10 $T=372940 106900 0 0 $X=372470 $Y=106670
X11453 2 digital_ldo_top_VIA10 $T=372940 110980 0 0 $X=372470 $Y=110750
X11454 2 digital_ldo_top_VIA10 $T=372940 115060 0 0 $X=372470 $Y=114830
X11455 2 digital_ldo_top_VIA10 $T=372940 119140 0 0 $X=372470 $Y=118910
X11456 2 digital_ldo_top_VIA10 $T=372940 123220 0 0 $X=372470 $Y=122990
X11457 2 digital_ldo_top_VIA10 $T=372940 127300 0 0 $X=372470 $Y=127070
X11458 3 digital_ldo_top_VIA10 $T=376620 11700 0 0 $X=376150 $Y=11470
X11459 3 digital_ldo_top_VIA10 $T=376620 15780 0 0 $X=376150 $Y=15550
X11460 3 digital_ldo_top_VIA10 $T=376620 19860 0 0 $X=376150 $Y=19630
X11461 3 digital_ldo_top_VIA10 $T=376620 23940 0 0 $X=376150 $Y=23710
X11462 3 digital_ldo_top_VIA10 $T=376620 28020 0 0 $X=376150 $Y=27790
X11463 3 digital_ldo_top_VIA10 $T=376620 32100 0 0 $X=376150 $Y=31870
X11464 3 digital_ldo_top_VIA10 $T=376620 36180 0 0 $X=376150 $Y=35950
X11465 3 digital_ldo_top_VIA10 $T=376620 40260 0 0 $X=376150 $Y=40030
X11466 3 digital_ldo_top_VIA10 $T=376620 44340 0 0 $X=376150 $Y=44110
X11467 3 digital_ldo_top_VIA10 $T=376620 48420 0 0 $X=376150 $Y=48190
X11468 3 digital_ldo_top_VIA10 $T=376620 52500 0 0 $X=376150 $Y=52270
X11469 3 digital_ldo_top_VIA10 $T=376620 56580 0 0 $X=376150 $Y=56350
X11470 3 digital_ldo_top_VIA10 $T=376620 60660 0 0 $X=376150 $Y=60430
X11471 3 digital_ldo_top_VIA10 $T=376620 64740 0 0 $X=376150 $Y=64510
X11472 3 digital_ldo_top_VIA10 $T=376620 68820 0 0 $X=376150 $Y=68590
X11473 3 digital_ldo_top_VIA10 $T=376620 72900 0 0 $X=376150 $Y=72670
X11474 3 digital_ldo_top_VIA10 $T=376620 76980 0 0 $X=376150 $Y=76750
X11475 3 digital_ldo_top_VIA10 $T=376620 81060 0 0 $X=376150 $Y=80830
X11476 3 digital_ldo_top_VIA10 $T=376620 85140 0 0 $X=376150 $Y=84910
X11477 3 digital_ldo_top_VIA10 $T=376620 89220 0 0 $X=376150 $Y=88990
X11478 3 digital_ldo_top_VIA10 $T=376620 93300 0 0 $X=376150 $Y=93070
X11479 3 digital_ldo_top_VIA10 $T=376620 97380 0 0 $X=376150 $Y=97150
X11480 3 digital_ldo_top_VIA10 $T=376620 101460 0 0 $X=376150 $Y=101230
X11481 3 digital_ldo_top_VIA10 $T=376620 105540 0 0 $X=376150 $Y=105310
X11482 3 digital_ldo_top_VIA10 $T=376620 109620 0 0 $X=376150 $Y=109390
X11483 3 digital_ldo_top_VIA10 $T=376620 113700 0 0 $X=376150 $Y=113470
X11484 3 digital_ldo_top_VIA10 $T=376620 117780 0 0 $X=376150 $Y=117550
X11485 3 digital_ldo_top_VIA10 $T=376620 121860 0 0 $X=376150 $Y=121630
X11486 3 digital_ldo_top_VIA10 $T=376620 125940 0 0 $X=376150 $Y=125710
X11487 2 digital_ldo_top_VIA10 $T=378460 13060 0 0 $X=377990 $Y=12830
X11488 2 digital_ldo_top_VIA10 $T=378460 17140 0 0 $X=377990 $Y=16910
X11489 2 digital_ldo_top_VIA10 $T=378460 21220 0 0 $X=377990 $Y=20990
X11490 2 digital_ldo_top_VIA10 $T=378460 25300 0 0 $X=377990 $Y=25070
X11491 2 digital_ldo_top_VIA10 $T=378460 29380 0 0 $X=377990 $Y=29150
X11492 2 digital_ldo_top_VIA10 $T=378460 33460 0 0 $X=377990 $Y=33230
X11493 2 digital_ldo_top_VIA10 $T=378460 37540 0 0 $X=377990 $Y=37310
X11494 2 digital_ldo_top_VIA10 $T=378460 41620 0 0 $X=377990 $Y=41390
X11495 2 digital_ldo_top_VIA10 $T=378460 45700 0 0 $X=377990 $Y=45470
X11496 2 digital_ldo_top_VIA10 $T=378460 49780 0 0 $X=377990 $Y=49550
X11497 2 digital_ldo_top_VIA10 $T=378460 53860 0 0 $X=377990 $Y=53630
X11498 2 digital_ldo_top_VIA10 $T=378460 57940 0 0 $X=377990 $Y=57710
X11499 2 digital_ldo_top_VIA10 $T=378460 62020 0 0 $X=377990 $Y=61790
X11500 2 digital_ldo_top_VIA10 $T=378460 66100 0 0 $X=377990 $Y=65870
X11501 2 digital_ldo_top_VIA10 $T=378460 70180 0 0 $X=377990 $Y=69950
X11502 2 digital_ldo_top_VIA10 $T=378460 74260 0 0 $X=377990 $Y=74030
X11503 2 digital_ldo_top_VIA10 $T=378460 78340 0 0 $X=377990 $Y=78110
X11504 2 digital_ldo_top_VIA10 $T=378460 82420 0 0 $X=377990 $Y=82190
X11505 2 digital_ldo_top_VIA10 $T=378460 86500 0 0 $X=377990 $Y=86270
X11506 2 digital_ldo_top_VIA10 $T=378460 90580 0 0 $X=377990 $Y=90350
X11507 2 digital_ldo_top_VIA10 $T=378460 94660 0 0 $X=377990 $Y=94430
X11508 2 digital_ldo_top_VIA10 $T=378460 98740 0 0 $X=377990 $Y=98510
X11509 2 digital_ldo_top_VIA10 $T=378460 102820 0 0 $X=377990 $Y=102590
X11510 2 digital_ldo_top_VIA10 $T=378460 106900 0 0 $X=377990 $Y=106670
X11511 2 digital_ldo_top_VIA10 $T=378460 110980 0 0 $X=377990 $Y=110750
X11512 2 digital_ldo_top_VIA10 $T=378460 115060 0 0 $X=377990 $Y=114830
X11513 2 digital_ldo_top_VIA10 $T=378460 119140 0 0 $X=377990 $Y=118910
X11514 2 digital_ldo_top_VIA10 $T=378460 123220 0 0 $X=377990 $Y=122990
X11515 2 digital_ldo_top_VIA10 $T=378460 127300 0 0 $X=377990 $Y=127070
X11516 2 digital_ldo_top_VIA11 $T=307005 29380 0 0 $X=306840 $Y=29150
X11517 2 digital_ldo_top_VIA11 $T=307005 33460 0 0 $X=306840 $Y=33230
X11518 2 digital_ldo_top_VIA11 $T=307005 37540 0 0 $X=306840 $Y=37310
X11519 2 digital_ldo_top_VIA11 $T=307005 41620 0 0 $X=306840 $Y=41390
X11520 2 digital_ldo_top_VIA11 $T=307005 45700 0 0 $X=306840 $Y=45470
X11521 2 digital_ldo_top_VIA11 $T=307005 49780 0 0 $X=306840 $Y=49550
X11522 2 digital_ldo_top_VIA11 $T=307005 53860 0 0 $X=306840 $Y=53630
X11523 2 digital_ldo_top_VIA11 $T=307005 57940 0 0 $X=306840 $Y=57710
X11524 2 digital_ldo_top_VIA11 $T=307005 62020 0 0 $X=306840 $Y=61790
X11525 2 digital_ldo_top_VIA11 $T=307005 66100 0 0 $X=306840 $Y=65870
X11526 2 digital_ldo_top_VIA11 $T=307005 70180 0 0 $X=306840 $Y=69950
X11527 2 digital_ldo_top_VIA11 $T=307005 74260 0 0 $X=306840 $Y=74030
X11528 2 digital_ldo_top_VIA11 $T=307005 78340 0 0 $X=306840 $Y=78110
X11529 2 digital_ldo_top_VIA11 $T=307005 82420 0 0 $X=306840 $Y=82190
X11530 2 digital_ldo_top_VIA12 $T=14140 45700 0 0 $X=13430 $Y=44700
X11531 2 digital_ldo_top_VIA12 $T=14140 66100 0 0 $X=13430 $Y=65100
X11532 2 digital_ldo_top_VIA12 $T=19660 45700 0 0 $X=18950 $Y=44700
X11533 2 digital_ldo_top_VIA12 $T=19660 66100 0 0 $X=18950 $Y=65100
X11534 2 digital_ldo_top_VIA12 $T=25180 45700 0 0 $X=24470 $Y=44700
X11535 2 digital_ldo_top_VIA12 $T=25180 66100 0 0 $X=24470 $Y=65100
X11536 2 digital_ldo_top_VIA12 $T=30700 45700 0 0 $X=29990 $Y=44700
X11537 2 digital_ldo_top_VIA12 $T=30700 66100 0 0 $X=29990 $Y=65100
X11538 2 digital_ldo_top_VIA12 $T=36220 45700 0 0 $X=35510 $Y=44700
X11539 2 digital_ldo_top_VIA12 $T=36220 66100 0 0 $X=35510 $Y=65100
X11540 2 digital_ldo_top_VIA12 $T=41740 45700 0 0 $X=41030 $Y=44700
X11541 2 digital_ldo_top_VIA12 $T=41740 66100 0 0 $X=41030 $Y=65100
X11542 2 digital_ldo_top_VIA12 $T=47260 45700 0 0 $X=46550 $Y=44700
X11543 2 digital_ldo_top_VIA12 $T=47260 66100 0 0 $X=46550 $Y=65100
X11544 2 digital_ldo_top_VIA12 $T=52780 45700 0 0 $X=52070 $Y=44700
X11545 2 digital_ldo_top_VIA12 $T=52780 66100 0 0 $X=52070 $Y=65100
X11546 2 digital_ldo_top_VIA12 $T=58300 45700 0 0 $X=57590 $Y=44700
X11547 2 digital_ldo_top_VIA12 $T=58300 66100 0 0 $X=57590 $Y=65100
X11548 2 digital_ldo_top_VIA12 $T=63820 45700 0 0 $X=63110 $Y=44700
X11549 2 digital_ldo_top_VIA12 $T=63820 66100 0 0 $X=63110 $Y=65100
X11550 2 digital_ldo_top_VIA12 $T=69340 45700 0 0 $X=68630 $Y=44700
X11551 2 digital_ldo_top_VIA12 $T=69340 66100 0 0 $X=68630 $Y=65100
X11552 2 digital_ldo_top_VIA12 $T=74860 45700 0 0 $X=74150 $Y=44700
X11553 2 digital_ldo_top_VIA12 $T=74860 66100 0 0 $X=74150 $Y=65100
X11554 2 digital_ldo_top_VIA12 $T=80380 25300 0 0 $X=79670 $Y=24300
X11555 2 digital_ldo_top_VIA12 $T=80380 45700 0 0 $X=79670 $Y=44700
X11556 2 digital_ldo_top_VIA12 $T=80380 66100 0 0 $X=79670 $Y=65100
X11557 2 digital_ldo_top_VIA12 $T=85900 25300 0 0 $X=85190 $Y=24300
X11558 2 digital_ldo_top_VIA12 $T=85900 45700 0 0 $X=85190 $Y=44700
X11559 2 digital_ldo_top_VIA12 $T=85900 66100 0 0 $X=85190 $Y=65100
X11560 2 digital_ldo_top_VIA12 $T=91420 25300 0 0 $X=90710 $Y=24300
X11561 2 digital_ldo_top_VIA12 $T=91420 45700 0 0 $X=90710 $Y=44700
X11562 2 digital_ldo_top_VIA12 $T=91420 66100 0 0 $X=90710 $Y=65100
X11563 2 digital_ldo_top_VIA12 $T=96940 25300 0 0 $X=96230 $Y=24300
X11564 2 digital_ldo_top_VIA12 $T=96940 45700 0 0 $X=96230 $Y=44700
X11565 2 digital_ldo_top_VIA12 $T=96940 66100 0 0 $X=96230 $Y=65100
X11566 2 digital_ldo_top_VIA12 $T=102460 25300 0 0 $X=101750 $Y=24300
X11567 2 digital_ldo_top_VIA12 $T=102460 45700 0 0 $X=101750 $Y=44700
X11568 2 digital_ldo_top_VIA12 $T=102460 66100 0 0 $X=101750 $Y=65100
X11569 2 digital_ldo_top_VIA12 $T=107980 25300 0 0 $X=107270 $Y=24300
X11570 2 digital_ldo_top_VIA12 $T=113500 25300 0 0 $X=112790 $Y=24300
X11571 2 digital_ldo_top_VIA12 $T=119020 25300 0 0 $X=118310 $Y=24300
X11572 2 digital_ldo_top_VIA12 $T=124540 25300 0 0 $X=123830 $Y=24300
X11573 2 digital_ldo_top_VIA12 $T=130060 25300 0 0 $X=129350 $Y=24300
X11574 2 digital_ldo_top_VIA12 $T=135580 25300 0 0 $X=134870 $Y=24300
X11575 2 digital_ldo_top_VIA12 $T=146620 25300 0 0 $X=145910 $Y=24300
X11576 2 digital_ldo_top_VIA12 $T=152140 25300 0 0 $X=151430 $Y=24300
X11577 2 digital_ldo_top_VIA12 $T=157660 25300 0 0 $X=156950 $Y=24300
X11578 2 digital_ldo_top_VIA12 $T=163180 25300 0 0 $X=162470 $Y=24300
X11579 2 digital_ldo_top_VIA12 $T=168700 25300 0 0 $X=167990 $Y=24300
X11580 2 digital_ldo_top_VIA12 $T=174220 25300 0 0 $X=173510 $Y=24300
X11581 2 digital_ldo_top_VIA12 $T=185260 25300 0 0 $X=184550 $Y=24300
X11582 2 digital_ldo_top_VIA12 $T=190780 25300 0 0 $X=190070 $Y=24300
X11583 2 digital_ldo_top_VIA12 $T=196300 25300 0 0 $X=195590 $Y=24300
X11584 2 digital_ldo_top_VIA12 $T=201820 25300 0 0 $X=201110 $Y=24300
X11585 2 digital_ldo_top_VIA12 $T=207340 25300 0 0 $X=206630 $Y=24300
X11586 2 digital_ldo_top_VIA12 $T=212860 25300 0 0 $X=212150 $Y=24300
X11587 2 digital_ldo_top_VIA12 $T=223900 25300 0 0 $X=223190 $Y=24300
X11588 2 digital_ldo_top_VIA12 $T=229420 25300 0 0 $X=228710 $Y=24300
X11589 2 digital_ldo_top_VIA12 $T=234940 25300 0 0 $X=234230 $Y=24300
X11590 2 digital_ldo_top_VIA12 $T=240460 25300 0 0 $X=239750 $Y=24300
X11591 2 digital_ldo_top_VIA12 $T=245980 25300 0 0 $X=245270 $Y=24300
X11592 2 digital_ldo_top_VIA12 $T=251500 25300 0 0 $X=250790 $Y=24300
X11593 2 digital_ldo_top_VIA12 $T=262540 25300 0 0 $X=261830 $Y=24300
X11594 2 digital_ldo_top_VIA12 $T=267820 25300 0 0 $X=267110 $Y=24300
X11595 2 digital_ldo_top_VIA12 $T=273580 25300 0 0 $X=272870 $Y=24300
X11596 2 digital_ldo_top_VIA12 $T=279100 25300 0 0 $X=278390 $Y=24300
X11597 2 digital_ldo_top_VIA12 $T=284620 25300 0 0 $X=283910 $Y=24300
X11598 2 digital_ldo_top_VIA12 $T=290140 25300 0 0 $X=289430 $Y=24300
X11599 2 digital_ldo_top_VIA12 $T=295900 25300 0 0 $X=295190 $Y=24300
X11600 2 digital_ldo_top_VIA12 $T=301180 25300 0 0 $X=300470 $Y=24300
X11601 2 digital_ldo_top_VIA12 $T=350860 45700 0 0 $X=350150 $Y=44700
X11602 2 digital_ldo_top_VIA12 $T=350860 66100 0 0 $X=350150 $Y=65100
X11603 2 digital_ldo_top_VIA12 $T=356380 45700 0 0 $X=355670 $Y=44700
X11604 2 digital_ldo_top_VIA12 $T=356380 66100 0 0 $X=355670 $Y=65100
X11605 2 digital_ldo_top_VIA12 $T=361900 45700 0 0 $X=361190 $Y=44700
X11606 2 digital_ldo_top_VIA12 $T=361900 66100 0 0 $X=361190 $Y=65100
X11607 2 digital_ldo_top_VIA12 $T=367420 45700 0 0 $X=366710 $Y=44700
X11608 2 digital_ldo_top_VIA12 $T=367420 66100 0 0 $X=366710 $Y=65100
X11609 2 digital_ldo_top_VIA12 $T=372940 45700 0 0 $X=372230 $Y=44700
X11610 2 digital_ldo_top_VIA12 $T=372940 66100 0 0 $X=372230 $Y=65100
X11611 2 digital_ldo_top_VIA12 $T=378460 45700 0 0 $X=377750 $Y=44700
X11612 2 digital_ldo_top_VIA12 $T=378460 66100 0 0 $X=377750 $Y=65100
X11613 2 digital_ldo_top_VIA13 $T=307710 45700 0 0 $X=307000 $Y=44700
X11614 2 digital_ldo_top_VIA13 $T=307710 66100 0 0 $X=307000 $Y=65100
X11615 3 digital_ldo_top_VIA15 $T=26795 23940 0 0 $X=26580 $Y=23710
X11616 3 digital_ldo_top_VIA15 $T=86795 23940 0 0 $X=86580 $Y=23710
X11617 3 digital_ldo_top_VIA15 $T=86795 32100 0 0 $X=86580 $Y=31870
X11618 3 digital_ldo_top_VIA15 $T=86795 36180 0 0 $X=86580 $Y=35950
X11619 3 digital_ldo_top_VIA16 $T=26795 20205 0 0 $X=26580 $Y=20040
X11620 3 digital_ldo_top_VIA16 $T=86795 20205 0 0 $X=86580 $Y=20040
X11621 3 digital_ldo_top_VIA18 $T=116150 84955 0 0 $X=115900 $Y=84790
X11622 3 digital_ldo_top_VIA18 $T=118910 84955 0 0 $X=118660 $Y=84790
X11623 3 digital_ldo_top_VIA18 $T=124430 84955 0 0 $X=124180 $Y=84790
X11624 3 digital_ldo_top_VIA18 $T=127190 84955 0 0 $X=126940 $Y=84790
X11625 3 digital_ldo_top_VIA18 $T=129950 84955 0 0 $X=129700 $Y=84790
X11626 3 digital_ldo_top_VIA18 $T=135470 84955 0 0 $X=135220 $Y=84790
X11627 3 digital_ldo_top_VIA18 $T=138230 84955 0 0 $X=137980 $Y=84790
X11628 3 digital_ldo_top_VIA18 $T=140990 84955 0 0 $X=140740 $Y=84790
X11629 3 digital_ldo_top_VIA18 $T=146510 84955 0 0 $X=146260 $Y=84790
X11630 3 digital_ldo_top_VIA18 $T=149270 84955 0 0 $X=149020 $Y=84790
X11631 3 digital_ldo_top_VIA18 $T=152030 84955 0 0 $X=151780 $Y=84790
X11632 3 digital_ldo_top_VIA18 $T=157550 84955 0 0 $X=157300 $Y=84790
X11633 3 digital_ldo_top_VIA18 $T=160310 84955 0 0 $X=160060 $Y=84790
X11634 3 digital_ldo_top_VIA18 $T=163070 84955 0 0 $X=162820 $Y=84790
X11635 3 digital_ldo_top_VIA18 $T=168590 84955 0 0 $X=168340 $Y=84790
X11636 3 digital_ldo_top_VIA18 $T=171350 84955 0 0 $X=171100 $Y=84790
X11637 3 digital_ldo_top_VIA18 $T=174110 84955 0 0 $X=173860 $Y=84790
X11638 3 digital_ldo_top_VIA18 $T=179630 84955 0 0 $X=179380 $Y=84790
X11639 3 digital_ldo_top_VIA18 $T=182390 84955 0 0 $X=182140 $Y=84790
X11640 3 digital_ldo_top_VIA18 $T=185150 84955 0 0 $X=184900 $Y=84790
X11641 3 digital_ldo_top_VIA18 $T=190670 84955 0 0 $X=190420 $Y=84790
X11642 3 digital_ldo_top_VIA18 $T=193430 84955 0 0 $X=193180 $Y=84790
X11643 3 digital_ldo_top_VIA18 $T=196190 84955 0 0 $X=195940 $Y=84790
X11644 3 digital_ldo_top_VIA18 $T=201710 84955 0 0 $X=201460 $Y=84790
X11645 3 digital_ldo_top_VIA18 $T=204470 84955 0 0 $X=204220 $Y=84790
X11646 3 digital_ldo_top_VIA18 $T=207230 84955 0 0 $X=206980 $Y=84790
X11647 3 digital_ldo_top_VIA18 $T=212750 84955 0 0 $X=212500 $Y=84790
X11648 3 digital_ldo_top_VIA18 $T=215510 84955 0 0 $X=215260 $Y=84790
X11649 3 digital_ldo_top_VIA18 $T=218270 84955 0 0 $X=218020 $Y=84790
X11650 3 digital_ldo_top_VIA18 $T=223790 84955 0 0 $X=223540 $Y=84790
X11651 3 digital_ldo_top_VIA18 $T=226550 84955 0 0 $X=226300 $Y=84790
X11652 3 digital_ldo_top_VIA18 $T=229310 84955 0 0 $X=229060 $Y=84790
X11653 3 digital_ldo_top_VIA18 $T=234830 84955 0 0 $X=234580 $Y=84790
X11654 3 digital_ldo_top_VIA18 $T=237590 84955 0 0 $X=237340 $Y=84790
X11655 3 digital_ldo_top_VIA18 $T=240350 84955 0 0 $X=240100 $Y=84790
X11656 3 digital_ldo_top_VIA18 $T=245870 84955 0 0 $X=245620 $Y=84790
X11657 3 digital_ldo_top_VIA18 $T=248630 84955 0 0 $X=248380 $Y=84790
X11658 3 digital_ldo_top_VIA18 $T=251390 84955 0 0 $X=251140 $Y=84790
X11659 3 digital_ldo_top_VIA18 $T=256910 84955 0 0 $X=256660 $Y=84790
X11660 3 digital_ldo_top_VIA18 $T=259670 84955 0 0 $X=259420 $Y=84790
X11661 3 digital_ldo_top_VIA18 $T=262430 84955 0 0 $X=262180 $Y=84790
X11662 3 digital_ldo_top_VIA18 $T=267950 84955 0 0 $X=267700 $Y=84790
X11663 3 digital_ldo_top_VIA18 $T=270710 84955 0 0 $X=270460 $Y=84790
X11664 3 digital_ldo_top_VIA18 $T=273470 84955 0 0 $X=273220 $Y=84790
X11665 3 digital_ldo_top_VIA18 $T=278990 84955 0 0 $X=278740 $Y=84790
X11666 3 digital_ldo_top_VIA18 $T=281750 84955 0 0 $X=281500 $Y=84790
X11667 3 digital_ldo_top_VIA18 $T=284510 84955 0 0 $X=284260 $Y=84790
X11668 3 digital_ldo_top_VIA18 $T=290030 84955 0 0 $X=289780 $Y=84790
X11669 3 digital_ldo_top_VIA18 $T=292790 84955 0 0 $X=292540 $Y=84790
X11670 2 MASCO__Y1 $T=305990 24300 0 0 $X=305990 $Y=24300
X11671 2 MASCO__Y1 $T=311510 44700 0 0 $X=311510 $Y=44700
X11672 2 MASCO__Y1 $T=311510 65100 0 0 $X=311510 $Y=65100
X11673 3 MASCO__Y1 $T=342790 17500 0 0 $X=342790 $Y=17500
X11674 3 MASCO__Y1 $T=342790 37900 0 0 $X=342790 $Y=37900
X11675 3 MASCO__Y1 $T=342790 58300 0 0 $X=342790 $Y=58300
X11676 3 MASCO__Y1 $T=342790 78700 0 0 $X=342790 $Y=78700
X11677 3 MASCO__Y1 $T=342790 99100 0 0 $X=342790 $Y=99100
X11678 3 MASCO__Y1 $T=342790 119500 0 0 $X=342790 $Y=119500
X11679 2 MASCO__Y1 $T=344630 24300 0 0 $X=344630 $Y=24300
X11680 2 MASCO__Y1 $T=344630 85500 0 0 $X=344630 $Y=85500
X11681 2 MASCO__Y1 $T=344630 105900 0 0 $X=344630 $Y=105900
X11682 2 MASCO__Y1 $T=344630 126300 0 0 $X=344630 $Y=126300
X11683 3 MASCO__Y2 $T=11590 17500 0 0 $X=11590 $Y=17500
X11684 3 MASCO__Y2 $T=11590 37900 0 0 $X=11590 $Y=37900
X11685 3 MASCO__Y2 $T=11590 58300 0 0 $X=11590 $Y=58300
X11686 3 MASCO__Y2 $T=11590 78700 0 0 $X=11590 $Y=78700
X11687 3 MASCO__Y2 $T=11590 99100 0 0 $X=11590 $Y=99100
X11688 3 MASCO__Y2 $T=11590 119500 0 0 $X=11590 $Y=119500
X11689 2 MASCO__Y2 $T=13430 24300 0 0 $X=13430 $Y=24300
X11690 2 MASCO__Y2 $T=13430 85500 0 0 $X=13430 $Y=85500
X11691 2 MASCO__Y2 $T=13430 105900 0 0 $X=13430 $Y=105900
X11692 2 MASCO__Y2 $T=13430 126300 0 0 $X=13430 $Y=126300
X11693 3 MASCO__Y2 $T=77830 17500 0 0 $X=77830 $Y=17500
X11694 3 MASCO__Y2 $T=77830 37900 0 0 $X=77830 $Y=37900
X11695 3 MASCO__Y2 $T=77830 58300 0 0 $X=77830 $Y=58300
X11696 3 MASCO__Y2 $T=77830 78700 0 0 $X=77830 $Y=78700
X11697 3 MASCO__Y2 $T=77830 99100 0 0 $X=77830 $Y=99100
X11698 3 MASCO__Y2 $T=77830 119500 0 0 $X=77830 $Y=119500
X11699 2 MASCO__Y2 $T=79670 85500 0 0 $X=79670 $Y=85500
X11700 2 MASCO__Y2 $T=79670 105900 0 0 $X=79670 $Y=105900
X11701 2 MASCO__Y2 $T=79670 126300 0 0 $X=79670 $Y=126300
X11702 3 MASCO__Y2 $T=144070 17500 0 0 $X=144070 $Y=17500
X11703 3 MASCO__Y2 $T=144070 37900 0 0 $X=144070 $Y=37900
X11704 3 MASCO__Y2 $T=144070 58300 0 0 $X=144070 $Y=58300
X11705 3 MASCO__Y2 $T=144070 78700 0 0 $X=144070 $Y=78700
X11706 3 MASCO__Y2 $T=144070 99100 0 0 $X=144070 $Y=99100
X11707 3 MASCO__Y2 $T=144070 119500 0 0 $X=144070 $Y=119500
X11708 2 MASCO__Y2 $T=145910 85500 0 0 $X=145910 $Y=85500
X11709 2 MASCO__Y2 $T=145910 105900 0 0 $X=145910 $Y=105900
X11710 2 MASCO__Y2 $T=145910 126300 0 0 $X=145910 $Y=126300
X11711 3 MASCO__Y2 $T=210310 17500 0 0 $X=210310 $Y=17500
X11712 3 MASCO__Y2 $T=210310 37900 0 0 $X=210310 $Y=37900
X11713 3 MASCO__Y2 $T=210310 58300 0 0 $X=210310 $Y=58300
X11714 3 MASCO__Y2 $T=210310 78700 0 0 $X=210310 $Y=78700
X11715 3 MASCO__Y2 $T=210310 99100 0 0 $X=210310 $Y=99100
X11716 3 MASCO__Y2 $T=210310 119500 0 0 $X=210310 $Y=119500
X11717 2 MASCO__Y2 $T=212150 85500 0 0 $X=212150 $Y=85500
X11718 2 MASCO__Y2 $T=212150 105900 0 0 $X=212150 $Y=105900
X11719 2 MASCO__Y2 $T=212150 126300 0 0 $X=212150 $Y=126300
X11720 3 MASCO__Y2 $T=276550 17500 0 0 $X=276550 $Y=17500
X11721 3 MASCO__Y2 $T=276550 37900 0 0 $X=276550 $Y=37900
X11722 3 MASCO__Y2 $T=276550 58300 0 0 $X=276550 $Y=58300
X11723 3 MASCO__Y2 $T=276550 78700 0 0 $X=276550 $Y=78700
X11724 3 MASCO__Y2 $T=276550 99100 0 0 $X=276550 $Y=99100
X11725 3 MASCO__Y2 $T=276550 119500 0 0 $X=276550 $Y=119500
X11726 2 MASCO__Y2 $T=278390 85500 0 0 $X=278390 $Y=85500
X11727 2 MASCO__Y2 $T=278390 105900 0 0 $X=278390 $Y=105900
X11728 2 MASCO__Y2 $T=278390 126300 0 0 $X=278390 $Y=126300
X11729 2 3 MASCO__B31 $T=13030 9760 0 0 $X=13030 $Y=9760
X11730 2 3 MASCO__B31 $T=13030 15200 0 0 $X=13030 $Y=15200
X11731 2 3 MASCO__B31 $T=13030 20640 0 0 $X=13030 $Y=20640
X11732 2 3 MASCO__B31 $T=13030 26080 0 0 $X=13030 $Y=26080
X11733 2 3 MASCO__B31 $T=13030 31520 0 0 $X=13030 $Y=31520
X11734 2 3 MASCO__B31 $T=13030 36960 0 0 $X=13030 $Y=36960
X11735 2 3 MASCO__B31 $T=13030 42400 0 0 $X=13030 $Y=42400
X11736 2 3 MASCO__B31 $T=13030 47840 0 0 $X=13030 $Y=47840
X11737 2 3 MASCO__B31 $T=13030 53280 0 0 $X=13030 $Y=53280
X11738 2 3 MASCO__B31 $T=13030 58720 0 0 $X=13030 $Y=58720
X11739 2 3 MASCO__B31 $T=13030 64160 0 0 $X=13030 $Y=64160
X11740 2 3 MASCO__B31 $T=13030 69600 0 0 $X=13030 $Y=69600
X11741 2 3 MASCO__B31 $T=13030 75040 0 0 $X=13030 $Y=75040
X11742 2 3 MASCO__B31 $T=13030 80480 0 0 $X=13030 $Y=80480
X11743 2 3 MASCO__B31 $T=13030 85920 0 0 $X=13030 $Y=85920
X11744 2 3 MASCO__B31 $T=13030 91360 0 0 $X=13030 $Y=91360
X11745 2 3 MASCO__B31 $T=13030 96800 0 0 $X=13030 $Y=96800
X11746 2 3 MASCO__B31 $T=13030 102240 0 0 $X=13030 $Y=102240
X11747 2 3 MASCO__B31 $T=13030 107680 0 0 $X=13030 $Y=107680
X11748 2 3 MASCO__B31 $T=13030 113120 0 0 $X=13030 $Y=113120
X11749 2 3 MASCO__B31 $T=13030 118560 0 0 $X=13030 $Y=118560
X11750 2 3 MASCO__B31 $T=13030 124000 0 0 $X=13030 $Y=124000
X11751 2 3 MASCO__B31 $T=61790 53280 0 0 $X=61790 $Y=53280
X11752 2 3 MASCO__B31 $T=99970 26080 0 0 $X=99970 $Y=26080
X11753 2 3 MASCO__B31 $T=99970 31520 0 0 $X=99970 $Y=31520
X11754 2 3 MASCO__B31 $T=99970 36960 0 0 $X=99970 $Y=36960
X11755 2 3 MASCO__B31 $T=101350 124000 0 0 $X=101350 $Y=124000
X11756 2 3 MASCO__B31 $T=130790 124000 0 0 $X=130790 $Y=124000
X11757 2 3 MASCO__B31 $T=160230 124000 0 0 $X=160230 $Y=124000
X11758 2 3 MASCO__B31 $T=189670 9760 0 0 $X=189670 $Y=9760
X11759 2 3 MASCO__B31 $T=189670 124000 0 0 $X=189670 $Y=124000
X11760 2 3 MASCO__B31 $T=219110 124000 0 0 $X=219110 $Y=124000
X11761 2 3 MASCO__B31 $T=233830 9760 0 0 $X=233830 $Y=9760
X11762 2 3 MASCO__B31 $T=248550 124000 0 0 $X=248550 $Y=124000
X11763 2 3 MASCO__B31 $T=277990 124000 0 0 $X=277990 $Y=124000
X11764 2 3 MASCO__B31 $T=307430 124000 0 0 $X=307430 $Y=124000
X11765 2 3 MASCO__B31 $T=320310 20640 0 0 $X=320310 $Y=20640
X11766 2 3 MASCO__B31 $T=320310 26080 0 0 $X=320310 $Y=26080
X11767 2 3 MASCO__B31 $T=320310 31520 0 0 $X=320310 $Y=31520
X11768 2 3 MASCO__B31 $T=320310 36960 0 0 $X=320310 $Y=36960
X11769 2 3 MASCO__B31 $T=320310 42400 0 0 $X=320310 $Y=42400
X11770 2 3 MASCO__B31 $T=366310 47840 0 0 $X=366310 $Y=47840
X11771 2 3 MASCO__B31 $T=366310 53280 0 0 $X=366310 $Y=53280
X11772 2 3 MASCO__B31 $T=366310 58720 0 0 $X=366310 $Y=58720
X11773 2 3 MASCO__B31 $T=366310 64160 0 0 $X=366310 $Y=64160
X11774 2 3 MASCO__B31 $T=366310 69600 0 0 $X=366310 $Y=69600
X11775 2 3 MASCO__B31 $T=366310 75040 0 0 $X=366310 $Y=75040
X11776 2 3 MASCO__B31 $T=366310 80480 0 0 $X=366310 $Y=80480
X11777 2 3 MASCO__B31 $T=366310 85920 0 0 $X=366310 $Y=85920
X11778 2 3 MASCO__B31 $T=366310 91360 0 0 $X=366310 $Y=91360
X11779 2 3 MASCO__B31 $T=366310 96800 0 0 $X=366310 $Y=96800
X11780 2 3 MASCO__B31 $T=366310 102240 0 0 $X=366310 $Y=102240
X11781 2 3 MASCO__B31 $T=366310 107680 0 0 $X=366310 $Y=107680
X11782 2 3 MASCO__B31 $T=366310 113120 0 0 $X=366310 $Y=113120
X11783 2 3 MASCO__B31 $T=366310 118560 0 0 $X=366310 $Y=118560
X11784 2 3 MASCO__B31 $T=366310 124000 0 0 $X=366310 $Y=124000
X11785 2 3 MASCO__B31 $T=377350 47840 0 0 $X=377350 $Y=47840
X11786 2 3 MASCO__B31 $T=377350 53280 0 0 $X=377350 $Y=53280
X11787 2 3 MASCO__B31 $T=377350 58720 0 0 $X=377350 $Y=58720
X11788 2 3 MASCO__B31 $T=377350 64160 0 0 $X=377350 $Y=64160
X11789 2 3 MASCO__B31 $T=377350 69600 0 0 $X=377350 $Y=69600
X11790 2 3 MASCO__B31 $T=377350 75040 0 0 $X=377350 $Y=75040
X11791 2 3 MASCO__B31 $T=377350 80480 0 0 $X=377350 $Y=80480
X11792 2 3 MASCO__B31 $T=377350 85920 0 0 $X=377350 $Y=85920
X11793 2 3 MASCO__B31 $T=377350 91360 0 0 $X=377350 $Y=91360
X11794 2 3 MASCO__B31 $T=377350 96800 0 0 $X=377350 $Y=96800
X11795 2 3 MASCO__B31 $T=377350 102240 0 0 $X=377350 $Y=102240
X11796 2 3 MASCO__B31 $T=377350 107680 0 0 $X=377350 $Y=107680
X11797 2 3 MASCO__B31 $T=377350 113120 0 0 $X=377350 $Y=113120
X11798 2 3 MASCO__B31 $T=377350 118560 0 0 $X=377350 $Y=118560
X11799 2 3 MASCO__B31 $T=377350 124000 0 0 $X=377350 $Y=124000
X11800 3 2 MASCO__B32 $T=90770 26080 0 0 $X=90770 $Y=26080
X11801 3 2 MASCO__B32 $T=90770 31520 0 0 $X=90770 $Y=31520
X11802 3 2 MASCO__B32 $T=90770 36960 0 0 $X=90770 $Y=36960
X11803 3 2 MASCO__B32 $T=368150 47840 0 0 $X=368150 $Y=47840
X11804 3 2 MASCO__B32 $T=368150 53280 0 0 $X=368150 $Y=53280
X11805 3 2 MASCO__B32 $T=368150 58720 0 0 $X=368150 $Y=58720
X11806 3 2 MASCO__B32 $T=368150 64160 0 0 $X=368150 $Y=64160
X11807 3 2 MASCO__B32 $T=368150 69600 0 0 $X=368150 $Y=69600
X11808 3 2 MASCO__B32 $T=368150 75040 0 0 $X=368150 $Y=75040
X11809 3 2 MASCO__B32 $T=368150 80480 0 0 $X=368150 $Y=80480
X11810 3 2 MASCO__B32 $T=368150 85920 0 0 $X=368150 $Y=85920
X11811 3 2 MASCO__B32 $T=368150 91360 0 0 $X=368150 $Y=91360
X11812 3 2 MASCO__B32 $T=368150 96800 0 0 $X=368150 $Y=96800
X11813 3 2 MASCO__B32 $T=368150 102240 0 0 $X=368150 $Y=102240
X11814 3 2 MASCO__B32 $T=368150 107680 0 0 $X=368150 $Y=107680
X11815 3 2 MASCO__B32 $T=368150 113120 0 0 $X=368150 $Y=113120
X11816 3 2 MASCO__B32 $T=368150 118560 0 0 $X=368150 $Y=118560
X11817 3 2 MASCO__B32 $T=368150 124000 0 0 $X=368150 $Y=124000
X11818 3 2 MASCO__B33 $T=29130 34240 0 0 $X=29130 $Y=34240
X11819 3 2 MASCO__B33 $T=29130 39680 0 0 $X=29130 $Y=39680
X11820 3 2 MASCO__B33 $T=29130 45120 0 0 $X=29130 $Y=45120
X11821 3 2 MASCO__B33 $T=29130 50560 0 0 $X=29130 $Y=50560
X11822 3 2 MASCO__B33 $T=29130 56000 0 0 $X=29130 $Y=56000
X11823 3 2 MASCO__B33 $T=29130 61440 0 0 $X=29130 $Y=61440
X11824 3 2 MASCO__B33 $T=29130 66880 0 0 $X=29130 $Y=66880
X11825 3 2 MASCO__B33 $T=29130 72320 0 0 $X=29130 $Y=72320
X11826 3 2 MASCO__B33 $T=29130 77760 0 0 $X=29130 $Y=77760
X11827 3 2 MASCO__B33 $T=29130 83200 0 0 $X=29130 $Y=83200
X11828 3 2 MASCO__B33 $T=29130 88640 0 0 $X=29130 $Y=88640
X11829 3 2 MASCO__B33 $T=29130 94080 0 0 $X=29130 $Y=94080
X11830 3 2 MASCO__B33 $T=29130 99520 0 0 $X=29130 $Y=99520
X11831 3 2 MASCO__B33 $T=29130 104960 0 0 $X=29130 $Y=104960
X11832 3 2 MASCO__B33 $T=29130 110400 0 0 $X=29130 $Y=110400
X11833 3 2 MASCO__B33 $T=29130 115840 0 0 $X=29130 $Y=115840
X11834 3 2 MASCO__B33 $T=29130 121280 0 0 $X=29130 $Y=121280
X11835 3 2 MASCO__B33 $T=88010 45120 0 0 $X=88010 $Y=45120
X11836 3 2 MASCO__B33 $T=88010 50560 0 0 $X=88010 $Y=50560
X11837 3 2 MASCO__B33 $T=88010 56000 0 0 $X=88010 $Y=56000
X11838 3 2 MASCO__B33 $T=323530 50560 0 0 $X=323530 $Y=50560
X11839 3 2 MASCO__B33 $T=323530 56000 0 0 $X=323530 $Y=56000
X11840 3 2 MASCO__B33 $T=323530 61440 0 0 $X=323530 $Y=61440
X11841 3 2 MASCO__B33 $T=323530 66880 0 0 $X=323530 $Y=66880
X11842 3 2 MASCO__B33 $T=323530 72320 0 0 $X=323530 $Y=72320
X11843 3 2 MASCO__B33 $T=323530 77760 0 0 $X=323530 $Y=77760
X11844 3 2 MASCO__B33 $T=323530 83200 0 0 $X=323530 $Y=83200
X11845 3 2 MASCO__B33 $T=323530 88640 0 0 $X=323530 $Y=88640
X11846 3 2 MASCO__B33 $T=323530 94080 0 0 $X=323530 $Y=94080
X11847 3 2 MASCO__B33 $T=323530 99520 0 0 $X=323530 $Y=99520
X11848 3 2 MASCO__B33 $T=323530 104960 0 0 $X=323530 $Y=104960
X11849 3 2 MASCO__B33 $T=323530 110400 0 0 $X=323530 $Y=110400
X11850 3 2 MASCO__B33 $T=323530 115840 0 0 $X=323530 $Y=115840
X11851 3 2 MASCO__B33 $T=323530 121280 0 0 $X=323530 $Y=121280
X11852 3 2 MASCO__B33 $T=367690 12480 0 0 $X=367690 $Y=12480
X11853 3 2 MASCO__B33 $T=367690 17920 0 0 $X=367690 $Y=17920
X11854 3 2 MASCO__B33 $T=367690 23360 0 0 $X=367690 $Y=23360
X11855 3 2 MASCO__B33 $T=367690 28800 0 0 $X=367690 $Y=28800
X11856 3 2 MASCO__B33 $T=367690 34240 0 0 $X=367690 $Y=34240
X11857 3 2 MASCO__B33 $T=367690 39680 0 0 $X=367690 $Y=39680
X11858 3 2 MASCO__B35 $T=93990 64160 0 0 $X=93990 $Y=64160
X11859 3 2 MASCO__B35 $T=93990 69600 0 0 $X=93990 $Y=69600
X11860 3 2 MASCO__B35 $T=93990 75040 0 0 $X=93990 $Y=75040
X11861 3 2 MASCO__B35 $T=93990 80480 0 0 $X=93990 $Y=80480
X11862 3 2 MASCO__B35 $T=93990 85920 0 0 $X=93990 $Y=85920
X11863 3 2 MASCO__B35 $T=93990 124000 0 0 $X=93990 $Y=124000
X11864 3 2 MASCO__B35 $T=123430 124000 0 0 $X=123430 $Y=124000
X11865 3 2 MASCO__B35 $T=152870 124000 0 0 $X=152870 $Y=124000
X11866 3 2 MASCO__B35 $T=182310 9760 0 0 $X=182310 $Y=9760
X11867 3 2 MASCO__B35 $T=182310 124000 0 0 $X=182310 $Y=124000
X11868 3 2 MASCO__B35 $T=211750 124000 0 0 $X=211750 $Y=124000
X11869 3 2 MASCO__B35 $T=241190 124000 0 0 $X=241190 $Y=124000
X11870 3 2 MASCO__B35 $T=270630 124000 0 0 $X=270630 $Y=124000
X11871 3 2 MASCO__B35 $T=300070 124000 0 0 $X=300070 $Y=124000
X11872 3 2 MASCO__B35 $T=358950 124000 0 0 $X=358950 $Y=124000
X11873 3 2 MASCO__B37 $T=88010 64160 0 0 $X=88010 $Y=64160
X11874 3 2 MASCO__B37 $T=88010 69600 0 0 $X=88010 $Y=69600
X11875 3 2 MASCO__B37 $T=88010 75040 0 0 $X=88010 $Y=75040
X11876 3 2 MASCO__B37 $T=88010 80480 0 0 $X=88010 $Y=80480
X11877 3 2 MASCO__B37 $T=88010 85920 0 0 $X=88010 $Y=85920
X11878 3 2 MASCO__B37 $T=88010 91360 0 0 $X=88010 $Y=91360
X11879 3 2 MASCO__B37 $T=88010 96800 0 0 $X=88010 $Y=96800
X11880 3 2 MASCO__B37 $T=88010 102240 0 0 $X=88010 $Y=102240
X11881 3 2 MASCO__B37 $T=88010 107680 0 0 $X=88010 $Y=107680
X11882 3 2 MASCO__B37 $T=88010 113120 0 0 $X=88010 $Y=113120
X11883 3 2 MASCO__B37 $T=88010 118560 0 0 $X=88010 $Y=118560
X11884 3 2 MASCO__B37 $T=88010 124000 0 0 $X=88010 $Y=124000
X11885 3 2 MASCO__B37 $T=102730 9760 0 0 $X=102730 $Y=9760
X11886 3 2 MASCO__B37 $T=117450 124000 0 0 $X=117450 $Y=124000
X11887 3 2 MASCO__B37 $T=146890 91360 0 0 $X=146890 $Y=91360
X11888 3 2 MASCO__B37 $T=146890 96800 0 0 $X=146890 $Y=96800
X11889 3 2 MASCO__B37 $T=146890 102240 0 0 $X=146890 $Y=102240
X11890 3 2 MASCO__B37 $T=146890 107680 0 0 $X=146890 $Y=107680
X11891 3 2 MASCO__B37 $T=146890 113120 0 0 $X=146890 $Y=113120
X11892 3 2 MASCO__B37 $T=146890 118560 0 0 $X=146890 $Y=118560
X11893 3 2 MASCO__B37 $T=146890 124000 0 0 $X=146890 $Y=124000
X11894 3 2 MASCO__B37 $T=161610 9760 0 0 $X=161610 $Y=9760
X11895 3 2 MASCO__B37 $T=176330 9760 0 0 $X=176330 $Y=9760
X11896 3 2 MASCO__B37 $T=176330 124000 0 0 $X=176330 $Y=124000
X11897 3 2 MASCO__B37 $T=205770 91360 0 0 $X=205770 $Y=91360
X11898 3 2 MASCO__B37 $T=205770 96800 0 0 $X=205770 $Y=96800
X11899 3 2 MASCO__B37 $T=205770 102240 0 0 $X=205770 $Y=102240
X11900 3 2 MASCO__B37 $T=205770 107680 0 0 $X=205770 $Y=107680
X11901 3 2 MASCO__B37 $T=205770 113120 0 0 $X=205770 $Y=113120
X11902 3 2 MASCO__B37 $T=205770 118560 0 0 $X=205770 $Y=118560
X11903 3 2 MASCO__B37 $T=205770 124000 0 0 $X=205770 $Y=124000
X11904 3 2 MASCO__B37 $T=235210 124000 0 0 $X=235210 $Y=124000
X11905 3 2 MASCO__B37 $T=249930 9760 0 0 $X=249930 $Y=9760
X11906 3 2 MASCO__B37 $T=264650 91360 0 0 $X=264650 $Y=91360
X11907 3 2 MASCO__B37 $T=264650 96800 0 0 $X=264650 $Y=96800
X11908 3 2 MASCO__B37 $T=264650 102240 0 0 $X=264650 $Y=102240
X11909 3 2 MASCO__B37 $T=264650 107680 0 0 $X=264650 $Y=107680
X11910 3 2 MASCO__B37 $T=264650 113120 0 0 $X=264650 $Y=113120
X11911 3 2 MASCO__B37 $T=264650 118560 0 0 $X=264650 $Y=118560
X11912 3 2 MASCO__B37 $T=264650 124000 0 0 $X=264650 $Y=124000
X11913 3 2 MASCO__B37 $T=294090 124000 0 0 $X=294090 $Y=124000
X11914 3 2 MASCO__B37 $T=308810 9760 0 0 $X=308810 $Y=9760
X11915 3 2 MASCO__B37 $T=352970 124000 0 0 $X=352970 $Y=124000
X11916 3 2 MASCO__B39 $T=35110 34240 0 0 $X=35110 $Y=34240
X11917 3 2 MASCO__B39 $T=35110 39680 0 0 $X=35110 $Y=39680
X11918 3 2 MASCO__B39 $T=35110 45120 0 0 $X=35110 $Y=45120
X11919 3 2 MASCO__B39 $T=35110 50560 0 0 $X=35110 $Y=50560
X11920 3 2 MASCO__B39 $T=35110 56000 0 0 $X=35110 $Y=56000
X11921 3 2 MASCO__B39 $T=61790 34240 0 0 $X=61790 $Y=34240
X11922 3 2 MASCO__B39 $T=61790 39680 0 0 $X=61790 $Y=39680
X11923 3 2 MASCO__B39 $T=61790 45120 0 0 $X=61790 $Y=45120
X11924 3 2 MASCO__B39 $T=71910 34240 0 0 $X=71910 $Y=34240
X11925 3 2 MASCO__B39 $T=71910 39680 0 0 $X=71910 $Y=39680
X11926 3 2 MASCO__B39 $T=71910 45120 0 0 $X=71910 $Y=45120
X11927 3 2 MASCO__B39 $T=71910 50560 0 0 $X=71910 $Y=50560
X11928 3 2 MASCO__B39 $T=71910 56000 0 0 $X=71910 $Y=56000
X11929 3 2 MASCO__B39 $T=99970 17920 0 0 $X=99970 $Y=17920
X11930 3 2 MASCO__B39 $T=145510 12480 0 0 $X=145510 $Y=12480
X11931 3 2 MASCO__B39 $T=336870 50560 0 0 $X=336870 $Y=50560
X11932 3 2 MASCO__B39 $T=336870 56000 0 0 $X=336870 $Y=56000
X11933 3 2 MASCO__B39 $T=336870 61440 0 0 $X=336870 $Y=61440
X11934 3 2 MASCO__B39 $T=336870 66880 0 0 $X=336870 $Y=66880
X11935 3 2 MASCO__B39 $T=336870 72320 0 0 $X=336870 $Y=72320
X11936 3 2 MASCO__B39 $T=336870 77760 0 0 $X=336870 $Y=77760
X11937 3 2 MASCO__B39 $T=336870 83200 0 0 $X=336870 $Y=83200
X11938 3 2 MASCO__B39 $T=336870 88640 0 0 $X=336870 $Y=88640
X11939 3 2 MASCO__B39 $T=336870 94080 0 0 $X=336870 $Y=94080
X11940 3 2 MASCO__B39 $T=336870 99520 0 0 $X=336870 $Y=99520
X11941 3 2 MASCO__B39 $T=336870 104960 0 0 $X=336870 $Y=104960
X11942 3 2 MASCO__B39 $T=336870 110400 0 0 $X=336870 $Y=110400
X11943 3 2 MASCO__B39 $T=336870 115840 0 0 $X=336870 $Y=115840
X11944 3 2 MASCO__B39 $T=336870 121280 0 0 $X=336870 $Y=121280
X11945 3 2 MASCO__B40 $T=93990 45120 0 0 $X=93990 $Y=45120
X11946 3 2 MASCO__B40 $T=93990 50560 0 0 $X=93990 $Y=50560
X11947 3 2 MASCO__B40 $T=93990 56000 0 0 $X=93990 $Y=56000
X11948 3 2 MASCO__B40 $T=329510 50560 0 0 $X=329510 $Y=50560
X11949 3 2 MASCO__B40 $T=329510 56000 0 0 $X=329510 $Y=56000
X11950 3 2 MASCO__B40 $T=329510 61440 0 0 $X=329510 $Y=61440
X11951 3 2 MASCO__B40 $T=329510 66880 0 0 $X=329510 $Y=66880
X11952 3 2 MASCO__B40 $T=329510 72320 0 0 $X=329510 $Y=72320
X11953 3 2 MASCO__B40 $T=329510 77760 0 0 $X=329510 $Y=77760
X11954 3 2 MASCO__B40 $T=329510 83200 0 0 $X=329510 $Y=83200
X11955 3 2 MASCO__B40 $T=329510 88640 0 0 $X=329510 $Y=88640
X11956 3 2 MASCO__B40 $T=329510 94080 0 0 $X=329510 $Y=94080
X11957 3 2 MASCO__B40 $T=329510 99520 0 0 $X=329510 $Y=99520
X11958 3 2 MASCO__B40 $T=329510 104960 0 0 $X=329510 $Y=104960
X11959 3 2 MASCO__B40 $T=329510 110400 0 0 $X=329510 $Y=110400
X11960 3 2 MASCO__B40 $T=329510 115840 0 0 $X=329510 $Y=115840
X11961 3 2 MASCO__B40 $T=329510 121280 0 0 $X=329510 $Y=121280
X11962 3 2 MASCO__B63 $T=14870 34240 0 0 $X=14870 $Y=34240
X11963 3 2 MASCO__B63 $T=14870 45120 0 0 $X=14870 $Y=45120
X11964 3 2 MASCO__B63 $T=14870 56000 0 0 $X=14870 $Y=56000
X11965 3 2 MASCO__B63 $T=14870 66880 0 0 $X=14870 $Y=66880
X11966 3 2 MASCO__B63 $T=14870 77760 0 0 $X=14870 $Y=77760
X11967 3 2 MASCO__B63 $T=14870 88640 0 0 $X=14870 $Y=88640
X11968 3 2 MASCO__B63 $T=14870 99520 0 0 $X=14870 $Y=99520
X11969 3 2 MASCO__B63 $T=14870 110400 0 0 $X=14870 $Y=110400
X11970 3 2 MASCO__B63 $T=73750 45120 0 0 $X=73750 $Y=45120
X11971 3 2 MASCO__B63 $T=338710 50560 0 0 $X=338710 $Y=50560
X11972 3 2 MASCO__B63 $T=338710 61440 0 0 $X=338710 $Y=61440
X11973 3 2 MASCO__B63 $T=338710 72320 0 0 $X=338710 $Y=72320
X11974 3 2 MASCO__B63 $T=338710 83200 0 0 $X=338710 $Y=83200
X11975 3 2 MASCO__B63 $T=338710 94080 0 0 $X=338710 $Y=94080
X11976 3 2 MASCO__B63 $T=338710 104960 0 0 $X=338710 $Y=104960
X11977 3 2 MASCO__B63 $T=338710 115840 0 0 $X=338710 $Y=115840
X11978 3 2 MASCO__B63 $T=353430 12480 0 0 $X=353430 $Y=12480
X11979 3 2 MASCO__B63 $T=353430 23360 0 0 $X=353430 $Y=23360
X11980 3 2 MASCO__B63 $T=353430 34240 0 0 $X=353430 $Y=34240
X11981 3 2 MASCO__B64 $T=58570 64160 0 0 $X=58570 $Y=64160
X11982 3 2 MASCO__B64 $T=58570 75040 0 0 $X=58570 $Y=75040
X11983 3 2 MASCO__B64 $T=58570 85920 0 0 $X=58570 $Y=85920
X11984 3 2 MASCO__B64 $T=58570 96800 0 0 $X=58570 $Y=96800
X11985 3 2 MASCO__B64 $T=58570 107680 0 0 $X=58570 $Y=107680
X11986 3 2 MASCO__B64 $T=58570 118560 0 0 $X=58570 $Y=118560
X11987 3 2 MASCO__B64 $T=117450 91360 0 0 $X=117450 $Y=91360
X11988 3 2 MASCO__B64 $T=117450 102240 0 0 $X=117450 $Y=102240
X11989 3 2 MASCO__B64 $T=117450 113120 0 0 $X=117450 $Y=113120
X11990 3 2 MASCO__B64 $T=176330 91360 0 0 $X=176330 $Y=91360
X11991 3 2 MASCO__B64 $T=176330 102240 0 0 $X=176330 $Y=102240
X11992 3 2 MASCO__B64 $T=176330 113120 0 0 $X=176330 $Y=113120
X11993 3 2 MASCO__B64 $T=235210 91360 0 0 $X=235210 $Y=91360
X11994 3 2 MASCO__B64 $T=235210 102240 0 0 $X=235210 $Y=102240
X11995 3 2 MASCO__B64 $T=235210 113120 0 0 $X=235210 $Y=113120
X11996 3 2 MASCO__B64 $T=294090 91360 0 0 $X=294090 $Y=91360
X11997 3 2 MASCO__B64 $T=294090 102240 0 0 $X=294090 $Y=102240
X11998 3 2 MASCO__B64 $T=294090 113120 0 0 $X=294090 $Y=113120
X11999 3 2 MASCO__B64 $T=352970 47840 0 0 $X=352970 $Y=47840
X12000 3 2 MASCO__B64 $T=352970 58720 0 0 $X=352970 $Y=58720
X12001 3 2 MASCO__B64 $T=352970 69600 0 0 $X=352970 $Y=69600
X12002 3 2 MASCO__B64 $T=352970 80480 0 0 $X=352970 $Y=80480
X12003 3 2 MASCO__B64 $T=352970 91360 0 0 $X=352970 $Y=91360
X12004 3 2 MASCO__B64 $T=352970 102240 0 0 $X=352970 $Y=102240
X12005 3 2 MASCO__B64 $T=352970 113120 0 0 $X=352970 $Y=113120
X12006 3 2 MASCO__B65 $T=71910 64160 0 0 $X=71910 $Y=64160
X12007 3 2 MASCO__B65 $T=71910 75040 0 0 $X=71910 $Y=75040
X12008 3 2 MASCO__B65 $T=71910 85920 0 0 $X=71910 $Y=85920
X12009 3 2 MASCO__B65 $T=71910 96800 0 0 $X=71910 $Y=96800
X12010 3 2 MASCO__B65 $T=71910 107680 0 0 $X=71910 $Y=107680
X12011 3 2 MASCO__B65 $T=71910 118560 0 0 $X=71910 $Y=118560
X12012 3 2 MASCO__B65 $T=130790 91360 0 0 $X=130790 $Y=91360
X12013 3 2 MASCO__B65 $T=130790 102240 0 0 $X=130790 $Y=102240
X12014 3 2 MASCO__B65 $T=130790 113120 0 0 $X=130790 $Y=113120
X12015 3 2 MASCO__B65 $T=189670 91360 0 0 $X=189670 $Y=91360
X12016 3 2 MASCO__B65 $T=189670 102240 0 0 $X=189670 $Y=102240
X12017 3 2 MASCO__B65 $T=189670 113120 0 0 $X=189670 $Y=113120
X12018 3 2 MASCO__B65 $T=248550 91360 0 0 $X=248550 $Y=91360
X12019 3 2 MASCO__B65 $T=248550 102240 0 0 $X=248550 $Y=102240
X12020 3 2 MASCO__B65 $T=248550 113120 0 0 $X=248550 $Y=113120
X12021 3 2 MASCO__B65 $T=307430 20640 0 0 $X=307430 $Y=20640
X12022 3 2 MASCO__B65 $T=307430 31520 0 0 $X=307430 $Y=31520
X12023 3 2 MASCO__B65 $T=307430 42400 0 0 $X=307430 $Y=42400
X12024 3 2 MASCO__B65 $T=307430 53280 0 0 $X=307430 $Y=53280
X12025 3 2 MASCO__B65 $T=307430 64160 0 0 $X=307430 $Y=64160
X12026 3 2 MASCO__B65 $T=307430 75040 0 0 $X=307430 $Y=75040
X12027 3 2 MASCO__B65 $T=307430 91360 0 0 $X=307430 $Y=91360
X12028 3 2 MASCO__B65 $T=307430 102240 0 0 $X=307430 $Y=102240
X12029 3 2 MASCO__B65 $T=307430 113120 0 0 $X=307430 $Y=113120
X12030 3 2 MASCO__B66 $T=44310 64160 0 0 $X=44310 $Y=64160
X12031 3 2 MASCO__B66 $T=44310 75040 0 0 $X=44310 $Y=75040
X12032 3 2 MASCO__B66 $T=44310 85920 0 0 $X=44310 $Y=85920
X12033 3 2 MASCO__B66 $T=44310 96800 0 0 $X=44310 $Y=96800
X12034 3 2 MASCO__B66 $T=44310 107680 0 0 $X=44310 $Y=107680
X12035 3 2 MASCO__B66 $T=44310 118560 0 0 $X=44310 $Y=118560
X12036 3 2 MASCO__B66 $T=103190 91360 0 0 $X=103190 $Y=91360
X12037 3 2 MASCO__B66 $T=103190 102240 0 0 $X=103190 $Y=102240
X12038 3 2 MASCO__B66 $T=103190 113120 0 0 $X=103190 $Y=113120
X12039 3 2 MASCO__B66 $T=162070 91360 0 0 $X=162070 $Y=91360
X12040 3 2 MASCO__B66 $T=162070 102240 0 0 $X=162070 $Y=102240
X12041 3 2 MASCO__B66 $T=162070 113120 0 0 $X=162070 $Y=113120
X12042 3 2 MASCO__B66 $T=220950 91360 0 0 $X=220950 $Y=91360
X12043 3 2 MASCO__B66 $T=220950 102240 0 0 $X=220950 $Y=102240
X12044 3 2 MASCO__B66 $T=220950 113120 0 0 $X=220950 $Y=113120
X12045 3 2 MASCO__B66 $T=279830 91360 0 0 $X=279830 $Y=91360
X12046 3 2 MASCO__B66 $T=279830 102240 0 0 $X=279830 $Y=102240
X12047 3 2 MASCO__B66 $T=279830 113120 0 0 $X=279830 $Y=113120
X12048 3 2 MASCO__B67 $T=35110 64160 0 0 $X=35110 $Y=64160
X12049 3 2 MASCO__B67 $T=35110 75040 0 0 $X=35110 $Y=75040
X12050 3 2 MASCO__B67 $T=35110 85920 0 0 $X=35110 $Y=85920
X12051 3 2 MASCO__B67 $T=35110 96800 0 0 $X=35110 $Y=96800
X12052 3 2 MASCO__B67 $T=35110 107680 0 0 $X=35110 $Y=107680
X12053 3 2 MASCO__B67 $T=35110 118560 0 0 $X=35110 $Y=118560
X12054 3 2 MASCO__B67 $T=93990 91360 0 0 $X=93990 $Y=91360
X12055 3 2 MASCO__B67 $T=93990 102240 0 0 $X=93990 $Y=102240
X12056 3 2 MASCO__B67 $T=93990 113120 0 0 $X=93990 $Y=113120
X12057 3 2 MASCO__B67 $T=152870 91360 0 0 $X=152870 $Y=91360
X12058 3 2 MASCO__B67 $T=152870 102240 0 0 $X=152870 $Y=102240
X12059 3 2 MASCO__B67 $T=152870 113120 0 0 $X=152870 $Y=113120
X12060 3 2 MASCO__B67 $T=211750 91360 0 0 $X=211750 $Y=91360
X12061 3 2 MASCO__B67 $T=211750 102240 0 0 $X=211750 $Y=102240
X12062 3 2 MASCO__B67 $T=211750 113120 0 0 $X=211750 $Y=113120
X12063 3 2 MASCO__B67 $T=270630 91360 0 0 $X=270630 $Y=91360
X12064 3 2 MASCO__B67 $T=270630 102240 0 0 $X=270630 $Y=102240
X12065 3 2 MASCO__B67 $T=270630 113120 0 0 $X=270630 $Y=113120
.ends digital_ldo_top
