VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DigitalLDOLogic
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN DigitalLDOLogic 0 0 ;
  SIZE 200.1 BY 70.04 ;
  SYMMETRY X Y ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 129.45 13.475 131.23 13.855 ;
        RECT 120.865 13.475 122.675 13.855 ;
      LAYER met1 ;
        RECT 130.25 13.64 130.57 13.9 ;
        RECT 129.805 13.655 130.57 13.885 ;
        RECT 121.985 13.7 130.57 13.84 ;
        RECT 121.985 13.655 122.735 13.885 ;
      LAYER met3 ;
        RECT 189.585 1.325 189.915 1.655 ;
        RECT 188.68 1.34 189.915 1.64 ;
        RECT 188.68 0.73 188.98 1.64 ;
        RECT 129.8 0.73 188.98 1.03 ;
        RECT 129.785 1.935 130.115 2.265 ;
        RECT 129.8 0.73 130.1 2.265 ;
      LAYER met2 ;
        RECT 189.61 1.305 189.89 1.675 ;
        RECT 189.68 0 189.82 1.675 ;
        RECT 130.28 13.61 130.54 13.93 ;
        RECT 130.34 2.03 130.48 13.93 ;
        RECT 129.81 2.03 130.48 2.17 ;
        RECT 129.81 1.915 130.09 2.285 ;
      LAYER via ;
        RECT 130.335 13.695 130.485 13.845 ;
      LAYER via2 ;
        RECT 129.85 2 130.05 2.2 ;
        RECT 189.65 1.39 189.85 1.59 ;
      LAYER mcon ;
        RECT 122.045 13.685 122.215 13.855 ;
        RECT 122.505 13.685 122.675 13.855 ;
        RECT 129.865 13.685 130.035 13.855 ;
        RECT 130.325 13.685 130.495 13.855 ;
    END
  END clk
  PIN comp_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 170.765 13.565 171.105 13.935 ;
        RECT 148.225 22.135 148.555 22.385 ;
        RECT 142.225 22.105 142.58 22.475 ;
      LAYER met1 ;
        RECT 171.65 13.64 171.97 13.9 ;
        RECT 166.13 13.7 171.97 13.84 ;
        RECT 170.745 13.655 171.035 13.885 ;
        RECT 166.13 13.64 166.45 13.9 ;
        RECT 166.13 22.48 166.45 22.74 ;
        RECT 165.3 22.54 166.45 22.68 ;
        RECT 165.3 22.2 165.44 22.68 ;
        RECT 155.18 22.2 165.44 22.34 ;
        RECT 148.28 22.54 155.32 22.68 ;
        RECT 155.18 22.2 155.32 22.68 ;
        RECT 148.205 22.155 148.495 22.385 ;
        RECT 148.28 22.155 148.42 22.68 ;
        RECT 147.36 22.2 148.495 22.34 ;
        RECT 144.6 22.37 147.5 22.51 ;
        RECT 147.36 22.2 147.5 22.51 ;
        RECT 143.68 22.54 144.74 22.68 ;
        RECT 144.6 22.37 144.74 22.68 ;
        RECT 143.68 22.2 143.82 22.68 ;
        RECT 142.225 22.2 143.82 22.34 ;
        RECT 142.225 22.155 142.515 22.385 ;
      LAYER met2 ;
        RECT 171.68 13.61 171.94 13.93 ;
        RECT 171.74 13.02 171.88 13.93 ;
        RECT 171.28 13.02 171.88 13.16 ;
        RECT 171.28 8.94 171.42 13.16 ;
        RECT 170.82 8.94 171.42 9.08 ;
        RECT 170.82 0 170.96 9.08 ;
        RECT 166.16 22.45 166.42 22.77 ;
        RECT 166.16 13.61 166.42 13.93 ;
        RECT 166.22 13.61 166.36 22.77 ;
      LAYER via ;
        RECT 166.215 22.535 166.365 22.685 ;
        RECT 166.215 13.695 166.365 13.845 ;
        RECT 171.735 13.695 171.885 13.845 ;
      LAYER mcon ;
        RECT 142.285 22.185 142.455 22.355 ;
        RECT 148.265 22.185 148.435 22.355 ;
        RECT 170.805 13.685 170.975 13.855 ;
    END
  END comp_in
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.855 20.995 22.025 23.205 ;
        RECT 19.335 22.555 22.025 22.725 ;
        RECT 21.77 21.845 22.025 22.725 ;
        RECT 19.335 21.845 22.025 22.015 ;
        RECT 21.015 22.555 21.185 23.205 ;
        RECT 21.015 20.995 21.185 22.015 ;
        RECT 20.175 22.555 20.345 23.205 ;
        RECT 20.175 20.995 20.345 22.015 ;
        RECT 19.335 22.555 19.505 23.205 ;
        RECT 19.335 20.995 19.505 22.015 ;
      LAYER met1 ;
        RECT 19.405 21.815 19.695 22.045 ;
        RECT 10.28 21.86 19.695 22 ;
        RECT 10.19 21.46 10.51 21.72 ;
        RECT 10.28 21.46 10.42 22 ;
      LAYER met2 ;
        RECT 10.22 21.43 10.48 21.75 ;
        RECT 10.28 0 10.42 21.75 ;
      LAYER via ;
        RECT 10.275 21.515 10.425 21.665 ;
      LAYER mcon ;
        RECT 19.465 21.845 19.635 22.015 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.615 18.275 24.785 20.485 ;
        RECT 22.095 19.465 24.785 19.635 ;
        RECT 24.53 18.755 24.785 19.635 ;
        RECT 22.095 18.755 24.785 18.925 ;
        RECT 23.775 19.465 23.945 20.485 ;
        RECT 23.775 18.275 23.945 18.925 ;
        RECT 22.935 19.465 23.105 20.485 ;
        RECT 22.935 18.275 23.105 18.925 ;
        RECT 22.095 19.465 22.265 20.485 ;
        RECT 22.095 18.275 22.265 18.925 ;
      LAYER met1 ;
        RECT 22.165 19.435 22.455 19.665 ;
        RECT 19.85 19.48 22.455 19.62 ;
        RECT 19.85 19.42 20.17 19.68 ;
      LAYER met2 ;
        RECT 19.88 19.39 20.14 19.71 ;
        RECT 19.94 0 20.08 19.71 ;
      LAYER via ;
        RECT 19.935 19.475 20.085 19.625 ;
      LAYER mcon ;
        RECT 22.225 19.465 22.395 19.635 ;
    END
  END out[16]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 33.395 22.555 33.565 23.205 ;
        RECT 30.875 21.845 33.565 22.015 ;
        RECT 33.395 20.995 33.565 22.015 ;
        RECT 30.875 22.555 33.565 22.725 ;
        RECT 32.555 22.555 32.725 23.205 ;
        RECT 32.555 20.995 32.725 22.015 ;
        RECT 31.715 22.555 31.885 23.205 ;
        RECT 31.715 20.995 31.885 22.015 ;
        RECT 30.875 21.845 31.13 22.725 ;
        RECT 30.875 20.995 31.045 23.205 ;
      LAYER met1 ;
        RECT 30.89 21.8 31.21 22.06 ;
      LAYER met2 ;
        RECT 30.92 21.77 31.18 22.09 ;
        RECT 30.52 21.86 31.18 22 ;
        RECT 30.52 20.84 30.89 20.98 ;
        RECT 30.75 14.72 30.89 20.98 ;
        RECT 30.52 14.72 30.89 14.86 ;
        RECT 30.52 20.84 30.66 22 ;
        RECT 30.52 8.94 30.66 14.86 ;
        RECT 29.6 8.94 30.66 9.08 ;
        RECT 29.6 0 29.74 9.08 ;
      LAYER via ;
        RECT 30.975 21.855 31.125 22.005 ;
      LAYER mcon ;
        RECT 30.965 21.845 31.135 22.015 ;
    END
  END out[17]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 41.675 22.555 41.845 23.205 ;
        RECT 39.155 21.845 41.845 22.015 ;
        RECT 41.675 20.995 41.845 22.015 ;
        RECT 39.155 22.555 41.845 22.725 ;
        RECT 40.835 22.555 41.005 23.205 ;
        RECT 40.835 20.995 41.005 22.015 ;
        RECT 39.995 22.555 40.165 23.205 ;
        RECT 39.995 20.995 40.165 22.015 ;
        RECT 39.155 21.845 39.41 22.725 ;
        RECT 39.155 20.995 39.325 23.205 ;
      LAYER met1 ;
        RECT 39.17 21.8 39.49 22.06 ;
      LAYER met2 ;
        RECT 39.2 21.77 39.46 22.09 ;
        RECT 39.26 20.84 39.4 22.09 ;
        RECT 39.03 20.84 39.4 20.98 ;
        RECT 39.03 13.7 39.17 20.98 ;
        RECT 38.8 13.7 39.17 13.84 ;
        RECT 38.8 0 38.94 13.84 ;
      LAYER via ;
        RECT 39.255 21.855 39.405 22.005 ;
      LAYER mcon ;
        RECT 39.245 21.845 39.415 22.015 ;
    END
  END out[18]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 48.575 24.905 48.745 25.925 ;
        RECT 46.055 24.195 48.745 24.365 ;
        RECT 48.575 23.715 48.745 24.365 ;
        RECT 46.055 24.905 48.745 25.075 ;
        RECT 47.735 24.905 47.905 25.925 ;
        RECT 47.735 23.715 47.905 24.365 ;
        RECT 46.895 24.905 47.065 25.925 ;
        RECT 46.895 23.715 47.065 24.365 ;
        RECT 46.055 24.565 46.315 24.735 ;
        RECT 46.055 24.195 46.31 25.075 ;
        RECT 46.055 23.715 46.225 25.925 ;
      LAYER met1 ;
        RECT 50.21 23.84 50.53 24.1 ;
        RECT 48 23.9 50.53 24.04 ;
        RECT 47.08 24.24 48.14 24.38 ;
        RECT 48 23.9 48.14 24.38 ;
        RECT 46.085 24.58 47.22 24.72 ;
        RECT 47.08 24.24 47.22 24.72 ;
        RECT 46.085 24.535 46.375 24.765 ;
      LAYER met2 ;
        RECT 50.24 23.81 50.5 24.13 ;
        RECT 50.3 17.78 50.44 24.13 ;
        RECT 49.84 17.78 50.44 17.92 ;
        RECT 49.84 8.94 49.98 17.92 ;
        RECT 48.46 8.94 49.98 9.08 ;
        RECT 48.46 0 48.6 9.08 ;
      LAYER via ;
        RECT 50.295 23.895 50.445 24.045 ;
      LAYER mcon ;
        RECT 46.145 24.565 46.315 24.735 ;
    END
  END out[19]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 64.215 17.115 64.385 17.765 ;
        RECT 61.695 16.405 64.385 16.575 ;
        RECT 64.215 15.555 64.385 16.575 ;
        RECT 61.695 17.115 64.385 17.285 ;
        RECT 63.375 17.115 63.545 17.765 ;
        RECT 63.375 15.555 63.545 16.575 ;
        RECT 62.535 17.115 62.705 17.765 ;
        RECT 62.535 15.555 62.705 16.575 ;
        RECT 61.695 16.405 61.95 17.285 ;
        RECT 61.695 15.555 61.865 17.765 ;
      LAYER met1 ;
        RECT 61.725 16.375 62.015 16.605 ;
        RECT 58.49 16.42 62.015 16.56 ;
        RECT 58.49 16.36 58.81 16.62 ;
      LAYER met2 ;
        RECT 58.52 16.33 58.78 16.65 ;
        RECT 58.12 16.42 58.78 16.56 ;
        RECT 58.12 8.94 58.26 16.56 ;
        RECT 57.66 8.94 58.26 9.08 ;
        RECT 57.66 0 57.8 9.08 ;
      LAYER via ;
        RECT 58.575 16.415 58.725 16.565 ;
      LAYER mcon ;
        RECT 61.785 16.405 61.955 16.575 ;
    END
  END out[20]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 70.155 37.315 70.325 39.525 ;
        RECT 67.635 38.875 70.325 39.045 ;
        RECT 70.07 38.165 70.325 39.045 ;
        RECT 67.635 38.165 70.325 38.335 ;
        RECT 69.315 38.875 69.485 39.525 ;
        RECT 69.315 37.315 69.485 38.335 ;
        RECT 68.475 38.875 68.645 39.525 ;
        RECT 68.475 37.315 68.645 38.335 ;
        RECT 67.635 38.875 67.805 39.525 ;
        RECT 67.635 37.315 67.805 38.335 ;
      LAYER met1 ;
        RECT 67.705 38.135 67.995 38.365 ;
        RECT 67.78 37.84 67.92 38.365 ;
        RECT 66.77 37.84 67.92 37.98 ;
        RECT 66.77 37.78 67.09 38.04 ;
      LAYER met2 ;
        RECT 66.86 31.38 67.46 31.52 ;
        RECT 67.32 12.68 67.46 31.52 ;
        RECT 66.86 9.28 67.46 9.42 ;
        RECT 67.32 0 67.46 9.42 ;
        RECT 66.86 12.68 67.46 12.82 ;
        RECT 66.8 37.75 67.06 38.07 ;
        RECT 66.86 31.38 67 38.07 ;
        RECT 66.86 9.28 67 12.82 ;
      LAYER via ;
        RECT 66.855 37.835 67.005 37.985 ;
      LAYER mcon ;
        RECT 67.765 38.165 67.935 38.335 ;
    END
  END out[21]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 81.655 10.115 81.825 12.325 ;
        RECT 79.135 11.675 81.825 11.845 ;
        RECT 81.57 10.965 81.825 11.845 ;
        RECT 79.135 10.965 81.825 11.135 ;
        RECT 80.815 11.675 80.985 12.325 ;
        RECT 80.815 10.115 80.985 11.135 ;
        RECT 79.975 11.675 80.145 12.325 ;
        RECT 79.975 10.115 80.145 11.135 ;
        RECT 79.135 11.675 79.305 12.325 ;
        RECT 79.135 10.115 79.305 11.135 ;
      LAYER met1 ;
        RECT 79.205 10.935 79.495 11.165 ;
        RECT 77.81 10.98 79.495 11.12 ;
        RECT 77.81 10.92 78.13 11.18 ;
      LAYER met2 ;
        RECT 77.84 10.89 78.1 11.21 ;
        RECT 77.9 8.94 78.04 11.21 ;
        RECT 76.52 8.94 78.04 9.08 ;
        RECT 76.52 0 76.66 9.08 ;
      LAYER via ;
        RECT 77.895 10.975 78.045 11.125 ;
      LAYER mcon ;
        RECT 79.265 10.965 79.435 11.135 ;
    END
  END out[22]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 85.835 22.555 86.005 23.205 ;
        RECT 83.315 21.845 86.005 22.015 ;
        RECT 85.835 20.995 86.005 22.015 ;
        RECT 83.315 22.555 86.005 22.725 ;
        RECT 84.995 22.555 85.165 23.205 ;
        RECT 84.995 20.995 85.165 22.015 ;
        RECT 84.155 22.555 84.325 23.205 ;
        RECT 84.155 20.995 84.325 22.015 ;
        RECT 83.315 21.845 83.57 22.725 ;
        RECT 83.315 20.995 83.485 23.205 ;
      LAYER met1 ;
        RECT 86.09 21.8 86.41 22.06 ;
        RECT 85.645 21.86 86.41 22 ;
        RECT 85.645 21.815 85.935 22.045 ;
      LAYER met2 ;
        RECT 86.18 20.5 86.78 20.64 ;
        RECT 86.64 16.42 86.78 20.64 ;
        RECT 86.18 16.42 86.78 16.56 ;
        RECT 86.12 21.77 86.38 22.09 ;
        RECT 86.18 20.5 86.32 22.09 ;
        RECT 86.18 0 86.32 16.56 ;
      LAYER via ;
        RECT 86.175 21.855 86.325 22.005 ;
      LAYER mcon ;
        RECT 85.705 21.845 85.875 22.015 ;
    END
  END out[23]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 94.995 10.115 95.165 12.325 ;
        RECT 92.475 11.675 95.165 11.845 ;
        RECT 94.91 10.965 95.165 11.845 ;
        RECT 92.475 10.965 95.165 11.135 ;
        RECT 94.155 11.675 94.325 12.325 ;
        RECT 94.155 10.115 94.325 11.135 ;
        RECT 93.315 11.675 93.485 12.325 ;
        RECT 93.315 10.115 93.485 11.135 ;
        RECT 92.475 11.675 92.645 12.325 ;
        RECT 92.475 10.115 92.645 11.135 ;
      LAYER met1 ;
        RECT 94.37 10.92 94.69 11.18 ;
      LAYER met2 ;
        RECT 95.38 0 95.52 0.485 ;
        RECT 94.46 0.17 95.52 0.31 ;
        RECT 94.4 10.89 94.66 11.21 ;
        RECT 94.46 0.17 94.6 11.21 ;
      LAYER via ;
        RECT 94.455 10.975 94.605 11.125 ;
      LAYER mcon ;
        RECT 94.445 10.965 94.615 11.135 ;
    END
  END out[24]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 107.875 10.115 108.045 12.325 ;
        RECT 105.355 11.675 108.045 11.845 ;
        RECT 107.79 10.965 108.045 11.845 ;
        RECT 105.355 10.965 108.045 11.135 ;
        RECT 107.035 11.675 107.205 12.325 ;
        RECT 107.035 10.115 107.205 11.135 ;
        RECT 106.195 11.675 106.365 12.325 ;
        RECT 106.195 10.115 106.365 11.135 ;
        RECT 105.355 11.675 105.525 12.325 ;
        RECT 105.355 10.115 105.525 11.135 ;
      LAYER met1 ;
        RECT 108.17 10.92 108.49 11.18 ;
        RECT 107.725 10.98 108.49 11.12 ;
        RECT 107.725 10.935 108.015 11.165 ;
      LAYER met2 ;
        RECT 108.2 10.89 108.46 11.21 ;
        RECT 108.26 0.78 108.4 11.21 ;
        RECT 105.04 0.78 108.4 0.92 ;
        RECT 105.04 0 105.18 0.92 ;
      LAYER via ;
        RECT 108.255 10.975 108.405 11.125 ;
      LAYER mcon ;
        RECT 107.785 10.965 107.955 11.135 ;
    END
  END out[25]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 116.615 23.715 116.785 25.925 ;
        RECT 114.095 24.905 116.785 25.075 ;
        RECT 116.53 24.195 116.785 25.075 ;
        RECT 114.095 24.195 116.785 24.365 ;
        RECT 115.775 24.905 115.945 25.925 ;
        RECT 115.775 23.715 115.945 24.365 ;
        RECT 114.935 24.905 115.105 25.925 ;
        RECT 114.935 23.715 115.105 24.365 ;
        RECT 114.095 24.905 114.265 25.925 ;
        RECT 114.095 23.715 114.265 24.365 ;
      LAYER met1 ;
        RECT 114.165 24.875 114.455 25.105 ;
        RECT 114.24 23.9 114.38 25.105 ;
        RECT 113.69 23.9 114.38 24.04 ;
        RECT 113.69 23.84 114.01 24.1 ;
      LAYER met2 ;
        RECT 113.72 23.9 114.38 24.04 ;
        RECT 114.24 0 114.38 24.04 ;
        RECT 113.72 23.81 113.98 24.13 ;
      LAYER via ;
        RECT 113.775 23.895 113.925 24.045 ;
      LAYER mcon ;
        RECT 114.225 24.905 114.395 25.075 ;
    END
  END out[26]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 122.595 10.115 122.765 12.325 ;
        RECT 120.075 11.675 122.765 11.845 ;
        RECT 122.51 10.965 122.765 11.845 ;
        RECT 120.075 10.965 122.765 11.135 ;
        RECT 121.755 11.675 121.925 12.325 ;
        RECT 121.755 10.115 121.925 11.135 ;
        RECT 120.915 11.675 121.085 12.325 ;
        RECT 120.915 10.115 121.085 11.135 ;
        RECT 120.075 11.675 120.245 12.325 ;
        RECT 120.075 10.115 120.245 11.135 ;
      LAYER met1 ;
        RECT 121.97 10.92 122.29 11.18 ;
      LAYER met2 ;
        RECT 122.06 0.78 124.04 0.92 ;
        RECT 123.9 0 124.04 0.92 ;
        RECT 122 10.89 122.26 11.21 ;
        RECT 122.06 0.78 122.2 11.21 ;
      LAYER via ;
        RECT 122.055 10.975 122.205 11.125 ;
      LAYER mcon ;
        RECT 122.045 10.965 122.215 11.135 ;
    END
  END out[27]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 137.315 10.115 137.485 12.325 ;
        RECT 134.795 11.675 137.485 11.845 ;
        RECT 137.23 10.965 137.485 11.845 ;
        RECT 134.795 10.965 137.485 11.135 ;
        RECT 136.475 11.675 136.645 12.325 ;
        RECT 136.475 10.115 136.645 11.135 ;
        RECT 135.635 11.675 135.805 12.325 ;
        RECT 135.635 10.115 135.805 11.135 ;
        RECT 134.795 11.675 134.965 12.325 ;
        RECT 134.795 10.115 134.965 11.135 ;
      LAYER met1 ;
        RECT 134.865 10.935 135.155 11.165 ;
        RECT 133.1 10.98 135.155 11.12 ;
        RECT 133.01 10.24 133.33 10.5 ;
        RECT 133.1 10.24 133.24 11.12 ;
      LAYER met2 ;
        RECT 133.04 10.21 133.3 10.53 ;
        RECT 133.1 0 133.24 10.53 ;
      LAYER via ;
        RECT 133.095 10.295 133.245 10.445 ;
      LAYER mcon ;
        RECT 134.925 10.965 135.095 11.135 ;
    END
  END out[28]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 157.555 10.115 157.725 12.325 ;
        RECT 155.035 11.675 157.725 11.845 ;
        RECT 157.47 10.965 157.725 11.845 ;
        RECT 155.035 10.965 157.725 11.135 ;
        RECT 156.715 11.675 156.885 12.325 ;
        RECT 156.715 10.115 156.885 11.135 ;
        RECT 155.875 11.675 156.045 12.325 ;
        RECT 155.875 10.115 156.045 11.135 ;
        RECT 155.035 11.675 155.205 12.325 ;
        RECT 155.035 10.115 155.205 11.135 ;
      LAYER met1 ;
        RECT 155.565 10.935 155.855 11.165 ;
        RECT 155.64 10.64 155.78 11.165 ;
        RECT 151.5 10.64 155.78 10.78 ;
        RECT 145.06 10.98 151.64 11.12 ;
        RECT 151.5 10.64 151.64 11.12 ;
        RECT 145.06 10.64 145.2 11.12 ;
        RECT 144.05 10.64 145.2 10.78 ;
        RECT 144.05 10.58 144.37 10.84 ;
      LAYER met2 ;
        RECT 144.08 10.55 144.34 10.87 ;
        RECT 144.14 1.46 144.28 10.87 ;
        RECT 142.76 1.46 144.28 1.6 ;
        RECT 142.76 0 142.9 1.6 ;
      LAYER via ;
        RECT 144.135 10.635 144.285 10.785 ;
      LAYER mcon ;
        RECT 155.625 10.965 155.795 11.135 ;
    END
  END out[29]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 172.275 10.115 172.445 12.325 ;
        RECT 169.755 11.675 172.445 11.845 ;
        RECT 172.19 10.965 172.445 11.845 ;
        RECT 172.185 11.305 172.445 11.475 ;
        RECT 169.755 10.965 172.445 11.135 ;
        RECT 171.435 11.675 171.605 12.325 ;
        RECT 171.435 10.115 171.605 11.135 ;
        RECT 170.595 11.675 170.765 12.325 ;
        RECT 170.595 10.115 170.765 11.135 ;
        RECT 169.755 11.675 169.925 12.325 ;
        RECT 169.755 10.115 169.925 11.135 ;
      LAYER met1 ;
        RECT 172.125 11.275 172.415 11.505 ;
        RECT 171.65 11.32 172.415 11.46 ;
        RECT 171.65 11.26 171.97 11.52 ;
        RECT 171.65 8.2 171.97 8.46 ;
        RECT 151.87 8.26 171.97 8.4 ;
        RECT 151.87 8.2 152.19 8.46 ;
      LAYER met2 ;
        RECT 171.68 11.23 171.94 11.55 ;
        RECT 171.68 8.17 171.94 8.49 ;
        RECT 171.74 8.17 171.88 11.55 ;
        RECT 151.9 8.17 152.16 8.49 ;
        RECT 151.96 0 152.1 8.49 ;
      LAYER via ;
        RECT 151.955 8.255 152.105 8.405 ;
        RECT 171.735 11.315 171.885 11.465 ;
        RECT 171.735 8.255 171.885 8.405 ;
      LAYER mcon ;
        RECT 172.185 11.305 172.355 11.475 ;
    END
  END out[30]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 181.475 10.115 181.645 12.325 ;
        RECT 178.955 11.675 181.645 11.845 ;
        RECT 181.39 10.965 181.645 11.845 ;
        RECT 178.955 10.965 181.645 11.135 ;
        RECT 180.635 11.675 180.805 12.325 ;
        RECT 180.635 10.115 180.805 11.135 ;
        RECT 179.795 11.675 179.965 12.325 ;
        RECT 179.795 10.115 179.965 11.135 ;
        RECT 178.955 11.675 179.125 12.325 ;
        RECT 178.955 10.115 179.125 11.135 ;
      LAYER met1 ;
        RECT 179.025 10.935 179.315 11.165 ;
        RECT 164.84 10.98 179.315 11.12 ;
        RECT 164.84 10.47 164.98 11.12 ;
        RECT 161.62 10.47 164.98 10.61 ;
        RECT 161.62 10.3 161.76 10.61 ;
        RECT 160.61 10.3 161.76 10.44 ;
        RECT 160.61 10.24 160.93 10.5 ;
      LAYER met2 ;
        RECT 161.16 8.94 161.76 9.08 ;
        RECT 161.62 0 161.76 9.08 ;
        RECT 160.64 10.3 161.3 10.44 ;
        RECT 161.16 8.94 161.3 10.44 ;
        RECT 160.64 10.21 160.9 10.53 ;
      LAYER via ;
        RECT 160.695 10.295 160.845 10.445 ;
      LAYER mcon ;
        RECT 179.085 10.965 179.255 11.135 ;
    END
  END out[31]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 182.725 11.225 183.065 11.595 ;
        RECT 144.065 22.105 144.42 22.475 ;
      LAYER met1 ;
        RECT 182.69 11.26 183.01 11.52 ;
        RECT 178.64 11.32 183.01 11.46 ;
        RECT 162.54 11.66 178.78 11.8 ;
        RECT 178.64 11.32 178.78 11.8 ;
        RECT 159.32 11.83 162.68 11.97 ;
        RECT 162.54 11.66 162.68 11.97 ;
        RECT 159.32 11.66 159.46 11.97 ;
        RECT 157.02 11.66 159.46 11.8 ;
        RECT 152.88 11.83 157.16 11.97 ;
        RECT 157.02 11.66 157.16 11.97 ;
        RECT 151.5 12 153.02 12.14 ;
        RECT 152.88 11.83 153.02 12.14 ;
        RECT 151.5 11.66 151.64 12.14 ;
        RECT 145.06 11.66 151.64 11.8 ;
        RECT 144.05 12 145.2 12.14 ;
        RECT 145.06 11.66 145.2 12.14 ;
        RECT 144.05 11.94 144.37 12.2 ;
        RECT 144.05 22.14 144.37 22.4 ;
      LAYER met2 ;
        RECT 182.72 11.23 182.98 11.55 ;
        RECT 182.78 0.78 182.92 11.55 ;
        RECT 180.48 0.78 182.92 0.92 ;
        RECT 180.48 0 180.62 0.92 ;
        RECT 144.08 22.11 144.34 22.43 ;
        RECT 144.08 11.91 144.34 12.23 ;
        RECT 144.14 11.91 144.28 22.43 ;
      LAYER via ;
        RECT 144.135 22.195 144.285 22.345 ;
        RECT 144.135 11.995 144.285 12.145 ;
        RECT 182.775 11.315 182.925 11.465 ;
      LAYER mcon ;
        RECT 144.125 22.185 144.295 22.355 ;
        RECT 182.765 11.305 182.935 11.475 ;
    END
  END rst
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 10.185 1.325 10.515 1.655 ;
        RECT 10.2 0 10.5 1.655 ;
      LAYER li1 ;
        RECT 20.015 10.115 20.185 12.325 ;
        RECT 17.495 11.675 20.185 11.845 ;
        RECT 19.93 10.965 20.185 11.845 ;
        RECT 17.495 10.965 20.185 11.135 ;
        RECT 19.175 11.675 19.345 12.325 ;
        RECT 19.175 10.115 19.345 11.135 ;
        RECT 18.335 11.675 18.505 12.325 ;
        RECT 18.335 10.115 18.505 11.135 ;
        RECT 17.495 11.675 17.665 12.325 ;
        RECT 17.495 10.115 17.665 11.135 ;
      LAYER met1 ;
        RECT 17.565 10.935 17.855 11.165 ;
        RECT 17.09 10.98 17.855 11.12 ;
        RECT 17.09 10.92 17.41 11.18 ;
      LAYER met3 ;
        RECT 17.085 1.325 17.415 1.655 ;
        RECT 10.16 1.34 17.415 1.64 ;
        RECT 10.16 1.33 10.54 1.65 ;
      LAYER met2 ;
        RECT 17.11 1.305 17.39 1.675 ;
        RECT 17.12 10.89 17.38 11.21 ;
        RECT 17.18 1.305 17.32 11.21 ;
      LAYER via ;
        RECT 17.175 10.975 17.325 11.125 ;
      LAYER via2 ;
        RECT 17.15 1.39 17.35 1.59 ;
      LAYER mcon ;
        RECT 17.625 10.965 17.795 11.135 ;
      LAYER via3 ;
        RECT 10.25 1.39 10.45 1.59 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.525 1.935 138.855 2.265 ;
        RECT 138.54 0 138.84 2.265 ;
      LAYER li1 ;
        RECT 142.835 12.835 143.005 15.045 ;
        RECT 140.315 14.025 143.005 14.195 ;
        RECT 142.75 13.315 143.005 14.195 ;
        RECT 140.315 13.315 143.005 13.485 ;
        RECT 141.995 14.025 142.165 15.045 ;
        RECT 141.995 12.835 142.165 13.485 ;
        RECT 141.155 14.025 141.325 15.045 ;
        RECT 141.155 12.835 141.325 13.485 ;
        RECT 140.315 14.025 140.485 15.045 ;
        RECT 140.315 12.835 140.485 13.485 ;
      LAYER met1 ;
        RECT 141.29 13.98 141.61 14.24 ;
      LAYER met3 ;
        RECT 141.285 1.935 141.615 2.265 ;
        RECT 138.5 1.95 141.615 2.25 ;
        RECT 138.5 1.94 138.88 2.26 ;
      LAYER met2 ;
        RECT 141.31 1.915 141.59 2.285 ;
        RECT 141.32 13.95 141.58 14.27 ;
        RECT 141.38 1.915 141.52 14.27 ;
      LAYER via ;
        RECT 141.375 14.035 141.525 14.185 ;
      LAYER via2 ;
        RECT 141.35 2 141.55 2.2 ;
      LAYER mcon ;
        RECT 141.365 14.025 141.535 14.195 ;
      LAYER via3 ;
        RECT 138.59 2 138.79 2.2 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.635 20.845 151.965 21.175 ;
        RECT 151.65 19.03 151.95 21.175 ;
        RECT 150.96 8.66 151.95 8.96 ;
        RECT 151.65 0 151.95 8.96 ;
        RECT 150.96 19.03 151.95 19.33 ;
        RECT 150.96 8.66 151.26 19.33 ;
      LAYER li1 ;
        RECT 153.455 22.555 153.625 23.205 ;
        RECT 150.935 21.845 153.625 22.015 ;
        RECT 153.455 20.995 153.625 22.015 ;
        RECT 150.935 22.555 153.625 22.725 ;
        RECT 152.615 22.555 152.785 23.205 ;
        RECT 152.615 20.995 152.785 22.015 ;
        RECT 151.775 22.555 151.945 23.205 ;
        RECT 151.775 20.995 151.945 22.015 ;
        RECT 150.935 21.845 151.19 22.725 ;
        RECT 150.935 20.995 151.105 23.205 ;
      LAYER met1 ;
        RECT 152.33 21.8 152.65 22.06 ;
      LAYER met3 ;
        RECT 152.325 20.845 152.655 21.175 ;
        RECT 151.61 20.86 152.655 21.16 ;
        RECT 151.61 20.85 151.99 21.17 ;
      LAYER met2 ;
        RECT 152.35 20.825 152.63 21.195 ;
        RECT 152.36 21.77 152.62 22.09 ;
        RECT 152.42 20.825 152.56 22.09 ;
      LAYER via ;
        RECT 152.415 21.855 152.565 22.005 ;
      LAYER via2 ;
        RECT 152.39 20.91 152.59 21.11 ;
      LAYER mcon ;
        RECT 152.405 21.845 152.575 22.015 ;
      LAYER via3 ;
        RECT 151.7 20.91 151.9 21.11 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 164.055 1.935 164.385 2.265 ;
        RECT 164.07 0 164.37 2.265 ;
      LAYER li1 ;
        RECT 166.755 10.115 166.925 12.325 ;
        RECT 164.235 11.675 166.925 11.845 ;
        RECT 166.67 10.965 166.925 11.845 ;
        RECT 164.235 10.965 166.925 11.135 ;
        RECT 165.915 11.675 166.085 12.325 ;
        RECT 165.915 10.115 166.085 11.135 ;
        RECT 165.075 11.675 165.245 12.325 ;
        RECT 165.075 10.115 165.245 11.135 ;
        RECT 164.235 11.675 164.405 12.325 ;
        RECT 164.235 10.115 164.405 11.135 ;
      LAYER met1 ;
        RECT 164.305 10.935 164.595 11.165 ;
        RECT 163.37 10.98 164.595 11.12 ;
        RECT 163.37 10.92 163.69 11.18 ;
      LAYER met3 ;
        RECT 164.03 1.94 164.41 2.26 ;
        RECT 163.365 1.95 164.41 2.25 ;
        RECT 163.365 1.935 163.695 2.265 ;
      LAYER met2 ;
        RECT 163.39 1.915 163.67 2.285 ;
        RECT 163.4 10.89 163.66 11.21 ;
        RECT 163.46 1.915 163.6 11.21 ;
      LAYER via ;
        RECT 163.455 10.975 163.605 11.125 ;
      LAYER via2 ;
        RECT 163.43 2 163.63 2.2 ;
      LAYER mcon ;
        RECT 164.365 10.965 164.535 11.135 ;
      LAYER via3 ;
        RECT 164.12 2 164.32 2.2 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 177.165 1.935 177.495 2.265 ;
        RECT 177.18 0 177.48 2.265 ;
      LAYER li1 ;
        RECT 175.495 20.995 175.665 23.205 ;
        RECT 172.975 22.555 175.665 22.725 ;
        RECT 175.41 21.845 175.665 22.725 ;
        RECT 172.975 21.845 175.665 22.015 ;
        RECT 174.655 22.555 174.825 23.205 ;
        RECT 174.655 20.995 174.825 22.015 ;
        RECT 173.815 22.555 173.985 23.205 ;
        RECT 173.815 20.995 173.985 22.015 ;
        RECT 172.975 22.555 173.145 23.205 ;
        RECT 172.975 20.995 173.145 22.015 ;
      LAYER met1 ;
        RECT 174.41 21.8 174.73 22.06 ;
      LAYER met3 ;
        RECT 177.14 1.94 177.52 2.26 ;
        RECT 174.405 1.95 177.52 2.25 ;
        RECT 174.405 1.935 174.735 2.265 ;
      LAYER met2 ;
        RECT 174.43 1.915 174.71 2.285 ;
        RECT 174.44 21.77 174.7 22.09 ;
        RECT 174.5 1.915 174.64 22.09 ;
      LAYER via ;
        RECT 174.495 21.855 174.645 22.005 ;
      LAYER via2 ;
        RECT 174.47 2 174.67 2.2 ;
      LAYER mcon ;
        RECT 174.485 21.845 174.655 22.015 ;
      LAYER via3 ;
        RECT 177.23 2 177.43 2.2 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 189.585 6.205 189.915 6.535 ;
        RECT 189.6 0 189.9 6.535 ;
      LAYER li1 ;
        RECT 175.495 29.155 175.665 31.365 ;
        RECT 172.975 30.345 175.665 30.515 ;
        RECT 175.41 29.635 175.665 30.515 ;
        RECT 175.405 29.635 175.665 29.835 ;
        RECT 172.975 29.635 175.665 29.805 ;
        RECT 174.655 30.345 174.825 31.365 ;
        RECT 174.655 29.155 174.825 29.805 ;
        RECT 173.815 30.345 173.985 31.365 ;
        RECT 173.815 29.155 173.985 29.805 ;
        RECT 172.975 30.345 173.145 31.365 ;
        RECT 172.975 29.155 173.145 29.805 ;
      LAYER met1 ;
        RECT 185.45 29.62 185.77 29.88 ;
        RECT 184.62 29.68 185.77 29.82 ;
        RECT 176.34 30.02 184.76 30.16 ;
        RECT 184.62 29.68 184.76 30.16 ;
        RECT 176.34 29.68 176.48 30.16 ;
        RECT 175.345 29.68 176.48 29.82 ;
        RECT 175.345 29.635 175.635 29.865 ;
      LAYER met3 ;
        RECT 189.56 6.21 189.94 6.53 ;
        RECT 185.445 6.22 189.94 6.52 ;
        RECT 185.445 6.205 185.775 6.535 ;
      LAYER met2 ;
        RECT 185.47 6.185 185.75 6.555 ;
        RECT 185.48 29.59 185.74 29.91 ;
        RECT 185.54 6.185 185.68 29.91 ;
      LAYER via ;
        RECT 185.535 29.675 185.685 29.825 ;
      LAYER via2 ;
        RECT 185.51 6.27 185.71 6.47 ;
      LAYER mcon ;
        RECT 175.405 29.665 175.575 29.835 ;
      LAYER via3 ;
        RECT 189.65 6.27 189.85 6.47 ;
    END
  END out[14]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.295 1.325 23.625 1.655 ;
        RECT 23.31 0 23.61 1.655 ;
      LAYER li1 ;
        RECT 28.295 10.115 28.465 12.325 ;
        RECT 25.775 11.675 28.465 11.845 ;
        RECT 28.21 10.965 28.465 11.845 ;
        RECT 25.775 10.965 28.465 11.135 ;
        RECT 27.455 11.675 27.625 12.325 ;
        RECT 27.455 10.115 27.625 11.135 ;
        RECT 26.615 11.675 26.785 12.325 ;
        RECT 26.615 10.115 26.785 11.135 ;
        RECT 25.775 11.675 25.945 12.325 ;
        RECT 25.775 10.115 25.945 11.135 ;
      LAYER met1 ;
        RECT 25.845 10.935 26.135 11.165 ;
        RECT 25.37 10.98 26.135 11.12 ;
        RECT 25.37 10.92 25.69 11.18 ;
      LAYER met3 ;
        RECT 25.365 1.325 25.695 1.655 ;
        RECT 23.27 1.34 25.695 1.64 ;
        RECT 23.27 1.33 23.65 1.65 ;
      LAYER met2 ;
        RECT 25.39 1.305 25.67 1.675 ;
        RECT 25.4 10.89 25.66 11.21 ;
        RECT 25.46 1.305 25.6 11.21 ;
      LAYER via ;
        RECT 25.455 10.975 25.605 11.125 ;
      LAYER via2 ;
        RECT 25.43 1.39 25.63 1.59 ;
      LAYER mcon ;
        RECT 25.905 10.965 26.075 11.135 ;
      LAYER via3 ;
        RECT 23.36 1.39 23.56 1.59 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.405 8.645 36.735 8.975 ;
        RECT 36.42 0 36.72 8.975 ;
      LAYER li1 ;
        RECT 41.175 10.115 41.345 12.325 ;
        RECT 38.655 11.675 41.345 11.845 ;
        RECT 41.09 10.965 41.345 11.845 ;
        RECT 38.655 10.965 41.345 11.135 ;
        RECT 40.335 11.675 40.505 12.325 ;
        RECT 40.335 10.115 40.505 11.135 ;
        RECT 39.495 11.675 39.665 12.325 ;
        RECT 39.495 10.115 39.665 11.135 ;
        RECT 38.655 11.675 38.825 12.325 ;
        RECT 38.655 10.115 38.825 11.135 ;
      LAYER met1 ;
        RECT 39.17 10.92 39.49 11.18 ;
      LAYER met3 ;
        RECT 39.165 10.475 39.495 10.805 ;
        RECT 37.8 10.49 39.495 10.79 ;
        RECT 37.8 8.66 38.1 10.79 ;
        RECT 36.38 8.66 38.1 8.96 ;
        RECT 36.38 8.65 36.76 8.97 ;
      LAYER met2 ;
        RECT 39.19 10.455 39.47 11.21 ;
      LAYER via ;
        RECT 39.255 10.975 39.405 11.125 ;
      LAYER via2 ;
        RECT 39.23 10.54 39.43 10.74 ;
      LAYER mcon ;
        RECT 39.245 10.965 39.415 11.135 ;
      LAYER via3 ;
        RECT 36.47 8.71 36.67 8.91 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.825 2.545 49.155 2.875 ;
        RECT 48.84 0 49.14 2.875 ;
      LAYER li1 ;
        RECT 51.295 10.115 51.465 12.325 ;
        RECT 48.775 11.675 51.465 11.845 ;
        RECT 51.21 10.965 51.465 11.845 ;
        RECT 51.205 11.305 51.465 11.475 ;
        RECT 48.775 10.965 51.465 11.135 ;
        RECT 50.455 11.675 50.625 12.325 ;
        RECT 50.455 10.115 50.625 11.135 ;
        RECT 49.615 11.675 49.785 12.325 ;
        RECT 49.615 10.115 49.785 11.135 ;
        RECT 48.775 11.675 48.945 12.325 ;
        RECT 48.775 10.115 48.945 11.135 ;
      LAYER met1 ;
        RECT 51.145 11.275 51.435 11.505 ;
        RECT 50.21 11.32 51.435 11.46 ;
        RECT 50.21 11.26 50.53 11.52 ;
      LAYER met3 ;
        RECT 50.205 2.545 50.535 2.875 ;
        RECT 48.8 2.56 50.535 2.86 ;
        RECT 48.8 2.55 49.18 2.87 ;
      LAYER met2 ;
        RECT 50.23 2.525 50.51 2.895 ;
        RECT 50.24 11.23 50.5 11.55 ;
        RECT 50.3 2.525 50.44 11.55 ;
      LAYER via ;
        RECT 50.295 11.315 50.445 11.465 ;
      LAYER via2 ;
        RECT 50.27 2.61 50.47 2.81 ;
      LAYER mcon ;
        RECT 51.205 11.305 51.375 11.475 ;
      LAYER via3 ;
        RECT 48.89 2.61 49.09 2.81 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.935 1.325 62.265 1.655 ;
        RECT 61.95 0 62.25 1.655 ;
      LAYER li1 ;
        RECT 64.635 10.115 64.805 12.325 ;
        RECT 62.115 11.675 64.805 11.845 ;
        RECT 64.55 10.965 64.805 11.845 ;
        RECT 62.115 10.965 64.805 11.135 ;
        RECT 63.795 11.675 63.965 12.325 ;
        RECT 63.795 10.115 63.965 11.135 ;
        RECT 62.955 11.675 63.125 12.325 ;
        RECT 62.955 10.115 63.125 11.135 ;
        RECT 62.115 11.675 62.285 12.325 ;
        RECT 62.115 10.115 62.285 11.135 ;
      LAYER met1 ;
        RECT 64.01 10.92 64.33 11.18 ;
      LAYER met3 ;
        RECT 64.005 1.325 64.335 1.655 ;
        RECT 61.91 1.34 64.335 1.64 ;
        RECT 61.91 1.33 62.29 1.65 ;
      LAYER met2 ;
        RECT 64.03 1.305 64.31 1.675 ;
        RECT 64.04 10.89 64.3 11.21 ;
        RECT 64.1 1.305 64.24 11.21 ;
      LAYER via ;
        RECT 64.095 10.975 64.245 11.125 ;
      LAYER via2 ;
        RECT 64.07 1.39 64.27 1.59 ;
      LAYER mcon ;
        RECT 64.085 10.965 64.255 11.135 ;
      LAYER via3 ;
        RECT 62 1.39 62.2 1.59 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.355 1.325 74.685 1.655 ;
        RECT 74.37 0 74.67 1.655 ;
      LAYER li1 ;
        RECT 72.455 10.115 72.625 12.325 ;
        RECT 69.935 11.675 72.625 11.845 ;
        RECT 72.37 10.965 72.625 11.845 ;
        RECT 69.935 10.965 72.625 11.135 ;
        RECT 71.615 11.675 71.785 12.325 ;
        RECT 71.615 10.115 71.785 11.135 ;
        RECT 70.775 11.675 70.945 12.325 ;
        RECT 70.775 10.115 70.945 11.135 ;
        RECT 69.935 11.675 70.105 12.325 ;
        RECT 69.935 10.115 70.105 11.135 ;
      LAYER met1 ;
        RECT 72.29 10.92 72.61 11.18 ;
      LAYER met3 ;
        RECT 74.33 1.33 74.71 1.65 ;
        RECT 72.285 1.34 74.71 1.64 ;
        RECT 72.285 1.325 72.615 1.655 ;
      LAYER met2 ;
        RECT 72.31 1.305 72.59 1.675 ;
        RECT 72.32 10.89 72.58 11.21 ;
        RECT 72.38 1.305 72.52 11.21 ;
      LAYER via ;
        RECT 72.375 10.975 72.525 11.125 ;
      LAYER via2 ;
        RECT 72.35 1.39 72.55 1.59 ;
      LAYER mcon ;
        RECT 72.365 10.965 72.535 11.135 ;
      LAYER via3 ;
        RECT 74.42 1.39 74.62 1.59 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.465 1.325 87.795 1.655 ;
        RECT 87.48 0 87.78 1.655 ;
      LAYER li1 ;
        RECT 87.175 10.115 87.345 12.325 ;
        RECT 84.655 11.675 87.345 11.845 ;
        RECT 87.09 10.965 87.345 11.845 ;
        RECT 84.655 10.965 87.345 11.135 ;
        RECT 86.335 11.675 86.505 12.325 ;
        RECT 86.335 10.115 86.505 11.135 ;
        RECT 85.495 11.675 85.665 12.325 ;
        RECT 85.495 10.115 85.665 11.135 ;
        RECT 84.655 11.675 84.825 12.325 ;
        RECT 84.655 10.115 84.825 11.135 ;
      LAYER met1 ;
        RECT 88.85 10.92 89.17 11.18 ;
        RECT 87.025 10.98 89.17 11.12 ;
        RECT 87.025 10.935 87.315 11.165 ;
      LAYER met3 ;
        RECT 88.845 1.325 89.175 1.655 ;
        RECT 87.44 1.34 89.175 1.64 ;
        RECT 87.44 1.33 87.82 1.65 ;
      LAYER met2 ;
        RECT 88.87 1.305 89.15 1.675 ;
        RECT 88.88 10.89 89.14 11.21 ;
        RECT 88.94 1.305 89.08 11.21 ;
      LAYER via ;
        RECT 88.935 10.975 89.085 11.125 ;
      LAYER via2 ;
        RECT 88.91 1.39 89.11 1.59 ;
      LAYER mcon ;
        RECT 87.085 10.965 87.255 11.135 ;
      LAYER via3 ;
        RECT 87.53 1.39 87.73 1.59 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.885 8.645 100.215 8.975 ;
        RECT 99.9 0 100.2 8.975 ;
      LAYER li1 ;
        RECT 101.435 10.115 101.605 12.325 ;
        RECT 98.915 11.675 101.605 11.845 ;
        RECT 101.35 10.965 101.605 11.845 ;
        RECT 98.915 10.965 101.605 11.135 ;
        RECT 100.595 11.675 100.765 12.325 ;
        RECT 100.595 10.115 100.765 11.135 ;
        RECT 99.755 11.675 99.925 12.325 ;
        RECT 99.755 10.115 99.925 11.135 ;
        RECT 98.915 11.675 99.085 12.325 ;
        RECT 98.915 10.115 99.085 11.135 ;
      LAYER met1 ;
        RECT 99.905 10.935 100.195 11.165 ;
        RECT 99.92 10.89 100.18 11.21 ;
      LAYER met3 ;
        RECT 99.86 8.65 100.24 8.97 ;
        RECT 99.885 8.645 100.215 8.975 ;
        RECT 99.44 8.66 100.24 8.96 ;
      LAYER met2 ;
        RECT 99.89 10.92 100.21 11.18 ;
        RECT 99.91 8.625 100.19 8.995 ;
        RECT 99.98 8.625 100.12 11.18 ;
      LAYER via ;
        RECT 99.975 10.975 100.125 11.125 ;
      LAYER via2 ;
        RECT 99.95 8.71 100.15 8.91 ;
      LAYER mcon ;
        RECT 99.965 10.965 100.135 11.135 ;
      LAYER via3 ;
        RECT 99.95 8.71 100.15 8.91 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.995 9.255 113.325 9.585 ;
        RECT 113.01 0 113.31 9.585 ;
      LAYER li1 ;
        RECT 113.435 11.675 113.605 12.325 ;
        RECT 110.915 10.965 113.605 11.135 ;
        RECT 113.435 10.115 113.605 11.135 ;
        RECT 110.915 11.675 113.605 11.845 ;
        RECT 112.595 11.675 112.765 12.325 ;
        RECT 112.595 10.115 112.765 11.135 ;
        RECT 111.755 11.675 111.925 12.325 ;
        RECT 111.755 10.115 111.925 11.135 ;
        RECT 110.915 10.965 111.17 11.845 ;
        RECT 110.915 10.115 111.085 12.325 ;
      LAYER met1 ;
        RECT 113.69 10.92 114.01 11.18 ;
        RECT 113.245 10.98 114.01 11.12 ;
        RECT 113.245 10.935 113.535 11.165 ;
      LAYER met3 ;
        RECT 113.225 9.255 113.555 9.585 ;
        RECT 112.97 9.26 113.555 9.58 ;
        RECT 112.755 9.27 113.555 9.57 ;
      LAYER met2 ;
        RECT 113.72 10.89 113.98 11.21 ;
        RECT 113.32 10.98 113.98 11.12 ;
        RECT 113.25 9.235 113.53 9.605 ;
        RECT 113.32 9.235 113.46 11.12 ;
      LAYER via ;
        RECT 113.775 10.975 113.925 11.125 ;
      LAYER via2 ;
        RECT 113.29 9.32 113.49 9.52 ;
      LAYER mcon ;
        RECT 113.305 10.965 113.475 11.135 ;
      LAYER via3 ;
        RECT 113.06 9.32 113.26 9.52 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 126.105 1.325 126.435 1.655 ;
        RECT 126.12 0 126.42 1.655 ;
      LAYER li1 ;
        RECT 128.575 10.115 128.745 12.325 ;
        RECT 126.055 11.675 128.745 11.845 ;
        RECT 128.49 10.965 128.745 11.845 ;
        RECT 126.055 10.965 128.745 11.135 ;
        RECT 127.735 11.675 127.905 12.325 ;
        RECT 127.735 10.115 127.905 11.135 ;
        RECT 126.895 11.675 127.065 12.325 ;
        RECT 126.895 10.115 127.065 11.135 ;
        RECT 126.055 11.675 126.225 12.325 ;
        RECT 126.055 10.115 126.225 11.135 ;
      LAYER met1 ;
        RECT 127.49 10.92 127.81 11.18 ;
      LAYER met3 ;
        RECT 127.485 1.325 127.815 1.655 ;
        RECT 126.08 1.34 127.815 1.64 ;
        RECT 126.08 1.33 126.46 1.65 ;
      LAYER met2 ;
        RECT 127.51 1.305 127.79 1.675 ;
        RECT 127.52 10.89 127.78 11.21 ;
        RECT 127.58 1.305 127.72 11.21 ;
      LAYER via ;
        RECT 127.575 10.975 127.725 11.125 ;
      LAYER via2 ;
        RECT 127.55 1.39 127.75 1.59 ;
      LAYER mcon ;
        RECT 127.565 10.965 127.735 11.135 ;
      LAYER via3 ;
        RECT 126.17 1.39 126.37 1.59 ;
    END
  END out[9]
  OBS
    LAYER mcon ;
      RECT 189.665 9.775 189.835 9.945 ;
      RECT 189.665 12.495 189.835 12.665 ;
      RECT 189.665 15.215 189.835 15.385 ;
      RECT 189.665 17.935 189.835 18.105 ;
      RECT 189.665 20.655 189.835 20.825 ;
      RECT 189.665 23.375 189.835 23.545 ;
      RECT 189.665 26.095 189.835 26.265 ;
      RECT 189.665 28.815 189.835 28.985 ;
      RECT 189.665 31.535 189.835 31.705 ;
      RECT 189.665 34.255 189.835 34.425 ;
      RECT 189.665 36.975 189.835 37.145 ;
      RECT 189.665 39.695 189.835 39.865 ;
      RECT 189.665 42.415 189.835 42.585 ;
      RECT 189.665 45.135 189.835 45.305 ;
      RECT 189.665 47.855 189.835 48.025 ;
      RECT 189.665 50.575 189.835 50.745 ;
      RECT 189.665 53.295 189.835 53.465 ;
      RECT 189.665 56.015 189.835 56.185 ;
      RECT 189.665 58.735 189.835 58.905 ;
      RECT 189.205 9.775 189.375 9.945 ;
      RECT 189.205 12.495 189.375 12.665 ;
      RECT 189.205 15.215 189.375 15.385 ;
      RECT 189.205 17.935 189.375 18.105 ;
      RECT 189.205 20.655 189.375 20.825 ;
      RECT 189.205 23.375 189.375 23.545 ;
      RECT 189.205 26.095 189.375 26.265 ;
      RECT 189.205 28.815 189.375 28.985 ;
      RECT 189.205 31.535 189.375 31.705 ;
      RECT 189.205 34.255 189.375 34.425 ;
      RECT 189.205 36.975 189.375 37.145 ;
      RECT 189.205 39.695 189.375 39.865 ;
      RECT 189.205 42.415 189.375 42.585 ;
      RECT 189.205 45.135 189.375 45.305 ;
      RECT 189.205 47.855 189.375 48.025 ;
      RECT 189.205 50.575 189.375 50.745 ;
      RECT 189.205 53.295 189.375 53.465 ;
      RECT 189.205 56.015 189.375 56.185 ;
      RECT 189.205 58.735 189.375 58.905 ;
      RECT 188.745 9.775 188.915 9.945 ;
      RECT 188.745 12.495 188.915 12.665 ;
      RECT 188.745 15.215 188.915 15.385 ;
      RECT 188.745 17.935 188.915 18.105 ;
      RECT 188.745 20.655 188.915 20.825 ;
      RECT 188.745 23.375 188.915 23.545 ;
      RECT 188.745 26.095 188.915 26.265 ;
      RECT 188.745 28.815 188.915 28.985 ;
      RECT 188.745 31.535 188.915 31.705 ;
      RECT 188.745 34.255 188.915 34.425 ;
      RECT 188.745 36.975 188.915 37.145 ;
      RECT 188.745 39.695 188.915 39.865 ;
      RECT 188.745 42.415 188.915 42.585 ;
      RECT 188.745 45.135 188.915 45.305 ;
      RECT 188.745 47.855 188.915 48.025 ;
      RECT 188.745 50.575 188.915 50.745 ;
      RECT 188.745 53.295 188.915 53.465 ;
      RECT 188.745 56.015 188.915 56.185 ;
      RECT 188.745 58.735 188.915 58.905 ;
      RECT 188.285 9.775 188.455 9.945 ;
      RECT 188.285 12.495 188.455 12.665 ;
      RECT 188.285 15.215 188.455 15.385 ;
      RECT 188.285 17.935 188.455 18.105 ;
      RECT 188.285 20.655 188.455 20.825 ;
      RECT 188.285 23.375 188.455 23.545 ;
      RECT 188.285 26.095 188.455 26.265 ;
      RECT 188.285 28.815 188.455 28.985 ;
      RECT 188.285 31.535 188.455 31.705 ;
      RECT 188.285 34.255 188.455 34.425 ;
      RECT 188.285 36.975 188.455 37.145 ;
      RECT 188.285 39.695 188.455 39.865 ;
      RECT 188.285 42.415 188.455 42.585 ;
      RECT 188.285 45.135 188.455 45.305 ;
      RECT 188.285 47.855 188.455 48.025 ;
      RECT 188.285 50.575 188.455 50.745 ;
      RECT 188.285 53.295 188.455 53.465 ;
      RECT 188.285 56.015 188.455 56.185 ;
      RECT 188.285 58.735 188.455 58.905 ;
      RECT 187.825 9.775 187.995 9.945 ;
      RECT 187.825 12.495 187.995 12.665 ;
      RECT 187.825 15.215 187.995 15.385 ;
      RECT 187.825 17.935 187.995 18.105 ;
      RECT 187.825 20.655 187.995 20.825 ;
      RECT 187.825 23.375 187.995 23.545 ;
      RECT 187.825 26.095 187.995 26.265 ;
      RECT 187.825 28.815 187.995 28.985 ;
      RECT 187.825 31.535 187.995 31.705 ;
      RECT 187.825 34.255 187.995 34.425 ;
      RECT 187.825 36.975 187.995 37.145 ;
      RECT 187.825 39.695 187.995 39.865 ;
      RECT 187.825 42.415 187.995 42.585 ;
      RECT 187.825 45.135 187.995 45.305 ;
      RECT 187.825 47.855 187.995 48.025 ;
      RECT 187.825 50.575 187.995 50.745 ;
      RECT 187.825 53.295 187.995 53.465 ;
      RECT 187.825 56.015 187.995 56.185 ;
      RECT 187.825 58.735 187.995 58.905 ;
      RECT 187.365 9.775 187.535 9.945 ;
      RECT 187.365 12.495 187.535 12.665 ;
      RECT 187.365 15.215 187.535 15.385 ;
      RECT 187.365 17.935 187.535 18.105 ;
      RECT 187.365 20.655 187.535 20.825 ;
      RECT 187.365 23.375 187.535 23.545 ;
      RECT 187.365 26.095 187.535 26.265 ;
      RECT 187.365 28.815 187.535 28.985 ;
      RECT 187.365 31.535 187.535 31.705 ;
      RECT 187.365 34.255 187.535 34.425 ;
      RECT 187.365 36.975 187.535 37.145 ;
      RECT 187.365 39.695 187.535 39.865 ;
      RECT 187.365 42.415 187.535 42.585 ;
      RECT 187.365 45.135 187.535 45.305 ;
      RECT 187.365 47.855 187.535 48.025 ;
      RECT 187.365 50.575 187.535 50.745 ;
      RECT 187.365 53.295 187.535 53.465 ;
      RECT 187.365 56.015 187.535 56.185 ;
      RECT 187.365 58.735 187.535 58.905 ;
      RECT 186.905 9.775 187.075 9.945 ;
      RECT 186.905 12.495 187.075 12.665 ;
      RECT 186.905 15.215 187.075 15.385 ;
      RECT 186.905 17.935 187.075 18.105 ;
      RECT 186.905 20.655 187.075 20.825 ;
      RECT 186.905 23.375 187.075 23.545 ;
      RECT 186.905 26.095 187.075 26.265 ;
      RECT 186.905 28.815 187.075 28.985 ;
      RECT 186.905 31.535 187.075 31.705 ;
      RECT 186.905 34.255 187.075 34.425 ;
      RECT 186.905 36.975 187.075 37.145 ;
      RECT 186.905 39.695 187.075 39.865 ;
      RECT 186.905 42.415 187.075 42.585 ;
      RECT 186.905 45.135 187.075 45.305 ;
      RECT 186.905 47.855 187.075 48.025 ;
      RECT 186.905 50.575 187.075 50.745 ;
      RECT 186.905 53.295 187.075 53.465 ;
      RECT 186.905 56.015 187.075 56.185 ;
      RECT 186.905 58.735 187.075 58.905 ;
      RECT 186.445 9.775 186.615 9.945 ;
      RECT 186.445 12.495 186.615 12.665 ;
      RECT 186.445 15.215 186.615 15.385 ;
      RECT 186.445 17.935 186.615 18.105 ;
      RECT 186.445 20.655 186.615 20.825 ;
      RECT 186.445 23.375 186.615 23.545 ;
      RECT 186.445 26.095 186.615 26.265 ;
      RECT 186.445 28.815 186.615 28.985 ;
      RECT 186.445 31.535 186.615 31.705 ;
      RECT 186.445 34.255 186.615 34.425 ;
      RECT 186.445 36.975 186.615 37.145 ;
      RECT 186.445 39.695 186.615 39.865 ;
      RECT 186.445 42.415 186.615 42.585 ;
      RECT 186.445 45.135 186.615 45.305 ;
      RECT 186.445 47.855 186.615 48.025 ;
      RECT 186.445 50.575 186.615 50.745 ;
      RECT 186.445 53.295 186.615 53.465 ;
      RECT 186.445 56.015 186.615 56.185 ;
      RECT 186.445 58.735 186.615 58.905 ;
      RECT 185.985 9.775 186.155 9.945 ;
      RECT 185.985 12.495 186.155 12.665 ;
      RECT 185.985 15.215 186.155 15.385 ;
      RECT 185.985 17.935 186.155 18.105 ;
      RECT 185.985 20.655 186.155 20.825 ;
      RECT 185.985 23.375 186.155 23.545 ;
      RECT 185.985 26.095 186.155 26.265 ;
      RECT 185.985 28.815 186.155 28.985 ;
      RECT 185.985 31.535 186.155 31.705 ;
      RECT 185.985 34.255 186.155 34.425 ;
      RECT 185.985 36.975 186.155 37.145 ;
      RECT 185.985 39.695 186.155 39.865 ;
      RECT 185.985 42.415 186.155 42.585 ;
      RECT 185.985 45.135 186.155 45.305 ;
      RECT 185.985 47.855 186.155 48.025 ;
      RECT 185.985 50.575 186.155 50.745 ;
      RECT 185.985 53.295 186.155 53.465 ;
      RECT 185.985 56.015 186.155 56.185 ;
      RECT 185.985 58.735 186.155 58.905 ;
      RECT 185.525 9.775 185.695 9.945 ;
      RECT 185.525 12.495 185.695 12.665 ;
      RECT 185.525 15.215 185.695 15.385 ;
      RECT 185.525 17.935 185.695 18.105 ;
      RECT 185.525 20.655 185.695 20.825 ;
      RECT 185.525 23.375 185.695 23.545 ;
      RECT 185.525 26.095 185.695 26.265 ;
      RECT 185.525 28.815 185.695 28.985 ;
      RECT 185.525 31.535 185.695 31.705 ;
      RECT 185.525 34.255 185.695 34.425 ;
      RECT 185.525 36.975 185.695 37.145 ;
      RECT 185.525 39.695 185.695 39.865 ;
      RECT 185.525 42.415 185.695 42.585 ;
      RECT 185.525 45.135 185.695 45.305 ;
      RECT 185.525 47.855 185.695 48.025 ;
      RECT 185.525 50.575 185.695 50.745 ;
      RECT 185.525 53.295 185.695 53.465 ;
      RECT 185.525 56.015 185.695 56.185 ;
      RECT 185.525 58.735 185.695 58.905 ;
      RECT 185.065 9.775 185.235 9.945 ;
      RECT 185.065 12.495 185.235 12.665 ;
      RECT 185.065 15.215 185.235 15.385 ;
      RECT 185.065 17.935 185.235 18.105 ;
      RECT 185.065 20.655 185.235 20.825 ;
      RECT 185.065 23.375 185.235 23.545 ;
      RECT 185.065 26.095 185.235 26.265 ;
      RECT 185.065 28.815 185.235 28.985 ;
      RECT 185.065 31.535 185.235 31.705 ;
      RECT 185.065 34.255 185.235 34.425 ;
      RECT 185.065 36.975 185.235 37.145 ;
      RECT 185.065 39.695 185.235 39.865 ;
      RECT 185.065 42.415 185.235 42.585 ;
      RECT 185.065 45.135 185.235 45.305 ;
      RECT 185.065 47.855 185.235 48.025 ;
      RECT 185.065 50.575 185.235 50.745 ;
      RECT 185.065 53.295 185.235 53.465 ;
      RECT 185.065 56.015 185.235 56.185 ;
      RECT 185.065 58.735 185.235 58.905 ;
      RECT 184.605 9.775 184.775 9.945 ;
      RECT 184.605 12.495 184.775 12.665 ;
      RECT 184.605 15.215 184.775 15.385 ;
      RECT 184.605 17.935 184.775 18.105 ;
      RECT 184.605 20.655 184.775 20.825 ;
      RECT 184.605 23.375 184.775 23.545 ;
      RECT 184.605 26.095 184.775 26.265 ;
      RECT 184.605 28.815 184.775 28.985 ;
      RECT 184.605 31.535 184.775 31.705 ;
      RECT 184.605 34.255 184.775 34.425 ;
      RECT 184.605 36.975 184.775 37.145 ;
      RECT 184.605 39.695 184.775 39.865 ;
      RECT 184.605 42.415 184.775 42.585 ;
      RECT 184.605 45.135 184.775 45.305 ;
      RECT 184.605 47.855 184.775 48.025 ;
      RECT 184.605 50.575 184.775 50.745 ;
      RECT 184.605 53.295 184.775 53.465 ;
      RECT 184.605 56.015 184.775 56.185 ;
      RECT 184.605 58.735 184.775 58.905 ;
      RECT 184.145 9.775 184.315 9.945 ;
      RECT 184.145 12.495 184.315 12.665 ;
      RECT 184.145 15.215 184.315 15.385 ;
      RECT 184.145 15.725 184.315 15.895 ;
      RECT 184.145 17.935 184.315 18.105 ;
      RECT 184.145 20.655 184.315 20.825 ;
      RECT 184.145 23.375 184.315 23.545 ;
      RECT 184.145 26.095 184.315 26.265 ;
      RECT 184.145 28.815 184.315 28.985 ;
      RECT 184.145 31.535 184.315 31.705 ;
      RECT 184.145 34.255 184.315 34.425 ;
      RECT 184.145 36.975 184.315 37.145 ;
      RECT 184.145 39.695 184.315 39.865 ;
      RECT 184.145 42.415 184.315 42.585 ;
      RECT 184.145 45.135 184.315 45.305 ;
      RECT 184.145 47.855 184.315 48.025 ;
      RECT 184.145 50.575 184.315 50.745 ;
      RECT 184.145 53.295 184.315 53.465 ;
      RECT 184.145 56.015 184.315 56.185 ;
      RECT 184.145 58.735 184.315 58.905 ;
      RECT 183.685 9.775 183.855 9.945 ;
      RECT 183.685 11.985 183.855 12.155 ;
      RECT 183.685 12.495 183.855 12.665 ;
      RECT 183.685 15.215 183.855 15.385 ;
      RECT 183.685 17.935 183.855 18.105 ;
      RECT 183.685 20.655 183.855 20.825 ;
      RECT 183.685 23.375 183.855 23.545 ;
      RECT 183.685 26.095 183.855 26.265 ;
      RECT 183.685 28.815 183.855 28.985 ;
      RECT 183.685 31.535 183.855 31.705 ;
      RECT 183.685 34.255 183.855 34.425 ;
      RECT 183.685 36.975 183.855 37.145 ;
      RECT 183.685 39.695 183.855 39.865 ;
      RECT 183.685 42.415 183.855 42.585 ;
      RECT 183.685 45.135 183.855 45.305 ;
      RECT 183.685 47.855 183.855 48.025 ;
      RECT 183.685 50.575 183.855 50.745 ;
      RECT 183.685 53.295 183.855 53.465 ;
      RECT 183.685 56.015 183.855 56.185 ;
      RECT 183.685 58.735 183.855 58.905 ;
      RECT 183.225 9.775 183.395 9.945 ;
      RECT 183.225 12.495 183.395 12.665 ;
      RECT 183.225 15.215 183.395 15.385 ;
      RECT 183.225 17.935 183.395 18.105 ;
      RECT 183.225 20.655 183.395 20.825 ;
      RECT 183.225 23.375 183.395 23.545 ;
      RECT 183.225 26.095 183.395 26.265 ;
      RECT 183.225 28.815 183.395 28.985 ;
      RECT 183.225 31.535 183.395 31.705 ;
      RECT 183.225 34.255 183.395 34.425 ;
      RECT 183.225 36.975 183.395 37.145 ;
      RECT 183.225 39.695 183.395 39.865 ;
      RECT 183.225 42.415 183.395 42.585 ;
      RECT 183.225 45.135 183.395 45.305 ;
      RECT 183.225 47.855 183.395 48.025 ;
      RECT 183.225 50.575 183.395 50.745 ;
      RECT 183.225 53.295 183.395 53.465 ;
      RECT 183.225 56.015 183.395 56.185 ;
      RECT 183.225 58.735 183.395 58.905 ;
      RECT 182.765 9.775 182.935 9.945 ;
      RECT 182.765 12.495 182.935 12.665 ;
      RECT 182.765 15.215 182.935 15.385 ;
      RECT 182.765 17.935 182.935 18.105 ;
      RECT 182.765 20.655 182.935 20.825 ;
      RECT 182.765 23.375 182.935 23.545 ;
      RECT 182.765 26.095 182.935 26.265 ;
      RECT 182.765 28.815 182.935 28.985 ;
      RECT 182.765 31.535 182.935 31.705 ;
      RECT 182.765 34.255 182.935 34.425 ;
      RECT 182.765 36.975 182.935 37.145 ;
      RECT 182.765 39.695 182.935 39.865 ;
      RECT 182.765 42.415 182.935 42.585 ;
      RECT 182.765 45.135 182.935 45.305 ;
      RECT 182.765 47.855 182.935 48.025 ;
      RECT 182.765 50.575 182.935 50.745 ;
      RECT 182.765 53.295 182.935 53.465 ;
      RECT 182.765 56.015 182.935 56.185 ;
      RECT 182.765 58.735 182.935 58.905 ;
      RECT 182.305 9.775 182.475 9.945 ;
      RECT 182.305 12.495 182.475 12.665 ;
      RECT 182.305 15.215 182.475 15.385 ;
      RECT 182.305 17.935 182.475 18.105 ;
      RECT 182.305 20.655 182.475 20.825 ;
      RECT 182.305 23.375 182.475 23.545 ;
      RECT 182.305 26.095 182.475 26.265 ;
      RECT 182.305 28.815 182.475 28.985 ;
      RECT 182.305 31.535 182.475 31.705 ;
      RECT 182.305 34.255 182.475 34.425 ;
      RECT 182.305 36.975 182.475 37.145 ;
      RECT 182.305 39.695 182.475 39.865 ;
      RECT 182.305 42.415 182.475 42.585 ;
      RECT 182.305 45.135 182.475 45.305 ;
      RECT 182.305 47.855 182.475 48.025 ;
      RECT 182.305 50.575 182.475 50.745 ;
      RECT 182.305 53.295 182.475 53.465 ;
      RECT 182.305 56.015 182.475 56.185 ;
      RECT 182.305 58.735 182.475 58.905 ;
      RECT 181.845 9.775 182.015 9.945 ;
      RECT 181.845 12.495 182.015 12.665 ;
      RECT 181.845 15.215 182.015 15.385 ;
      RECT 181.845 17.935 182.015 18.105 ;
      RECT 181.845 20.655 182.015 20.825 ;
      RECT 181.845 23.375 182.015 23.545 ;
      RECT 181.845 26.095 182.015 26.265 ;
      RECT 181.845 28.815 182.015 28.985 ;
      RECT 181.845 31.535 182.015 31.705 ;
      RECT 181.845 34.255 182.015 34.425 ;
      RECT 181.845 36.975 182.015 37.145 ;
      RECT 181.845 39.695 182.015 39.865 ;
      RECT 181.845 42.415 182.015 42.585 ;
      RECT 181.845 45.135 182.015 45.305 ;
      RECT 181.845 47.855 182.015 48.025 ;
      RECT 181.845 50.575 182.015 50.745 ;
      RECT 181.845 53.295 182.015 53.465 ;
      RECT 181.845 56.015 182.015 56.185 ;
      RECT 181.845 58.735 182.015 58.905 ;
      RECT 181.835 16.405 182.005 16.575 ;
      RECT 181.4 16.065 181.57 16.235 ;
      RECT 181.385 9.775 181.555 9.945 ;
      RECT 181.385 12.495 181.555 12.665 ;
      RECT 181.385 15.215 181.555 15.385 ;
      RECT 181.385 17.935 181.555 18.105 ;
      RECT 181.385 20.655 181.555 20.825 ;
      RECT 181.385 23.375 181.555 23.545 ;
      RECT 181.385 26.095 181.555 26.265 ;
      RECT 181.385 28.815 181.555 28.985 ;
      RECT 181.385 31.535 181.555 31.705 ;
      RECT 181.385 34.255 181.555 34.425 ;
      RECT 181.385 36.975 181.555 37.145 ;
      RECT 181.385 39.695 181.555 39.865 ;
      RECT 181.385 42.415 181.555 42.585 ;
      RECT 181.385 45.135 181.555 45.305 ;
      RECT 181.385 47.855 181.555 48.025 ;
      RECT 181.385 50.575 181.555 50.745 ;
      RECT 181.385 53.295 181.555 53.465 ;
      RECT 181.385 56.015 181.555 56.185 ;
      RECT 181.385 58.735 181.555 58.905 ;
      RECT 180.925 9.775 181.095 9.945 ;
      RECT 180.925 12.495 181.095 12.665 ;
      RECT 180.925 15.215 181.095 15.385 ;
      RECT 180.925 17.935 181.095 18.105 ;
      RECT 180.925 20.655 181.095 20.825 ;
      RECT 180.925 23.375 181.095 23.545 ;
      RECT 180.925 26.095 181.095 26.265 ;
      RECT 180.925 28.815 181.095 28.985 ;
      RECT 180.925 31.535 181.095 31.705 ;
      RECT 180.925 34.255 181.095 34.425 ;
      RECT 180.925 36.975 181.095 37.145 ;
      RECT 180.925 39.695 181.095 39.865 ;
      RECT 180.925 42.415 181.095 42.585 ;
      RECT 180.925 45.135 181.095 45.305 ;
      RECT 180.925 47.855 181.095 48.025 ;
      RECT 180.925 50.575 181.095 50.745 ;
      RECT 180.925 53.295 181.095 53.465 ;
      RECT 180.925 56.015 181.095 56.185 ;
      RECT 180.925 58.735 181.095 58.905 ;
      RECT 180.465 9.775 180.635 9.945 ;
      RECT 180.465 12.495 180.635 12.665 ;
      RECT 180.465 15.215 180.635 15.385 ;
      RECT 180.465 17.935 180.635 18.105 ;
      RECT 180.465 20.655 180.635 20.825 ;
      RECT 180.465 23.375 180.635 23.545 ;
      RECT 180.465 26.095 180.635 26.265 ;
      RECT 180.465 28.815 180.635 28.985 ;
      RECT 180.465 31.535 180.635 31.705 ;
      RECT 180.465 34.255 180.635 34.425 ;
      RECT 180.465 36.975 180.635 37.145 ;
      RECT 180.465 39.695 180.635 39.865 ;
      RECT 180.465 42.415 180.635 42.585 ;
      RECT 180.465 45.135 180.635 45.305 ;
      RECT 180.465 47.855 180.635 48.025 ;
      RECT 180.465 50.575 180.635 50.745 ;
      RECT 180.465 53.295 180.635 53.465 ;
      RECT 180.465 56.015 180.635 56.185 ;
      RECT 180.465 58.735 180.635 58.905 ;
      RECT 180.005 9.775 180.175 9.945 ;
      RECT 180.005 12.495 180.175 12.665 ;
      RECT 180.005 15.215 180.175 15.385 ;
      RECT 180.005 17.935 180.175 18.105 ;
      RECT 180.005 20.655 180.175 20.825 ;
      RECT 180.005 23.375 180.175 23.545 ;
      RECT 180.005 26.095 180.175 26.265 ;
      RECT 180.005 28.815 180.175 28.985 ;
      RECT 180.005 31.535 180.175 31.705 ;
      RECT 180.005 34.255 180.175 34.425 ;
      RECT 180.005 36.975 180.175 37.145 ;
      RECT 180.005 39.695 180.175 39.865 ;
      RECT 180.005 42.415 180.175 42.585 ;
      RECT 180.005 45.135 180.175 45.305 ;
      RECT 180.005 47.855 180.175 48.025 ;
      RECT 180.005 50.575 180.175 50.745 ;
      RECT 180.005 53.295 180.175 53.465 ;
      RECT 180.005 56.015 180.175 56.185 ;
      RECT 180.005 58.735 180.175 58.905 ;
      RECT 179.83 16.065 180 16.235 ;
      RECT 179.545 9.775 179.715 9.945 ;
      RECT 179.545 12.495 179.715 12.665 ;
      RECT 179.545 15.215 179.715 15.385 ;
      RECT 179.545 17.935 179.715 18.105 ;
      RECT 179.545 20.655 179.715 20.825 ;
      RECT 179.545 23.375 179.715 23.545 ;
      RECT 179.545 26.095 179.715 26.265 ;
      RECT 179.545 28.815 179.715 28.985 ;
      RECT 179.545 31.535 179.715 31.705 ;
      RECT 179.545 34.255 179.715 34.425 ;
      RECT 179.545 36.975 179.715 37.145 ;
      RECT 179.545 39.695 179.715 39.865 ;
      RECT 179.545 42.415 179.715 42.585 ;
      RECT 179.545 45.135 179.715 45.305 ;
      RECT 179.545 47.855 179.715 48.025 ;
      RECT 179.545 50.575 179.715 50.745 ;
      RECT 179.545 53.295 179.715 53.465 ;
      RECT 179.545 56.015 179.715 56.185 ;
      RECT 179.545 58.735 179.715 58.905 ;
      RECT 179.315 16.405 179.485 16.575 ;
      RECT 179.085 9.775 179.255 9.945 ;
      RECT 179.085 12.495 179.255 12.665 ;
      RECT 179.085 15.215 179.255 15.385 ;
      RECT 179.085 17.935 179.255 18.105 ;
      RECT 179.085 20.655 179.255 20.825 ;
      RECT 179.085 23.375 179.255 23.545 ;
      RECT 179.085 26.095 179.255 26.265 ;
      RECT 179.085 28.815 179.255 28.985 ;
      RECT 179.085 31.535 179.255 31.705 ;
      RECT 179.085 34.255 179.255 34.425 ;
      RECT 179.085 36.975 179.255 37.145 ;
      RECT 179.085 39.695 179.255 39.865 ;
      RECT 179.085 42.415 179.255 42.585 ;
      RECT 179.085 45.135 179.255 45.305 ;
      RECT 179.085 47.855 179.255 48.025 ;
      RECT 179.085 50.575 179.255 50.745 ;
      RECT 179.085 53.295 179.255 53.465 ;
      RECT 179.085 56.015 179.255 56.185 ;
      RECT 179.085 58.735 179.255 58.905 ;
      RECT 178.625 9.775 178.795 9.945 ;
      RECT 178.625 12.495 178.795 12.665 ;
      RECT 178.625 15.215 178.795 15.385 ;
      RECT 178.625 17.935 178.795 18.105 ;
      RECT 178.625 20.655 178.795 20.825 ;
      RECT 178.625 23.375 178.795 23.545 ;
      RECT 178.625 26.095 178.795 26.265 ;
      RECT 178.625 28.815 178.795 28.985 ;
      RECT 178.625 31.535 178.795 31.705 ;
      RECT 178.625 34.255 178.795 34.425 ;
      RECT 178.625 36.975 178.795 37.145 ;
      RECT 178.625 39.695 178.795 39.865 ;
      RECT 178.625 42.415 178.795 42.585 ;
      RECT 178.625 45.135 178.795 45.305 ;
      RECT 178.625 47.855 178.795 48.025 ;
      RECT 178.625 50.575 178.795 50.745 ;
      RECT 178.625 53.295 178.795 53.465 ;
      RECT 178.625 56.015 178.795 56.185 ;
      RECT 178.625 58.735 178.795 58.905 ;
      RECT 178.55 17.085 178.72 17.255 ;
      RECT 178.165 9.775 178.335 9.945 ;
      RECT 178.165 12.495 178.335 12.665 ;
      RECT 178.165 15.215 178.335 15.385 ;
      RECT 178.165 17.935 178.335 18.105 ;
      RECT 178.165 20.655 178.335 20.825 ;
      RECT 178.165 23.375 178.335 23.545 ;
      RECT 178.165 26.095 178.335 26.265 ;
      RECT 178.165 28.815 178.335 28.985 ;
      RECT 178.165 31.535 178.335 31.705 ;
      RECT 178.165 34.255 178.335 34.425 ;
      RECT 178.165 36.975 178.335 37.145 ;
      RECT 178.165 39.695 178.335 39.865 ;
      RECT 178.165 42.415 178.335 42.585 ;
      RECT 178.165 45.135 178.335 45.305 ;
      RECT 178.165 47.855 178.335 48.025 ;
      RECT 178.165 50.575 178.335 50.745 ;
      RECT 178.165 53.295 178.335 53.465 ;
      RECT 178.165 56.015 178.335 56.185 ;
      RECT 178.165 58.735 178.335 58.905 ;
      RECT 178.125 16.405 178.295 16.575 ;
      RECT 177.73 16.065 177.9 16.235 ;
      RECT 177.705 9.775 177.875 9.945 ;
      RECT 177.705 12.495 177.875 12.665 ;
      RECT 177.705 15.215 177.875 15.385 ;
      RECT 177.705 17.935 177.875 18.105 ;
      RECT 177.705 20.655 177.875 20.825 ;
      RECT 177.705 23.375 177.875 23.545 ;
      RECT 177.705 26.095 177.875 26.265 ;
      RECT 177.705 28.815 177.875 28.985 ;
      RECT 177.705 31.535 177.875 31.705 ;
      RECT 177.705 34.255 177.875 34.425 ;
      RECT 177.705 36.975 177.875 37.145 ;
      RECT 177.705 39.695 177.875 39.865 ;
      RECT 177.705 42.415 177.875 42.585 ;
      RECT 177.705 45.135 177.875 45.305 ;
      RECT 177.705 47.855 177.875 48.025 ;
      RECT 177.705 50.575 177.875 50.745 ;
      RECT 177.705 53.295 177.875 53.465 ;
      RECT 177.705 56.015 177.875 56.185 ;
      RECT 177.705 58.735 177.875 58.905 ;
      RECT 177.245 9.775 177.415 9.945 ;
      RECT 177.245 11.305 177.415 11.475 ;
      RECT 177.245 12.495 177.415 12.665 ;
      RECT 177.245 15.215 177.415 15.385 ;
      RECT 177.245 16.745 177.415 16.915 ;
      RECT 177.245 17.935 177.415 18.105 ;
      RECT 177.245 20.655 177.415 20.825 ;
      RECT 177.245 23.375 177.415 23.545 ;
      RECT 177.245 26.095 177.415 26.265 ;
      RECT 177.245 28.815 177.415 28.985 ;
      RECT 177.245 31.535 177.415 31.705 ;
      RECT 177.245 34.255 177.415 34.425 ;
      RECT 177.245 36.975 177.415 37.145 ;
      RECT 177.245 39.695 177.415 39.865 ;
      RECT 177.245 42.415 177.415 42.585 ;
      RECT 177.245 45.135 177.415 45.305 ;
      RECT 177.245 47.855 177.415 48.025 ;
      RECT 177.245 50.575 177.415 50.745 ;
      RECT 177.245 53.295 177.415 53.465 ;
      RECT 177.245 56.015 177.415 56.185 ;
      RECT 177.245 58.735 177.415 58.905 ;
      RECT 176.785 9.775 176.955 9.945 ;
      RECT 176.785 12.495 176.955 12.665 ;
      RECT 176.785 15.215 176.955 15.385 ;
      RECT 176.785 17.935 176.955 18.105 ;
      RECT 176.785 20.655 176.955 20.825 ;
      RECT 176.785 23.375 176.955 23.545 ;
      RECT 176.785 26.095 176.955 26.265 ;
      RECT 176.785 28.815 176.955 28.985 ;
      RECT 176.785 31.535 176.955 31.705 ;
      RECT 176.785 34.255 176.955 34.425 ;
      RECT 176.785 36.975 176.955 37.145 ;
      RECT 176.785 39.695 176.955 39.865 ;
      RECT 176.785 42.415 176.955 42.585 ;
      RECT 176.785 45.135 176.955 45.305 ;
      RECT 176.785 47.855 176.955 48.025 ;
      RECT 176.785 50.575 176.955 50.745 ;
      RECT 176.785 53.295 176.955 53.465 ;
      RECT 176.785 56.015 176.955 56.185 ;
      RECT 176.785 58.735 176.955 58.905 ;
      RECT 176.325 9.775 176.495 9.945 ;
      RECT 176.325 12.495 176.495 12.665 ;
      RECT 176.325 15.215 176.495 15.385 ;
      RECT 176.325 17.935 176.495 18.105 ;
      RECT 176.325 20.655 176.495 20.825 ;
      RECT 176.325 23.375 176.495 23.545 ;
      RECT 176.325 26.095 176.495 26.265 ;
      RECT 176.325 28.815 176.495 28.985 ;
      RECT 176.325 31.535 176.495 31.705 ;
      RECT 176.325 34.255 176.495 34.425 ;
      RECT 176.325 36.975 176.495 37.145 ;
      RECT 176.325 39.695 176.495 39.865 ;
      RECT 176.325 42.415 176.495 42.585 ;
      RECT 176.325 45.135 176.495 45.305 ;
      RECT 176.325 47.855 176.495 48.025 ;
      RECT 176.325 50.575 176.495 50.745 ;
      RECT 176.325 53.295 176.495 53.465 ;
      RECT 176.325 56.015 176.495 56.185 ;
      RECT 176.325 58.735 176.495 58.905 ;
      RECT 175.865 9.775 176.035 9.945 ;
      RECT 175.865 12.495 176.035 12.665 ;
      RECT 175.865 15.215 176.035 15.385 ;
      RECT 175.865 17.935 176.035 18.105 ;
      RECT 175.865 20.655 176.035 20.825 ;
      RECT 175.865 23.375 176.035 23.545 ;
      RECT 175.865 26.095 176.035 26.265 ;
      RECT 175.865 28.815 176.035 28.985 ;
      RECT 175.865 31.535 176.035 31.705 ;
      RECT 175.865 34.255 176.035 34.425 ;
      RECT 175.865 36.975 176.035 37.145 ;
      RECT 175.865 39.695 176.035 39.865 ;
      RECT 175.865 42.415 176.035 42.585 ;
      RECT 175.865 45.135 176.035 45.305 ;
      RECT 175.865 47.855 176.035 48.025 ;
      RECT 175.865 50.575 176.035 50.745 ;
      RECT 175.865 53.295 176.035 53.465 ;
      RECT 175.865 56.015 176.035 56.185 ;
      RECT 175.865 58.735 176.035 58.905 ;
      RECT 175.405 9.775 175.575 9.945 ;
      RECT 175.405 12.495 175.575 12.665 ;
      RECT 175.405 15.215 175.575 15.385 ;
      RECT 175.405 17.935 175.575 18.105 ;
      RECT 175.405 20.655 175.575 20.825 ;
      RECT 175.405 23.375 175.575 23.545 ;
      RECT 175.405 26.095 175.575 26.265 ;
      RECT 175.405 28.815 175.575 28.985 ;
      RECT 175.405 31.535 175.575 31.705 ;
      RECT 175.405 34.255 175.575 34.425 ;
      RECT 175.405 36.975 175.575 37.145 ;
      RECT 175.405 39.695 175.575 39.865 ;
      RECT 175.405 42.415 175.575 42.585 ;
      RECT 175.405 45.135 175.575 45.305 ;
      RECT 175.405 47.855 175.575 48.025 ;
      RECT 175.405 50.575 175.575 50.745 ;
      RECT 175.405 53.295 175.575 53.465 ;
      RECT 175.405 56.015 175.575 56.185 ;
      RECT 175.405 58.735 175.575 58.905 ;
      RECT 174.945 9.775 175.115 9.945 ;
      RECT 174.945 12.495 175.115 12.665 ;
      RECT 174.945 15.215 175.115 15.385 ;
      RECT 174.945 17.935 175.115 18.105 ;
      RECT 174.945 20.655 175.115 20.825 ;
      RECT 174.945 23.375 175.115 23.545 ;
      RECT 174.945 26.095 175.115 26.265 ;
      RECT 174.945 28.815 175.115 28.985 ;
      RECT 174.945 31.535 175.115 31.705 ;
      RECT 174.945 34.255 175.115 34.425 ;
      RECT 174.945 36.975 175.115 37.145 ;
      RECT 174.945 39.695 175.115 39.865 ;
      RECT 174.945 42.415 175.115 42.585 ;
      RECT 174.945 45.135 175.115 45.305 ;
      RECT 174.945 47.855 175.115 48.025 ;
      RECT 174.945 50.575 175.115 50.745 ;
      RECT 174.945 53.295 175.115 53.465 ;
      RECT 174.945 56.015 175.115 56.185 ;
      RECT 174.945 58.735 175.115 58.905 ;
      RECT 174.485 9.775 174.655 9.945 ;
      RECT 174.485 12.495 174.655 12.665 ;
      RECT 174.485 15.215 174.655 15.385 ;
      RECT 174.485 17.935 174.655 18.105 ;
      RECT 174.485 19.805 174.655 19.975 ;
      RECT 174.485 20.655 174.655 20.825 ;
      RECT 174.485 23.375 174.655 23.545 ;
      RECT 174.485 26.095 174.655 26.265 ;
      RECT 174.485 28.815 174.655 28.985 ;
      RECT 174.485 31.535 174.655 31.705 ;
      RECT 174.485 34.255 174.655 34.425 ;
      RECT 174.485 36.975 174.655 37.145 ;
      RECT 174.485 39.695 174.655 39.865 ;
      RECT 174.485 42.415 174.655 42.585 ;
      RECT 174.485 45.135 174.655 45.305 ;
      RECT 174.485 47.855 174.655 48.025 ;
      RECT 174.485 50.575 174.655 50.745 ;
      RECT 174.485 53.295 174.655 53.465 ;
      RECT 174.485 56.015 174.655 56.185 ;
      RECT 174.485 58.735 174.655 58.905 ;
      RECT 174.025 9.775 174.195 9.945 ;
      RECT 174.025 12.495 174.195 12.665 ;
      RECT 174.025 15.215 174.195 15.385 ;
      RECT 174.025 17.935 174.195 18.105 ;
      RECT 174.025 20.655 174.195 20.825 ;
      RECT 174.025 23.375 174.195 23.545 ;
      RECT 174.025 26.095 174.195 26.265 ;
      RECT 174.025 28.815 174.195 28.985 ;
      RECT 174.025 31.535 174.195 31.705 ;
      RECT 174.025 34.255 174.195 34.425 ;
      RECT 174.025 36.975 174.195 37.145 ;
      RECT 174.025 39.695 174.195 39.865 ;
      RECT 174.025 42.415 174.195 42.585 ;
      RECT 174.025 45.135 174.195 45.305 ;
      RECT 174.025 47.855 174.195 48.025 ;
      RECT 174.025 50.575 174.195 50.745 ;
      RECT 174.025 53.295 174.195 53.465 ;
      RECT 174.025 56.015 174.195 56.185 ;
      RECT 174.025 58.735 174.195 58.905 ;
      RECT 173.565 9.775 173.735 9.945 ;
      RECT 173.565 12.495 173.735 12.665 ;
      RECT 173.565 15.215 173.735 15.385 ;
      RECT 173.565 17.935 173.735 18.105 ;
      RECT 173.565 20.655 173.735 20.825 ;
      RECT 173.565 23.375 173.735 23.545 ;
      RECT 173.565 26.095 173.735 26.265 ;
      RECT 173.565 28.815 173.735 28.985 ;
      RECT 173.565 31.535 173.735 31.705 ;
      RECT 173.565 34.255 173.735 34.425 ;
      RECT 173.565 36.975 173.735 37.145 ;
      RECT 173.565 39.695 173.735 39.865 ;
      RECT 173.565 42.415 173.735 42.585 ;
      RECT 173.565 45.135 173.735 45.305 ;
      RECT 173.565 47.855 173.735 48.025 ;
      RECT 173.565 50.575 173.735 50.745 ;
      RECT 173.565 53.295 173.735 53.465 ;
      RECT 173.565 56.015 173.735 56.185 ;
      RECT 173.565 58.735 173.735 58.905 ;
      RECT 173.105 9.775 173.275 9.945 ;
      RECT 173.105 12.495 173.275 12.665 ;
      RECT 173.105 15.215 173.275 15.385 ;
      RECT 173.105 17.425 173.275 17.595 ;
      RECT 173.105 17.935 173.275 18.105 ;
      RECT 173.105 20.655 173.275 20.825 ;
      RECT 173.105 23.375 173.275 23.545 ;
      RECT 173.105 26.095 173.275 26.265 ;
      RECT 173.105 28.815 173.275 28.985 ;
      RECT 173.105 31.535 173.275 31.705 ;
      RECT 173.105 34.255 173.275 34.425 ;
      RECT 173.105 36.975 173.275 37.145 ;
      RECT 173.105 39.695 173.275 39.865 ;
      RECT 173.105 42.415 173.275 42.585 ;
      RECT 173.105 45.135 173.275 45.305 ;
      RECT 173.105 47.855 173.275 48.025 ;
      RECT 173.105 50.575 173.275 50.745 ;
      RECT 173.105 53.295 173.275 53.465 ;
      RECT 173.105 56.015 173.275 56.185 ;
      RECT 173.105 58.735 173.275 58.905 ;
      RECT 172.645 9.775 172.815 9.945 ;
      RECT 172.645 12.495 172.815 12.665 ;
      RECT 172.645 15.215 172.815 15.385 ;
      RECT 172.645 17.935 172.815 18.105 ;
      RECT 172.645 20.655 172.815 20.825 ;
      RECT 172.645 23.375 172.815 23.545 ;
      RECT 172.645 26.095 172.815 26.265 ;
      RECT 172.645 28.815 172.815 28.985 ;
      RECT 172.645 31.535 172.815 31.705 ;
      RECT 172.645 34.255 172.815 34.425 ;
      RECT 172.645 36.975 172.815 37.145 ;
      RECT 172.645 39.695 172.815 39.865 ;
      RECT 172.645 42.415 172.815 42.585 ;
      RECT 172.645 45.135 172.815 45.305 ;
      RECT 172.645 47.855 172.815 48.025 ;
      RECT 172.645 50.575 172.815 50.745 ;
      RECT 172.645 53.295 172.815 53.465 ;
      RECT 172.645 56.015 172.815 56.185 ;
      RECT 172.645 58.735 172.815 58.905 ;
      RECT 172.185 9.775 172.355 9.945 ;
      RECT 172.185 12.495 172.355 12.665 ;
      RECT 172.185 15.215 172.355 15.385 ;
      RECT 172.185 17.935 172.355 18.105 ;
      RECT 172.185 20.655 172.355 20.825 ;
      RECT 172.185 23.375 172.355 23.545 ;
      RECT 172.185 26.095 172.355 26.265 ;
      RECT 172.185 28.815 172.355 28.985 ;
      RECT 172.185 31.535 172.355 31.705 ;
      RECT 172.185 34.255 172.355 34.425 ;
      RECT 172.185 36.975 172.355 37.145 ;
      RECT 172.185 39.695 172.355 39.865 ;
      RECT 172.185 42.415 172.355 42.585 ;
      RECT 172.185 45.135 172.355 45.305 ;
      RECT 172.185 47.855 172.355 48.025 ;
      RECT 172.185 50.575 172.355 50.745 ;
      RECT 172.185 53.295 172.355 53.465 ;
      RECT 172.185 56.015 172.355 56.185 ;
      RECT 172.185 58.735 172.355 58.905 ;
      RECT 171.725 9.775 171.895 9.945 ;
      RECT 171.725 12.495 171.895 12.665 ;
      RECT 171.725 14.705 171.895 14.875 ;
      RECT 171.725 15.215 171.895 15.385 ;
      RECT 171.725 17.935 171.895 18.105 ;
      RECT 171.725 19.125 171.895 19.295 ;
      RECT 171.725 20.655 171.895 20.825 ;
      RECT 171.725 23.375 171.895 23.545 ;
      RECT 171.725 26.095 171.895 26.265 ;
      RECT 171.725 28.815 171.895 28.985 ;
      RECT 171.725 31.535 171.895 31.705 ;
      RECT 171.725 34.255 171.895 34.425 ;
      RECT 171.725 36.975 171.895 37.145 ;
      RECT 171.725 39.695 171.895 39.865 ;
      RECT 171.725 42.415 171.895 42.585 ;
      RECT 171.725 45.135 171.895 45.305 ;
      RECT 171.725 47.855 171.895 48.025 ;
      RECT 171.725 50.575 171.895 50.745 ;
      RECT 171.725 53.295 171.895 53.465 ;
      RECT 171.725 56.015 171.895 56.185 ;
      RECT 171.725 58.735 171.895 58.905 ;
      RECT 171.265 9.775 171.435 9.945 ;
      RECT 171.265 12.495 171.435 12.665 ;
      RECT 171.265 15.215 171.435 15.385 ;
      RECT 171.265 17.935 171.435 18.105 ;
      RECT 171.265 19.465 171.435 19.635 ;
      RECT 171.265 20.655 171.435 20.825 ;
      RECT 171.265 22.185 171.435 22.355 ;
      RECT 171.265 23.375 171.435 23.545 ;
      RECT 171.265 26.095 171.435 26.265 ;
      RECT 171.265 28.815 171.435 28.985 ;
      RECT 171.265 30.005 171.435 30.175 ;
      RECT 171.265 31.535 171.435 31.705 ;
      RECT 171.265 34.255 171.435 34.425 ;
      RECT 171.265 36.975 171.435 37.145 ;
      RECT 171.265 39.695 171.435 39.865 ;
      RECT 171.265 42.415 171.435 42.585 ;
      RECT 171.265 45.135 171.435 45.305 ;
      RECT 171.265 47.855 171.435 48.025 ;
      RECT 171.265 50.575 171.435 50.745 ;
      RECT 171.265 53.295 171.435 53.465 ;
      RECT 171.265 56.015 171.435 56.185 ;
      RECT 171.265 58.735 171.435 58.905 ;
      RECT 170.805 9.775 170.975 9.945 ;
      RECT 170.805 12.495 170.975 12.665 ;
      RECT 170.805 15.215 170.975 15.385 ;
      RECT 170.805 17.935 170.975 18.105 ;
      RECT 170.805 20.655 170.975 20.825 ;
      RECT 170.805 23.375 170.975 23.545 ;
      RECT 170.805 26.095 170.975 26.265 ;
      RECT 170.805 28.815 170.975 28.985 ;
      RECT 170.805 31.535 170.975 31.705 ;
      RECT 170.805 34.255 170.975 34.425 ;
      RECT 170.805 36.975 170.975 37.145 ;
      RECT 170.805 39.695 170.975 39.865 ;
      RECT 170.805 42.415 170.975 42.585 ;
      RECT 170.805 45.135 170.975 45.305 ;
      RECT 170.805 47.855 170.975 48.025 ;
      RECT 170.805 50.575 170.975 50.745 ;
      RECT 170.805 53.295 170.975 53.465 ;
      RECT 170.805 56.015 170.975 56.185 ;
      RECT 170.805 58.735 170.975 58.905 ;
      RECT 170.345 9.775 170.515 9.945 ;
      RECT 170.345 12.495 170.515 12.665 ;
      RECT 170.345 15.215 170.515 15.385 ;
      RECT 170.345 16.405 170.515 16.575 ;
      RECT 170.345 17.935 170.515 18.105 ;
      RECT 170.345 19.125 170.515 19.295 ;
      RECT 170.345 20.655 170.515 20.825 ;
      RECT 170.345 23.375 170.515 23.545 ;
      RECT 170.345 26.095 170.515 26.265 ;
      RECT 170.345 28.815 170.515 28.985 ;
      RECT 170.345 31.535 170.515 31.705 ;
      RECT 170.345 34.255 170.515 34.425 ;
      RECT 170.345 36.975 170.515 37.145 ;
      RECT 170.345 39.695 170.515 39.865 ;
      RECT 170.345 42.415 170.515 42.585 ;
      RECT 170.345 45.135 170.515 45.305 ;
      RECT 170.345 47.855 170.515 48.025 ;
      RECT 170.345 50.575 170.515 50.745 ;
      RECT 170.345 53.295 170.515 53.465 ;
      RECT 170.345 56.015 170.515 56.185 ;
      RECT 170.345 58.735 170.515 58.905 ;
      RECT 169.885 9.775 170.055 9.945 ;
      RECT 169.885 12.495 170.055 12.665 ;
      RECT 169.885 15.215 170.055 15.385 ;
      RECT 169.885 17.935 170.055 18.105 ;
      RECT 169.885 20.655 170.055 20.825 ;
      RECT 169.885 23.375 170.055 23.545 ;
      RECT 169.885 26.095 170.055 26.265 ;
      RECT 169.885 28.815 170.055 28.985 ;
      RECT 169.885 31.535 170.055 31.705 ;
      RECT 169.885 34.255 170.055 34.425 ;
      RECT 169.885 36.975 170.055 37.145 ;
      RECT 169.885 39.695 170.055 39.865 ;
      RECT 169.885 42.415 170.055 42.585 ;
      RECT 169.885 45.135 170.055 45.305 ;
      RECT 169.885 47.855 170.055 48.025 ;
      RECT 169.885 50.575 170.055 50.745 ;
      RECT 169.885 53.295 170.055 53.465 ;
      RECT 169.885 56.015 170.055 56.185 ;
      RECT 169.885 58.735 170.055 58.905 ;
      RECT 169.425 9.775 169.595 9.945 ;
      RECT 169.425 12.495 169.595 12.665 ;
      RECT 169.425 15.215 169.595 15.385 ;
      RECT 169.425 15.725 169.595 15.895 ;
      RECT 169.425 17.935 169.595 18.105 ;
      RECT 169.425 18.445 169.595 18.615 ;
      RECT 169.425 20.655 169.595 20.825 ;
      RECT 169.425 23.375 169.595 23.545 ;
      RECT 169.425 26.095 169.595 26.265 ;
      RECT 169.425 28.815 169.595 28.985 ;
      RECT 169.425 31.535 169.595 31.705 ;
      RECT 169.425 34.255 169.595 34.425 ;
      RECT 169.425 36.975 169.595 37.145 ;
      RECT 169.425 39.695 169.595 39.865 ;
      RECT 169.425 42.415 169.595 42.585 ;
      RECT 169.425 45.135 169.595 45.305 ;
      RECT 169.425 47.855 169.595 48.025 ;
      RECT 169.425 50.575 169.595 50.745 ;
      RECT 169.425 53.295 169.595 53.465 ;
      RECT 169.425 56.015 169.595 56.185 ;
      RECT 169.425 58.735 169.595 58.905 ;
      RECT 168.965 9.775 169.135 9.945 ;
      RECT 168.965 11.305 169.135 11.475 ;
      RECT 168.965 12.495 169.135 12.665 ;
      RECT 168.965 15.215 169.135 15.385 ;
      RECT 168.965 17.935 169.135 18.105 ;
      RECT 168.965 19.125 169.135 19.295 ;
      RECT 168.965 20.655 169.135 20.825 ;
      RECT 168.965 23.375 169.135 23.545 ;
      RECT 168.965 26.095 169.135 26.265 ;
      RECT 168.965 28.815 169.135 28.985 ;
      RECT 168.965 31.535 169.135 31.705 ;
      RECT 168.965 34.255 169.135 34.425 ;
      RECT 168.965 36.975 169.135 37.145 ;
      RECT 168.965 39.695 169.135 39.865 ;
      RECT 168.965 42.415 169.135 42.585 ;
      RECT 168.965 45.135 169.135 45.305 ;
      RECT 168.965 47.855 169.135 48.025 ;
      RECT 168.965 50.575 169.135 50.745 ;
      RECT 168.965 53.295 169.135 53.465 ;
      RECT 168.965 56.015 169.135 56.185 ;
      RECT 168.965 58.735 169.135 58.905 ;
      RECT 168.505 9.775 168.675 9.945 ;
      RECT 168.505 12.495 168.675 12.665 ;
      RECT 168.505 15.215 168.675 15.385 ;
      RECT 168.505 17.935 168.675 18.105 ;
      RECT 168.505 20.655 168.675 20.825 ;
      RECT 168.505 23.375 168.675 23.545 ;
      RECT 168.505 26.095 168.675 26.265 ;
      RECT 168.505 28.815 168.675 28.985 ;
      RECT 168.505 31.535 168.675 31.705 ;
      RECT 168.505 34.255 168.675 34.425 ;
      RECT 168.505 36.975 168.675 37.145 ;
      RECT 168.505 39.695 168.675 39.865 ;
      RECT 168.505 42.415 168.675 42.585 ;
      RECT 168.505 45.135 168.675 45.305 ;
      RECT 168.505 47.855 168.675 48.025 ;
      RECT 168.505 50.575 168.675 50.745 ;
      RECT 168.505 53.295 168.675 53.465 ;
      RECT 168.505 56.015 168.675 56.185 ;
      RECT 168.505 58.735 168.675 58.905 ;
      RECT 168.045 9.775 168.215 9.945 ;
      RECT 168.045 12.495 168.215 12.665 ;
      RECT 168.045 15.215 168.215 15.385 ;
      RECT 168.045 17.935 168.215 18.105 ;
      RECT 168.045 20.655 168.215 20.825 ;
      RECT 168.045 23.375 168.215 23.545 ;
      RECT 168.045 26.095 168.215 26.265 ;
      RECT 168.045 28.815 168.215 28.985 ;
      RECT 168.045 31.535 168.215 31.705 ;
      RECT 168.045 34.255 168.215 34.425 ;
      RECT 168.045 36.975 168.215 37.145 ;
      RECT 168.045 39.695 168.215 39.865 ;
      RECT 168.045 42.415 168.215 42.585 ;
      RECT 168.045 45.135 168.215 45.305 ;
      RECT 168.045 47.855 168.215 48.025 ;
      RECT 168.045 50.575 168.215 50.745 ;
      RECT 168.045 53.295 168.215 53.465 ;
      RECT 168.045 56.015 168.215 56.185 ;
      RECT 168.045 58.735 168.215 58.905 ;
      RECT 167.585 9.775 167.755 9.945 ;
      RECT 167.585 12.495 167.755 12.665 ;
      RECT 167.585 15.215 167.755 15.385 ;
      RECT 167.585 17.935 167.755 18.105 ;
      RECT 167.585 20.655 167.755 20.825 ;
      RECT 167.585 23.375 167.755 23.545 ;
      RECT 167.585 26.095 167.755 26.265 ;
      RECT 167.585 28.815 167.755 28.985 ;
      RECT 167.585 31.535 167.755 31.705 ;
      RECT 167.585 34.255 167.755 34.425 ;
      RECT 167.585 36.975 167.755 37.145 ;
      RECT 167.585 39.695 167.755 39.865 ;
      RECT 167.585 42.415 167.755 42.585 ;
      RECT 167.585 45.135 167.755 45.305 ;
      RECT 167.585 47.855 167.755 48.025 ;
      RECT 167.585 50.575 167.755 50.745 ;
      RECT 167.585 53.295 167.755 53.465 ;
      RECT 167.585 56.015 167.755 56.185 ;
      RECT 167.585 58.735 167.755 58.905 ;
      RECT 167.125 9.775 167.295 9.945 ;
      RECT 167.125 12.495 167.295 12.665 ;
      RECT 167.125 15.215 167.295 15.385 ;
      RECT 167.125 17.935 167.295 18.105 ;
      RECT 167.125 20.655 167.295 20.825 ;
      RECT 167.125 23.375 167.295 23.545 ;
      RECT 167.125 26.095 167.295 26.265 ;
      RECT 167.125 28.815 167.295 28.985 ;
      RECT 167.125 31.535 167.295 31.705 ;
      RECT 167.125 34.255 167.295 34.425 ;
      RECT 167.125 36.975 167.295 37.145 ;
      RECT 167.125 39.695 167.295 39.865 ;
      RECT 167.125 42.415 167.295 42.585 ;
      RECT 167.125 45.135 167.295 45.305 ;
      RECT 167.125 47.855 167.295 48.025 ;
      RECT 167.125 50.575 167.295 50.745 ;
      RECT 167.125 53.295 167.295 53.465 ;
      RECT 167.125 56.015 167.295 56.185 ;
      RECT 167.125 58.735 167.295 58.905 ;
      RECT 167.115 16.405 167.285 16.575 ;
      RECT 166.68 16.065 166.85 16.235 ;
      RECT 166.665 9.775 166.835 9.945 ;
      RECT 166.665 12.495 166.835 12.665 ;
      RECT 166.665 15.215 166.835 15.385 ;
      RECT 166.665 17.935 166.835 18.105 ;
      RECT 166.665 20.655 166.835 20.825 ;
      RECT 166.665 23.375 166.835 23.545 ;
      RECT 166.665 26.095 166.835 26.265 ;
      RECT 166.665 28.815 166.835 28.985 ;
      RECT 166.665 31.535 166.835 31.705 ;
      RECT 166.665 34.255 166.835 34.425 ;
      RECT 166.665 36.975 166.835 37.145 ;
      RECT 166.665 39.695 166.835 39.865 ;
      RECT 166.665 42.415 166.835 42.585 ;
      RECT 166.665 45.135 166.835 45.305 ;
      RECT 166.665 47.855 166.835 48.025 ;
      RECT 166.665 50.575 166.835 50.745 ;
      RECT 166.665 53.295 166.835 53.465 ;
      RECT 166.665 56.015 166.835 56.185 ;
      RECT 166.665 58.735 166.835 58.905 ;
      RECT 166.205 9.775 166.375 9.945 ;
      RECT 166.205 12.495 166.375 12.665 ;
      RECT 166.205 15.215 166.375 15.385 ;
      RECT 166.205 17.935 166.375 18.105 ;
      RECT 166.205 20.655 166.375 20.825 ;
      RECT 166.205 23.375 166.375 23.545 ;
      RECT 166.205 26.095 166.375 26.265 ;
      RECT 166.205 28.815 166.375 28.985 ;
      RECT 166.205 31.535 166.375 31.705 ;
      RECT 166.205 34.255 166.375 34.425 ;
      RECT 166.205 36.975 166.375 37.145 ;
      RECT 166.205 39.695 166.375 39.865 ;
      RECT 166.205 42.415 166.375 42.585 ;
      RECT 166.205 45.135 166.375 45.305 ;
      RECT 166.205 47.855 166.375 48.025 ;
      RECT 166.205 50.575 166.375 50.745 ;
      RECT 166.205 53.295 166.375 53.465 ;
      RECT 166.205 56.015 166.375 56.185 ;
      RECT 166.205 58.735 166.375 58.905 ;
      RECT 165.745 9.775 165.915 9.945 ;
      RECT 165.745 12.495 165.915 12.665 ;
      RECT 165.745 15.215 165.915 15.385 ;
      RECT 165.745 17.935 165.915 18.105 ;
      RECT 165.745 20.655 165.915 20.825 ;
      RECT 165.745 23.375 165.915 23.545 ;
      RECT 165.745 26.095 165.915 26.265 ;
      RECT 165.745 28.815 165.915 28.985 ;
      RECT 165.745 31.535 165.915 31.705 ;
      RECT 165.745 34.255 165.915 34.425 ;
      RECT 165.745 36.975 165.915 37.145 ;
      RECT 165.745 39.695 165.915 39.865 ;
      RECT 165.745 42.415 165.915 42.585 ;
      RECT 165.745 45.135 165.915 45.305 ;
      RECT 165.745 47.855 165.915 48.025 ;
      RECT 165.745 50.575 165.915 50.745 ;
      RECT 165.745 53.295 165.915 53.465 ;
      RECT 165.745 56.015 165.915 56.185 ;
      RECT 165.745 58.735 165.915 58.905 ;
      RECT 165.285 9.775 165.455 9.945 ;
      RECT 165.285 12.495 165.455 12.665 ;
      RECT 165.285 15.215 165.455 15.385 ;
      RECT 165.285 17.935 165.455 18.105 ;
      RECT 165.285 20.655 165.455 20.825 ;
      RECT 165.285 23.375 165.455 23.545 ;
      RECT 165.285 26.095 165.455 26.265 ;
      RECT 165.285 28.815 165.455 28.985 ;
      RECT 165.285 31.535 165.455 31.705 ;
      RECT 165.285 34.255 165.455 34.425 ;
      RECT 165.285 36.975 165.455 37.145 ;
      RECT 165.285 39.695 165.455 39.865 ;
      RECT 165.285 42.415 165.455 42.585 ;
      RECT 165.285 45.135 165.455 45.305 ;
      RECT 165.285 47.855 165.455 48.025 ;
      RECT 165.285 50.575 165.455 50.745 ;
      RECT 165.285 53.295 165.455 53.465 ;
      RECT 165.285 56.015 165.455 56.185 ;
      RECT 165.285 58.735 165.455 58.905 ;
      RECT 165.11 16.065 165.28 16.235 ;
      RECT 164.825 9.775 164.995 9.945 ;
      RECT 164.825 12.495 164.995 12.665 ;
      RECT 164.825 15.215 164.995 15.385 ;
      RECT 164.825 17.935 164.995 18.105 ;
      RECT 164.825 20.655 164.995 20.825 ;
      RECT 164.825 23.375 164.995 23.545 ;
      RECT 164.825 26.095 164.995 26.265 ;
      RECT 164.825 28.815 164.995 28.985 ;
      RECT 164.825 31.535 164.995 31.705 ;
      RECT 164.825 34.255 164.995 34.425 ;
      RECT 164.825 36.975 164.995 37.145 ;
      RECT 164.825 39.695 164.995 39.865 ;
      RECT 164.825 42.415 164.995 42.585 ;
      RECT 164.825 45.135 164.995 45.305 ;
      RECT 164.825 47.855 164.995 48.025 ;
      RECT 164.825 50.575 164.995 50.745 ;
      RECT 164.825 53.295 164.995 53.465 ;
      RECT 164.825 56.015 164.995 56.185 ;
      RECT 164.825 58.735 164.995 58.905 ;
      RECT 164.595 16.405 164.765 16.575 ;
      RECT 164.365 9.775 164.535 9.945 ;
      RECT 164.365 12.495 164.535 12.665 ;
      RECT 164.365 15.215 164.535 15.385 ;
      RECT 164.365 17.935 164.535 18.105 ;
      RECT 164.365 20.655 164.535 20.825 ;
      RECT 164.365 23.375 164.535 23.545 ;
      RECT 164.365 26.095 164.535 26.265 ;
      RECT 164.365 28.815 164.535 28.985 ;
      RECT 164.365 31.535 164.535 31.705 ;
      RECT 164.365 34.255 164.535 34.425 ;
      RECT 164.365 36.975 164.535 37.145 ;
      RECT 164.365 39.695 164.535 39.865 ;
      RECT 164.365 42.415 164.535 42.585 ;
      RECT 164.365 45.135 164.535 45.305 ;
      RECT 164.365 47.855 164.535 48.025 ;
      RECT 164.365 50.575 164.535 50.745 ;
      RECT 164.365 53.295 164.535 53.465 ;
      RECT 164.365 56.015 164.535 56.185 ;
      RECT 164.365 58.735 164.535 58.905 ;
      RECT 163.905 9.775 164.075 9.945 ;
      RECT 163.905 12.495 164.075 12.665 ;
      RECT 163.905 15.215 164.075 15.385 ;
      RECT 163.905 17.935 164.075 18.105 ;
      RECT 163.905 20.655 164.075 20.825 ;
      RECT 163.905 23.375 164.075 23.545 ;
      RECT 163.905 26.095 164.075 26.265 ;
      RECT 163.905 28.815 164.075 28.985 ;
      RECT 163.905 31.535 164.075 31.705 ;
      RECT 163.905 34.255 164.075 34.425 ;
      RECT 163.905 36.975 164.075 37.145 ;
      RECT 163.905 39.695 164.075 39.865 ;
      RECT 163.905 42.415 164.075 42.585 ;
      RECT 163.905 45.135 164.075 45.305 ;
      RECT 163.905 47.855 164.075 48.025 ;
      RECT 163.905 50.575 164.075 50.745 ;
      RECT 163.905 53.295 164.075 53.465 ;
      RECT 163.905 56.015 164.075 56.185 ;
      RECT 163.905 58.735 164.075 58.905 ;
      RECT 163.83 17.085 164 17.255 ;
      RECT 163.445 9.775 163.615 9.945 ;
      RECT 163.445 12.495 163.615 12.665 ;
      RECT 163.445 15.215 163.615 15.385 ;
      RECT 163.445 17.935 163.615 18.105 ;
      RECT 163.445 20.655 163.615 20.825 ;
      RECT 163.445 23.375 163.615 23.545 ;
      RECT 163.445 26.095 163.615 26.265 ;
      RECT 163.445 28.815 163.615 28.985 ;
      RECT 163.445 31.535 163.615 31.705 ;
      RECT 163.445 34.255 163.615 34.425 ;
      RECT 163.445 36.975 163.615 37.145 ;
      RECT 163.445 39.695 163.615 39.865 ;
      RECT 163.445 42.415 163.615 42.585 ;
      RECT 163.445 45.135 163.615 45.305 ;
      RECT 163.445 47.855 163.615 48.025 ;
      RECT 163.445 50.575 163.615 50.745 ;
      RECT 163.445 53.295 163.615 53.465 ;
      RECT 163.445 56.015 163.615 56.185 ;
      RECT 163.445 58.735 163.615 58.905 ;
      RECT 163.405 16.405 163.575 16.575 ;
      RECT 163.01 16.065 163.18 16.235 ;
      RECT 162.985 9.775 163.155 9.945 ;
      RECT 162.985 12.495 163.155 12.665 ;
      RECT 162.985 15.215 163.155 15.385 ;
      RECT 162.985 17.935 163.155 18.105 ;
      RECT 162.985 20.655 163.155 20.825 ;
      RECT 162.985 23.375 163.155 23.545 ;
      RECT 162.985 26.095 163.155 26.265 ;
      RECT 162.985 28.815 163.155 28.985 ;
      RECT 162.985 31.535 163.155 31.705 ;
      RECT 162.985 34.255 163.155 34.425 ;
      RECT 162.985 36.975 163.155 37.145 ;
      RECT 162.985 39.695 163.155 39.865 ;
      RECT 162.985 42.415 163.155 42.585 ;
      RECT 162.985 45.135 163.155 45.305 ;
      RECT 162.985 47.855 163.155 48.025 ;
      RECT 162.985 50.575 163.155 50.745 ;
      RECT 162.985 53.295 163.155 53.465 ;
      RECT 162.985 56.015 163.155 56.185 ;
      RECT 162.985 58.735 163.155 58.905 ;
      RECT 162.525 9.775 162.695 9.945 ;
      RECT 162.525 12.495 162.695 12.665 ;
      RECT 162.525 15.215 162.695 15.385 ;
      RECT 162.525 16.745 162.695 16.915 ;
      RECT 162.525 17.935 162.695 18.105 ;
      RECT 162.525 20.655 162.695 20.825 ;
      RECT 162.525 23.375 162.695 23.545 ;
      RECT 162.525 26.095 162.695 26.265 ;
      RECT 162.525 28.815 162.695 28.985 ;
      RECT 162.525 31.535 162.695 31.705 ;
      RECT 162.525 34.255 162.695 34.425 ;
      RECT 162.525 36.975 162.695 37.145 ;
      RECT 162.525 39.695 162.695 39.865 ;
      RECT 162.525 42.415 162.695 42.585 ;
      RECT 162.525 45.135 162.695 45.305 ;
      RECT 162.525 47.855 162.695 48.025 ;
      RECT 162.525 50.575 162.695 50.745 ;
      RECT 162.525 53.295 162.695 53.465 ;
      RECT 162.525 56.015 162.695 56.185 ;
      RECT 162.525 58.735 162.695 58.905 ;
      RECT 162.065 9.775 162.235 9.945 ;
      RECT 162.065 11.305 162.235 11.475 ;
      RECT 162.065 12.495 162.235 12.665 ;
      RECT 162.065 15.215 162.235 15.385 ;
      RECT 162.065 17.935 162.235 18.105 ;
      RECT 162.065 20.655 162.235 20.825 ;
      RECT 162.065 23.375 162.235 23.545 ;
      RECT 162.065 26.095 162.235 26.265 ;
      RECT 162.065 28.815 162.235 28.985 ;
      RECT 162.065 31.535 162.235 31.705 ;
      RECT 162.065 34.255 162.235 34.425 ;
      RECT 162.065 36.975 162.235 37.145 ;
      RECT 162.065 39.695 162.235 39.865 ;
      RECT 162.065 42.415 162.235 42.585 ;
      RECT 162.065 45.135 162.235 45.305 ;
      RECT 162.065 47.855 162.235 48.025 ;
      RECT 162.065 50.575 162.235 50.745 ;
      RECT 162.065 53.295 162.235 53.465 ;
      RECT 162.065 56.015 162.235 56.185 ;
      RECT 162.065 58.735 162.235 58.905 ;
      RECT 161.605 9.775 161.775 9.945 ;
      RECT 161.605 12.495 161.775 12.665 ;
      RECT 161.605 15.215 161.775 15.385 ;
      RECT 161.605 17.935 161.775 18.105 ;
      RECT 161.605 20.655 161.775 20.825 ;
      RECT 161.605 23.375 161.775 23.545 ;
      RECT 161.605 26.095 161.775 26.265 ;
      RECT 161.605 28.815 161.775 28.985 ;
      RECT 161.605 31.535 161.775 31.705 ;
      RECT 161.605 34.255 161.775 34.425 ;
      RECT 161.605 36.975 161.775 37.145 ;
      RECT 161.605 39.695 161.775 39.865 ;
      RECT 161.605 42.415 161.775 42.585 ;
      RECT 161.605 45.135 161.775 45.305 ;
      RECT 161.605 47.855 161.775 48.025 ;
      RECT 161.605 50.575 161.775 50.745 ;
      RECT 161.605 53.295 161.775 53.465 ;
      RECT 161.605 56.015 161.775 56.185 ;
      RECT 161.605 58.735 161.775 58.905 ;
      RECT 161.145 9.775 161.315 9.945 ;
      RECT 161.145 12.495 161.315 12.665 ;
      RECT 161.145 15.215 161.315 15.385 ;
      RECT 161.145 17.935 161.315 18.105 ;
      RECT 161.145 20.655 161.315 20.825 ;
      RECT 161.145 23.375 161.315 23.545 ;
      RECT 161.145 26.095 161.315 26.265 ;
      RECT 161.145 28.815 161.315 28.985 ;
      RECT 161.145 31.535 161.315 31.705 ;
      RECT 161.145 34.255 161.315 34.425 ;
      RECT 161.145 36.975 161.315 37.145 ;
      RECT 161.145 39.695 161.315 39.865 ;
      RECT 161.145 42.415 161.315 42.585 ;
      RECT 161.145 45.135 161.315 45.305 ;
      RECT 161.145 47.855 161.315 48.025 ;
      RECT 161.145 50.575 161.315 50.745 ;
      RECT 161.145 53.295 161.315 53.465 ;
      RECT 161.145 56.015 161.315 56.185 ;
      RECT 161.145 58.735 161.315 58.905 ;
      RECT 160.685 9.775 160.855 9.945 ;
      RECT 160.685 12.495 160.855 12.665 ;
      RECT 160.685 15.215 160.855 15.385 ;
      RECT 160.685 17.935 160.855 18.105 ;
      RECT 160.685 20.655 160.855 20.825 ;
      RECT 160.685 23.375 160.855 23.545 ;
      RECT 160.685 26.095 160.855 26.265 ;
      RECT 160.685 28.815 160.855 28.985 ;
      RECT 160.685 31.535 160.855 31.705 ;
      RECT 160.685 34.255 160.855 34.425 ;
      RECT 160.685 36.975 160.855 37.145 ;
      RECT 160.685 39.695 160.855 39.865 ;
      RECT 160.685 42.415 160.855 42.585 ;
      RECT 160.685 45.135 160.855 45.305 ;
      RECT 160.685 47.855 160.855 48.025 ;
      RECT 160.685 50.575 160.855 50.745 ;
      RECT 160.685 53.295 160.855 53.465 ;
      RECT 160.685 56.015 160.855 56.185 ;
      RECT 160.685 58.735 160.855 58.905 ;
      RECT 160.225 9.775 160.395 9.945 ;
      RECT 160.225 12.495 160.395 12.665 ;
      RECT 160.225 15.215 160.395 15.385 ;
      RECT 160.225 17.935 160.395 18.105 ;
      RECT 160.225 20.655 160.395 20.825 ;
      RECT 160.225 23.375 160.395 23.545 ;
      RECT 160.225 26.095 160.395 26.265 ;
      RECT 160.225 28.815 160.395 28.985 ;
      RECT 160.225 31.535 160.395 31.705 ;
      RECT 160.225 34.255 160.395 34.425 ;
      RECT 160.225 36.975 160.395 37.145 ;
      RECT 160.225 39.695 160.395 39.865 ;
      RECT 160.225 42.415 160.395 42.585 ;
      RECT 160.225 45.135 160.395 45.305 ;
      RECT 160.225 47.855 160.395 48.025 ;
      RECT 160.225 50.575 160.395 50.745 ;
      RECT 160.225 53.295 160.395 53.465 ;
      RECT 160.225 56.015 160.395 56.185 ;
      RECT 160.225 58.735 160.395 58.905 ;
      RECT 159.765 9.775 159.935 9.945 ;
      RECT 159.765 12.495 159.935 12.665 ;
      RECT 159.765 15.215 159.935 15.385 ;
      RECT 159.765 17.935 159.935 18.105 ;
      RECT 159.765 20.655 159.935 20.825 ;
      RECT 159.765 23.375 159.935 23.545 ;
      RECT 159.765 26.095 159.935 26.265 ;
      RECT 159.765 28.815 159.935 28.985 ;
      RECT 159.765 31.535 159.935 31.705 ;
      RECT 159.765 34.255 159.935 34.425 ;
      RECT 159.765 36.975 159.935 37.145 ;
      RECT 159.765 39.695 159.935 39.865 ;
      RECT 159.765 42.415 159.935 42.585 ;
      RECT 159.765 45.135 159.935 45.305 ;
      RECT 159.765 47.855 159.935 48.025 ;
      RECT 159.765 50.575 159.935 50.745 ;
      RECT 159.765 53.295 159.935 53.465 ;
      RECT 159.765 56.015 159.935 56.185 ;
      RECT 159.765 58.735 159.935 58.905 ;
      RECT 159.305 9.775 159.475 9.945 ;
      RECT 159.305 12.495 159.475 12.665 ;
      RECT 159.305 15.215 159.475 15.385 ;
      RECT 159.305 17.935 159.475 18.105 ;
      RECT 159.305 20.655 159.475 20.825 ;
      RECT 159.305 23.375 159.475 23.545 ;
      RECT 159.305 26.095 159.475 26.265 ;
      RECT 159.305 28.815 159.475 28.985 ;
      RECT 159.305 31.535 159.475 31.705 ;
      RECT 159.305 34.255 159.475 34.425 ;
      RECT 159.305 36.975 159.475 37.145 ;
      RECT 159.305 39.695 159.475 39.865 ;
      RECT 159.305 42.415 159.475 42.585 ;
      RECT 159.305 45.135 159.475 45.305 ;
      RECT 159.305 47.855 159.475 48.025 ;
      RECT 159.305 50.575 159.475 50.745 ;
      RECT 159.305 53.295 159.475 53.465 ;
      RECT 159.305 56.015 159.475 56.185 ;
      RECT 159.305 58.735 159.475 58.905 ;
      RECT 158.845 9.775 159.015 9.945 ;
      RECT 158.845 12.495 159.015 12.665 ;
      RECT 158.845 15.215 159.015 15.385 ;
      RECT 158.845 17.935 159.015 18.105 ;
      RECT 158.845 20.655 159.015 20.825 ;
      RECT 158.845 23.375 159.015 23.545 ;
      RECT 158.845 26.095 159.015 26.265 ;
      RECT 158.845 28.815 159.015 28.985 ;
      RECT 158.845 31.535 159.015 31.705 ;
      RECT 158.845 34.255 159.015 34.425 ;
      RECT 158.845 36.975 159.015 37.145 ;
      RECT 158.845 39.695 159.015 39.865 ;
      RECT 158.845 42.415 159.015 42.585 ;
      RECT 158.845 45.135 159.015 45.305 ;
      RECT 158.845 47.855 159.015 48.025 ;
      RECT 158.845 50.575 159.015 50.745 ;
      RECT 158.845 53.295 159.015 53.465 ;
      RECT 158.845 56.015 159.015 56.185 ;
      RECT 158.845 58.735 159.015 58.905 ;
      RECT 158.385 9.775 158.555 9.945 ;
      RECT 158.385 12.495 158.555 12.665 ;
      RECT 158.385 15.215 158.555 15.385 ;
      RECT 158.385 17.935 158.555 18.105 ;
      RECT 158.385 20.655 158.555 20.825 ;
      RECT 158.385 23.375 158.555 23.545 ;
      RECT 158.385 26.095 158.555 26.265 ;
      RECT 158.385 28.815 158.555 28.985 ;
      RECT 158.385 31.535 158.555 31.705 ;
      RECT 158.385 34.255 158.555 34.425 ;
      RECT 158.385 34.765 158.555 34.935 ;
      RECT 158.385 36.975 158.555 37.145 ;
      RECT 158.385 39.695 158.555 39.865 ;
      RECT 158.385 42.415 158.555 42.585 ;
      RECT 158.385 45.135 158.555 45.305 ;
      RECT 158.385 47.855 158.555 48.025 ;
      RECT 158.385 50.575 158.555 50.745 ;
      RECT 158.385 53.295 158.555 53.465 ;
      RECT 158.385 56.015 158.555 56.185 ;
      RECT 158.385 58.735 158.555 58.905 ;
      RECT 157.925 9.775 158.095 9.945 ;
      RECT 157.925 12.495 158.095 12.665 ;
      RECT 157.925 15.215 158.095 15.385 ;
      RECT 157.925 17.935 158.095 18.105 ;
      RECT 157.925 20.655 158.095 20.825 ;
      RECT 157.925 23.375 158.095 23.545 ;
      RECT 157.925 26.095 158.095 26.265 ;
      RECT 157.925 28.815 158.095 28.985 ;
      RECT 157.925 29.325 158.095 29.495 ;
      RECT 157.925 31.535 158.095 31.705 ;
      RECT 157.925 34.255 158.095 34.425 ;
      RECT 157.925 36.975 158.095 37.145 ;
      RECT 157.925 39.695 158.095 39.865 ;
      RECT 157.925 42.415 158.095 42.585 ;
      RECT 157.925 45.135 158.095 45.305 ;
      RECT 157.925 47.855 158.095 48.025 ;
      RECT 157.925 50.575 158.095 50.745 ;
      RECT 157.925 53.295 158.095 53.465 ;
      RECT 157.925 56.015 158.095 56.185 ;
      RECT 157.925 58.735 158.095 58.905 ;
      RECT 157.465 9.775 157.635 9.945 ;
      RECT 157.465 12.495 157.635 12.665 ;
      RECT 157.465 15.215 157.635 15.385 ;
      RECT 157.465 17.935 157.635 18.105 ;
      RECT 157.465 20.655 157.635 20.825 ;
      RECT 157.465 23.375 157.635 23.545 ;
      RECT 157.465 26.095 157.635 26.265 ;
      RECT 157.465 28.815 157.635 28.985 ;
      RECT 157.465 31.535 157.635 31.705 ;
      RECT 157.465 34.255 157.635 34.425 ;
      RECT 157.465 36.975 157.635 37.145 ;
      RECT 157.465 39.695 157.635 39.865 ;
      RECT 157.465 42.415 157.635 42.585 ;
      RECT 157.465 45.135 157.635 45.305 ;
      RECT 157.465 47.855 157.635 48.025 ;
      RECT 157.465 50.575 157.635 50.745 ;
      RECT 157.465 53.295 157.635 53.465 ;
      RECT 157.465 56.015 157.635 56.185 ;
      RECT 157.465 58.735 157.635 58.905 ;
      RECT 157.005 9.775 157.175 9.945 ;
      RECT 157.005 12.495 157.175 12.665 ;
      RECT 157.005 15.215 157.175 15.385 ;
      RECT 157.005 17.935 157.175 18.105 ;
      RECT 157.005 20.655 157.175 20.825 ;
      RECT 157.005 23.375 157.175 23.545 ;
      RECT 157.005 26.095 157.175 26.265 ;
      RECT 157.005 28.815 157.175 28.985 ;
      RECT 157.005 31.535 157.175 31.705 ;
      RECT 157.005 34.255 157.175 34.425 ;
      RECT 157.005 36.975 157.175 37.145 ;
      RECT 157.005 39.695 157.175 39.865 ;
      RECT 157.005 42.415 157.175 42.585 ;
      RECT 157.005 45.135 157.175 45.305 ;
      RECT 157.005 47.855 157.175 48.025 ;
      RECT 157.005 50.575 157.175 50.745 ;
      RECT 157.005 53.295 157.175 53.465 ;
      RECT 157.005 56.015 157.175 56.185 ;
      RECT 157.005 58.735 157.175 58.905 ;
      RECT 156.545 9.775 156.715 9.945 ;
      RECT 156.545 12.495 156.715 12.665 ;
      RECT 156.545 15.215 156.715 15.385 ;
      RECT 156.545 17.935 156.715 18.105 ;
      RECT 156.545 20.655 156.715 20.825 ;
      RECT 156.545 23.375 156.715 23.545 ;
      RECT 156.545 26.095 156.715 26.265 ;
      RECT 156.545 28.815 156.715 28.985 ;
      RECT 156.545 31.535 156.715 31.705 ;
      RECT 156.545 34.255 156.715 34.425 ;
      RECT 156.545 36.975 156.715 37.145 ;
      RECT 156.545 39.695 156.715 39.865 ;
      RECT 156.545 42.415 156.715 42.585 ;
      RECT 156.545 45.135 156.715 45.305 ;
      RECT 156.545 47.855 156.715 48.025 ;
      RECT 156.545 50.575 156.715 50.745 ;
      RECT 156.545 53.295 156.715 53.465 ;
      RECT 156.545 56.015 156.715 56.185 ;
      RECT 156.545 58.735 156.715 58.905 ;
      RECT 156.085 9.775 156.255 9.945 ;
      RECT 156.085 12.495 156.255 12.665 ;
      RECT 156.085 15.215 156.255 15.385 ;
      RECT 156.085 17.935 156.255 18.105 ;
      RECT 156.085 18.445 156.255 18.615 ;
      RECT 156.085 20.655 156.255 20.825 ;
      RECT 156.085 23.375 156.255 23.545 ;
      RECT 156.085 26.095 156.255 26.265 ;
      RECT 156.085 28.305 156.255 28.475 ;
      RECT 156.085 28.815 156.255 28.985 ;
      RECT 156.085 31.535 156.255 31.705 ;
      RECT 156.085 33.745 156.255 33.915 ;
      RECT 156.085 34.255 156.255 34.425 ;
      RECT 156.085 36.975 156.255 37.145 ;
      RECT 156.085 39.695 156.255 39.865 ;
      RECT 156.085 42.415 156.255 42.585 ;
      RECT 156.085 45.135 156.255 45.305 ;
      RECT 156.085 47.855 156.255 48.025 ;
      RECT 156.085 50.575 156.255 50.745 ;
      RECT 156.085 53.295 156.255 53.465 ;
      RECT 156.085 56.015 156.255 56.185 ;
      RECT 156.085 58.735 156.255 58.905 ;
      RECT 156.075 35.785 156.245 35.955 ;
      RECT 155.64 36.125 155.81 36.295 ;
      RECT 155.625 9.775 155.795 9.945 ;
      RECT 155.625 12.495 155.795 12.665 ;
      RECT 155.625 15.215 155.795 15.385 ;
      RECT 155.625 17.935 155.795 18.105 ;
      RECT 155.625 20.655 155.795 20.825 ;
      RECT 155.625 23.375 155.795 23.545 ;
      RECT 155.625 26.095 155.795 26.265 ;
      RECT 155.625 28.815 155.795 28.985 ;
      RECT 155.625 31.535 155.795 31.705 ;
      RECT 155.625 34.255 155.795 34.425 ;
      RECT 155.625 36.975 155.795 37.145 ;
      RECT 155.625 39.695 155.795 39.865 ;
      RECT 155.625 42.415 155.795 42.585 ;
      RECT 155.625 45.135 155.795 45.305 ;
      RECT 155.625 47.855 155.795 48.025 ;
      RECT 155.625 50.575 155.795 50.745 ;
      RECT 155.625 53.295 155.795 53.465 ;
      RECT 155.625 56.015 155.795 56.185 ;
      RECT 155.625 58.735 155.795 58.905 ;
      RECT 155.615 30.345 155.785 30.515 ;
      RECT 155.395 19.125 155.565 19.295 ;
      RECT 155.395 27.625 155.565 27.795 ;
      RECT 155.395 33.065 155.565 33.235 ;
      RECT 155.18 30.685 155.35 30.855 ;
      RECT 155.165 9.775 155.335 9.945 ;
      RECT 155.165 12.495 155.335 12.665 ;
      RECT 155.165 15.215 155.335 15.385 ;
      RECT 155.165 17.935 155.335 18.105 ;
      RECT 155.165 20.655 155.335 20.825 ;
      RECT 155.165 23.375 155.335 23.545 ;
      RECT 155.165 26.095 155.335 26.265 ;
      RECT 155.165 28.815 155.335 28.985 ;
      RECT 155.165 31.535 155.335 31.705 ;
      RECT 155.165 34.255 155.335 34.425 ;
      RECT 155.165 36.975 155.335 37.145 ;
      RECT 155.165 39.695 155.335 39.865 ;
      RECT 155.165 42.415 155.335 42.585 ;
      RECT 155.165 45.135 155.335 45.305 ;
      RECT 155.165 47.855 155.335 48.025 ;
      RECT 155.165 50.575 155.335 50.745 ;
      RECT 155.165 53.295 155.335 53.465 ;
      RECT 155.165 56.015 155.335 56.185 ;
      RECT 155.165 58.735 155.335 58.905 ;
      RECT 154.705 9.775 154.875 9.945 ;
      RECT 154.705 12.495 154.875 12.665 ;
      RECT 154.705 15.215 154.875 15.385 ;
      RECT 154.705 15.725 154.875 15.895 ;
      RECT 154.705 17.935 154.875 18.105 ;
      RECT 154.705 18.785 154.875 18.955 ;
      RECT 154.705 20.655 154.875 20.825 ;
      RECT 154.705 23.375 154.875 23.545 ;
      RECT 154.705 26.095 154.875 26.265 ;
      RECT 154.705 27.625 154.875 27.795 ;
      RECT 154.705 28.815 154.875 28.985 ;
      RECT 154.705 31.535 154.875 31.705 ;
      RECT 154.705 33.405 154.875 33.575 ;
      RECT 154.705 34.255 154.875 34.425 ;
      RECT 154.705 36.975 154.875 37.145 ;
      RECT 154.705 39.695 154.875 39.865 ;
      RECT 154.705 42.415 154.875 42.585 ;
      RECT 154.705 45.135 154.875 45.305 ;
      RECT 154.705 47.855 154.875 48.025 ;
      RECT 154.705 50.575 154.875 50.745 ;
      RECT 154.705 53.295 154.875 53.465 ;
      RECT 154.705 56.015 154.875 56.185 ;
      RECT 154.705 58.735 154.875 58.905 ;
      RECT 154.245 9.775 154.415 9.945 ;
      RECT 154.245 12.495 154.415 12.665 ;
      RECT 154.245 15.215 154.415 15.385 ;
      RECT 154.245 17.935 154.415 18.105 ;
      RECT 154.245 18.785 154.415 18.955 ;
      RECT 154.245 20.655 154.415 20.825 ;
      RECT 154.245 22.185 154.415 22.355 ;
      RECT 154.245 23.375 154.415 23.545 ;
      RECT 154.245 26.095 154.415 26.265 ;
      RECT 154.245 27.965 154.415 28.135 ;
      RECT 154.245 28.815 154.415 28.985 ;
      RECT 154.245 31.535 154.415 31.705 ;
      RECT 154.245 33.065 154.415 33.235 ;
      RECT 154.245 34.255 154.415 34.425 ;
      RECT 154.245 36.975 154.415 37.145 ;
      RECT 154.245 39.695 154.415 39.865 ;
      RECT 154.245 42.415 154.415 42.585 ;
      RECT 154.245 45.135 154.415 45.305 ;
      RECT 154.245 47.855 154.415 48.025 ;
      RECT 154.245 50.575 154.415 50.745 ;
      RECT 154.245 53.295 154.415 53.465 ;
      RECT 154.245 56.015 154.415 56.185 ;
      RECT 154.245 58.735 154.415 58.905 ;
      RECT 154.07 36.125 154.24 36.295 ;
      RECT 153.785 9.775 153.955 9.945 ;
      RECT 153.785 12.495 153.955 12.665 ;
      RECT 153.785 15.215 153.955 15.385 ;
      RECT 153.785 17.935 153.955 18.105 ;
      RECT 153.785 20.655 153.955 20.825 ;
      RECT 153.785 23.375 153.955 23.545 ;
      RECT 153.785 26.095 153.955 26.265 ;
      RECT 153.785 28.815 153.955 28.985 ;
      RECT 153.785 31.535 153.955 31.705 ;
      RECT 153.785 34.255 153.955 34.425 ;
      RECT 153.785 36.975 153.955 37.145 ;
      RECT 153.785 39.695 153.955 39.865 ;
      RECT 153.785 42.415 153.955 42.585 ;
      RECT 153.785 45.135 153.955 45.305 ;
      RECT 153.785 47.855 153.955 48.025 ;
      RECT 153.785 50.575 153.955 50.745 ;
      RECT 153.785 53.295 153.955 53.465 ;
      RECT 153.785 56.015 153.955 56.185 ;
      RECT 153.785 58.735 153.955 58.905 ;
      RECT 153.61 30.685 153.78 30.855 ;
      RECT 153.555 27.625 153.725 27.795 ;
      RECT 153.555 33.065 153.725 33.235 ;
      RECT 153.555 35.785 153.725 35.955 ;
      RECT 153.465 19.125 153.635 19.295 ;
      RECT 153.325 9.775 153.495 9.945 ;
      RECT 153.325 11.305 153.495 11.475 ;
      RECT 153.325 12.495 153.495 12.665 ;
      RECT 153.325 15.215 153.495 15.385 ;
      RECT 153.325 17.935 153.495 18.105 ;
      RECT 153.325 20.655 153.495 20.825 ;
      RECT 153.325 23.375 153.495 23.545 ;
      RECT 153.325 26.095 153.495 26.265 ;
      RECT 153.325 28.815 153.495 28.985 ;
      RECT 153.325 31.535 153.495 31.705 ;
      RECT 153.325 34.255 153.495 34.425 ;
      RECT 153.325 36.975 153.495 37.145 ;
      RECT 153.325 39.695 153.495 39.865 ;
      RECT 153.325 42.415 153.495 42.585 ;
      RECT 153.325 45.135 153.495 45.305 ;
      RECT 153.325 47.855 153.495 48.025 ;
      RECT 153.325 50.575 153.495 50.745 ;
      RECT 153.325 53.295 153.495 53.465 ;
      RECT 153.325 56.015 153.495 56.185 ;
      RECT 153.325 58.735 153.495 58.905 ;
      RECT 153.095 30.345 153.265 30.515 ;
      RECT 152.865 9.775 153.035 9.945 ;
      RECT 152.865 12.495 153.035 12.665 ;
      RECT 152.865 15.215 153.035 15.385 ;
      RECT 152.865 17.935 153.035 18.105 ;
      RECT 152.865 19.125 153.035 19.295 ;
      RECT 152.865 20.655 153.035 20.825 ;
      RECT 152.865 23.375 153.035 23.545 ;
      RECT 152.865 26.095 153.035 26.265 ;
      RECT 152.865 27.625 153.035 27.795 ;
      RECT 152.865 28.815 153.035 28.985 ;
      RECT 152.865 31.535 153.035 31.705 ;
      RECT 152.865 33.065 153.035 33.235 ;
      RECT 152.865 34.255 153.035 34.425 ;
      RECT 152.865 36.975 153.035 37.145 ;
      RECT 152.865 39.695 153.035 39.865 ;
      RECT 152.865 42.415 153.035 42.585 ;
      RECT 152.865 45.135 153.035 45.305 ;
      RECT 152.865 47.855 153.035 48.025 ;
      RECT 152.865 50.575 153.035 50.745 ;
      RECT 152.865 53.295 153.035 53.465 ;
      RECT 152.865 56.015 153.035 56.185 ;
      RECT 152.865 58.735 153.035 58.905 ;
      RECT 152.79 35.445 152.96 35.615 ;
      RECT 152.405 9.775 152.575 9.945 ;
      RECT 152.405 12.495 152.575 12.665 ;
      RECT 152.405 15.215 152.575 15.385 ;
      RECT 152.405 17.935 152.575 18.105 ;
      RECT 152.405 20.655 152.575 20.825 ;
      RECT 152.405 23.375 152.575 23.545 ;
      RECT 152.405 26.095 152.575 26.265 ;
      RECT 152.405 28.815 152.575 28.985 ;
      RECT 152.405 31.535 152.575 31.705 ;
      RECT 152.405 34.255 152.575 34.425 ;
      RECT 152.405 36.975 152.575 37.145 ;
      RECT 152.405 39.695 152.575 39.865 ;
      RECT 152.405 42.415 152.575 42.585 ;
      RECT 152.405 45.135 152.575 45.305 ;
      RECT 152.405 47.855 152.575 48.025 ;
      RECT 152.405 50.575 152.575 50.745 ;
      RECT 152.405 53.295 152.575 53.465 ;
      RECT 152.405 56.015 152.575 56.185 ;
      RECT 152.405 58.735 152.575 58.905 ;
      RECT 152.395 16.405 152.565 16.575 ;
      RECT 152.365 35.785 152.535 35.955 ;
      RECT 152.33 29.665 152.5 29.835 ;
      RECT 151.97 36.125 152.14 36.295 ;
      RECT 151.96 16.065 152.13 16.235 ;
      RECT 151.945 9.775 152.115 9.945 ;
      RECT 151.945 12.495 152.115 12.665 ;
      RECT 151.945 15.215 152.115 15.385 ;
      RECT 151.945 17.935 152.115 18.105 ;
      RECT 151.945 20.655 152.115 20.825 ;
      RECT 151.945 23.375 152.115 23.545 ;
      RECT 151.945 26.095 152.115 26.265 ;
      RECT 151.945 28.815 152.115 28.985 ;
      RECT 151.945 31.535 152.115 31.705 ;
      RECT 151.945 34.255 152.115 34.425 ;
      RECT 151.945 36.975 152.115 37.145 ;
      RECT 151.945 39.695 152.115 39.865 ;
      RECT 151.945 42.415 152.115 42.585 ;
      RECT 151.945 45.135 152.115 45.305 ;
      RECT 151.945 47.855 152.115 48.025 ;
      RECT 151.945 50.575 152.115 50.745 ;
      RECT 151.945 53.295 152.115 53.465 ;
      RECT 151.945 56.015 152.115 56.185 ;
      RECT 151.945 58.735 152.115 58.905 ;
      RECT 151.905 30.345 152.075 30.515 ;
      RECT 151.51 30.685 151.68 30.855 ;
      RECT 151.485 9.775 151.655 9.945 ;
      RECT 151.485 12.495 151.655 12.665 ;
      RECT 151.485 15.215 151.655 15.385 ;
      RECT 151.485 17.935 151.655 18.105 ;
      RECT 151.485 20.655 151.655 20.825 ;
      RECT 151.485 23.375 151.655 23.545 ;
      RECT 151.485 26.095 151.655 26.265 ;
      RECT 151.485 28.815 151.655 28.985 ;
      RECT 151.485 31.535 151.655 31.705 ;
      RECT 151.485 34.255 151.655 34.425 ;
      RECT 151.485 35.445 151.655 35.615 ;
      RECT 151.485 36.975 151.655 37.145 ;
      RECT 151.485 39.695 151.655 39.865 ;
      RECT 151.485 42.415 151.655 42.585 ;
      RECT 151.485 45.135 151.655 45.305 ;
      RECT 151.485 47.855 151.655 48.025 ;
      RECT 151.485 50.575 151.655 50.745 ;
      RECT 151.485 53.295 151.655 53.465 ;
      RECT 151.485 56.015 151.655 56.185 ;
      RECT 151.485 58.735 151.655 58.905 ;
      RECT 151.025 9.775 151.195 9.945 ;
      RECT 151.025 12.495 151.195 12.665 ;
      RECT 151.025 15.215 151.195 15.385 ;
      RECT 151.025 17.935 151.195 18.105 ;
      RECT 151.025 18.445 151.195 18.615 ;
      RECT 151.025 20.655 151.195 20.825 ;
      RECT 151.025 23.375 151.195 23.545 ;
      RECT 151.025 26.095 151.195 26.265 ;
      RECT 151.025 28.815 151.195 28.985 ;
      RECT 151.025 30.005 151.195 30.175 ;
      RECT 151.025 31.535 151.195 31.705 ;
      RECT 151.025 34.255 151.195 34.425 ;
      RECT 151.025 36.975 151.195 37.145 ;
      RECT 151.025 39.695 151.195 39.865 ;
      RECT 151.025 42.415 151.195 42.585 ;
      RECT 151.025 45.135 151.195 45.305 ;
      RECT 151.025 47.855 151.195 48.025 ;
      RECT 151.025 50.575 151.195 50.745 ;
      RECT 151.025 53.295 151.195 53.465 ;
      RECT 151.025 56.015 151.195 56.185 ;
      RECT 151.025 58.735 151.195 58.905 ;
      RECT 150.565 9.775 150.735 9.945 ;
      RECT 150.565 12.495 150.735 12.665 ;
      RECT 150.565 15.215 150.735 15.385 ;
      RECT 150.565 17.935 150.735 18.105 ;
      RECT 150.565 20.655 150.735 20.825 ;
      RECT 150.565 23.375 150.735 23.545 ;
      RECT 150.565 26.095 150.735 26.265 ;
      RECT 150.565 28.815 150.735 28.985 ;
      RECT 150.565 31.535 150.735 31.705 ;
      RECT 150.565 34.255 150.735 34.425 ;
      RECT 150.565 36.975 150.735 37.145 ;
      RECT 150.565 39.695 150.735 39.865 ;
      RECT 150.565 42.415 150.735 42.585 ;
      RECT 150.565 45.135 150.735 45.305 ;
      RECT 150.565 47.855 150.735 48.025 ;
      RECT 150.565 50.575 150.735 50.745 ;
      RECT 150.565 53.295 150.735 53.465 ;
      RECT 150.565 56.015 150.735 56.185 ;
      RECT 150.565 58.735 150.735 58.905 ;
      RECT 150.39 16.065 150.56 16.235 ;
      RECT 150.335 19.125 150.505 19.295 ;
      RECT 150.105 9.775 150.275 9.945 ;
      RECT 150.105 12.495 150.275 12.665 ;
      RECT 150.105 15.215 150.275 15.385 ;
      RECT 150.105 17.935 150.275 18.105 ;
      RECT 150.105 20.655 150.275 20.825 ;
      RECT 150.105 23.375 150.275 23.545 ;
      RECT 150.105 26.095 150.275 26.265 ;
      RECT 150.105 28.815 150.275 28.985 ;
      RECT 150.105 31.535 150.275 31.705 ;
      RECT 150.105 34.255 150.275 34.425 ;
      RECT 150.105 36.975 150.275 37.145 ;
      RECT 150.105 39.695 150.275 39.865 ;
      RECT 150.105 42.415 150.275 42.585 ;
      RECT 150.105 45.135 150.275 45.305 ;
      RECT 150.105 47.855 150.275 48.025 ;
      RECT 150.105 50.575 150.275 50.745 ;
      RECT 150.105 53.295 150.275 53.465 ;
      RECT 150.105 56.015 150.275 56.185 ;
      RECT 150.105 58.735 150.275 58.905 ;
      RECT 149.875 16.405 150.045 16.575 ;
      RECT 149.645 9.775 149.815 9.945 ;
      RECT 149.645 12.495 149.815 12.665 ;
      RECT 149.645 15.215 149.815 15.385 ;
      RECT 149.645 17.935 149.815 18.105 ;
      RECT 149.645 19.125 149.815 19.295 ;
      RECT 149.645 20.655 149.815 20.825 ;
      RECT 149.645 23.375 149.815 23.545 ;
      RECT 149.645 26.095 149.815 26.265 ;
      RECT 149.645 28.815 149.815 28.985 ;
      RECT 149.645 31.535 149.815 31.705 ;
      RECT 149.645 34.255 149.815 34.425 ;
      RECT 149.645 36.975 149.815 37.145 ;
      RECT 149.645 39.695 149.815 39.865 ;
      RECT 149.645 42.415 149.815 42.585 ;
      RECT 149.645 45.135 149.815 45.305 ;
      RECT 149.645 47.855 149.815 48.025 ;
      RECT 149.645 50.575 149.815 50.745 ;
      RECT 149.645 53.295 149.815 53.465 ;
      RECT 149.645 56.015 149.815 56.185 ;
      RECT 149.645 58.735 149.815 58.905 ;
      RECT 149.185 9.775 149.355 9.945 ;
      RECT 149.185 12.495 149.355 12.665 ;
      RECT 149.185 15.215 149.355 15.385 ;
      RECT 149.185 17.935 149.355 18.105 ;
      RECT 149.185 18.785 149.355 18.955 ;
      RECT 149.185 20.655 149.355 20.825 ;
      RECT 149.185 23.375 149.355 23.545 ;
      RECT 149.185 26.095 149.355 26.265 ;
      RECT 149.185 28.815 149.355 28.985 ;
      RECT 149.185 31.535 149.355 31.705 ;
      RECT 149.185 34.255 149.355 34.425 ;
      RECT 149.185 36.975 149.355 37.145 ;
      RECT 149.185 39.695 149.355 39.865 ;
      RECT 149.185 42.415 149.355 42.585 ;
      RECT 149.185 45.135 149.355 45.305 ;
      RECT 149.185 47.855 149.355 48.025 ;
      RECT 149.185 50.575 149.355 50.745 ;
      RECT 149.185 53.295 149.355 53.465 ;
      RECT 149.185 56.015 149.355 56.185 ;
      RECT 149.185 58.735 149.355 58.905 ;
      RECT 149.11 17.085 149.28 17.255 ;
      RECT 148.725 9.775 148.895 9.945 ;
      RECT 148.725 12.495 148.895 12.665 ;
      RECT 148.725 15.215 148.895 15.385 ;
      RECT 148.725 17.935 148.895 18.105 ;
      RECT 148.725 20.655 148.895 20.825 ;
      RECT 148.725 21.505 148.895 21.675 ;
      RECT 148.725 22.865 148.895 23.035 ;
      RECT 148.725 23.375 148.895 23.545 ;
      RECT 148.725 26.095 148.895 26.265 ;
      RECT 148.725 28.815 148.895 28.985 ;
      RECT 148.725 31.535 148.895 31.705 ;
      RECT 148.725 34.255 148.895 34.425 ;
      RECT 148.725 36.975 148.895 37.145 ;
      RECT 148.725 39.695 148.895 39.865 ;
      RECT 148.725 42.415 148.895 42.585 ;
      RECT 148.725 45.135 148.895 45.305 ;
      RECT 148.725 47.855 148.895 48.025 ;
      RECT 148.725 50.575 148.895 50.745 ;
      RECT 148.725 53.295 148.895 53.465 ;
      RECT 148.725 56.015 148.895 56.185 ;
      RECT 148.725 58.735 148.895 58.905 ;
      RECT 148.685 16.405 148.855 16.575 ;
      RECT 148.495 19.125 148.665 19.295 ;
      RECT 148.29 16.065 148.46 16.235 ;
      RECT 148.265 9.775 148.435 9.945 ;
      RECT 148.265 12.495 148.435 12.665 ;
      RECT 148.265 15.215 148.435 15.385 ;
      RECT 148.265 17.935 148.435 18.105 ;
      RECT 148.265 20.655 148.435 20.825 ;
      RECT 148.265 23.375 148.435 23.545 ;
      RECT 148.265 26.095 148.435 26.265 ;
      RECT 148.265 28.815 148.435 28.985 ;
      RECT 148.265 31.535 148.435 31.705 ;
      RECT 148.265 34.255 148.435 34.425 ;
      RECT 148.265 36.975 148.435 37.145 ;
      RECT 148.265 39.695 148.435 39.865 ;
      RECT 148.265 42.415 148.435 42.585 ;
      RECT 148.265 45.135 148.435 45.305 ;
      RECT 148.265 47.855 148.435 48.025 ;
      RECT 148.265 50.575 148.435 50.745 ;
      RECT 148.265 53.295 148.435 53.465 ;
      RECT 148.265 56.015 148.435 56.185 ;
      RECT 148.265 58.735 148.435 58.905 ;
      RECT 147.805 9.775 147.975 9.945 ;
      RECT 147.805 12.495 147.975 12.665 ;
      RECT 147.805 15.215 147.975 15.385 ;
      RECT 147.805 16.745 147.975 16.915 ;
      RECT 147.805 17.935 147.975 18.105 ;
      RECT 147.805 19.125 147.975 19.295 ;
      RECT 147.805 20.655 147.975 20.825 ;
      RECT 147.805 23.375 147.975 23.545 ;
      RECT 147.805 26.095 147.975 26.265 ;
      RECT 147.805 28.815 147.975 28.985 ;
      RECT 147.805 31.535 147.975 31.705 ;
      RECT 147.805 34.255 147.975 34.425 ;
      RECT 147.805 36.975 147.975 37.145 ;
      RECT 147.805 39.695 147.975 39.865 ;
      RECT 147.805 42.415 147.975 42.585 ;
      RECT 147.805 45.135 147.975 45.305 ;
      RECT 147.805 47.855 147.975 48.025 ;
      RECT 147.805 50.575 147.975 50.745 ;
      RECT 147.805 53.295 147.975 53.465 ;
      RECT 147.805 56.015 147.975 56.185 ;
      RECT 147.805 58.735 147.975 58.905 ;
      RECT 147.345 9.775 147.515 9.945 ;
      RECT 147.345 12.495 147.515 12.665 ;
      RECT 147.345 15.215 147.515 15.385 ;
      RECT 147.345 17.935 147.515 18.105 ;
      RECT 147.345 20.655 147.515 20.825 ;
      RECT 147.345 23.375 147.515 23.545 ;
      RECT 147.345 26.095 147.515 26.265 ;
      RECT 147.345 28.815 147.515 28.985 ;
      RECT 147.345 31.535 147.515 31.705 ;
      RECT 147.345 34.255 147.515 34.425 ;
      RECT 147.345 36.975 147.515 37.145 ;
      RECT 147.345 39.695 147.515 39.865 ;
      RECT 147.345 42.415 147.515 42.585 ;
      RECT 147.345 45.135 147.515 45.305 ;
      RECT 147.345 47.855 147.515 48.025 ;
      RECT 147.345 50.575 147.515 50.745 ;
      RECT 147.345 53.295 147.515 53.465 ;
      RECT 147.345 56.015 147.515 56.185 ;
      RECT 147.345 58.735 147.515 58.905 ;
      RECT 146.885 9.775 147.055 9.945 ;
      RECT 146.885 12.495 147.055 12.665 ;
      RECT 146.885 15.215 147.055 15.385 ;
      RECT 146.885 17.935 147.055 18.105 ;
      RECT 146.885 20.655 147.055 20.825 ;
      RECT 146.885 23.375 147.055 23.545 ;
      RECT 146.885 26.095 147.055 26.265 ;
      RECT 146.885 28.815 147.055 28.985 ;
      RECT 146.885 31.535 147.055 31.705 ;
      RECT 146.885 34.255 147.055 34.425 ;
      RECT 146.885 36.975 147.055 37.145 ;
      RECT 146.885 39.695 147.055 39.865 ;
      RECT 146.885 42.415 147.055 42.585 ;
      RECT 146.885 45.135 147.055 45.305 ;
      RECT 146.885 47.855 147.055 48.025 ;
      RECT 146.885 50.575 147.055 50.745 ;
      RECT 146.885 53.295 147.055 53.465 ;
      RECT 146.885 56.015 147.055 56.185 ;
      RECT 146.885 58.735 147.055 58.905 ;
      RECT 146.425 9.775 146.595 9.945 ;
      RECT 146.425 12.495 146.595 12.665 ;
      RECT 146.425 15.215 146.595 15.385 ;
      RECT 146.425 17.935 146.595 18.105 ;
      RECT 146.425 20.655 146.595 20.825 ;
      RECT 146.425 23.375 146.595 23.545 ;
      RECT 146.425 26.095 146.595 26.265 ;
      RECT 146.425 28.815 146.595 28.985 ;
      RECT 146.425 31.535 146.595 31.705 ;
      RECT 146.425 34.255 146.595 34.425 ;
      RECT 146.425 36.975 146.595 37.145 ;
      RECT 146.425 39.695 146.595 39.865 ;
      RECT 146.425 42.415 146.595 42.585 ;
      RECT 146.425 45.135 146.595 45.305 ;
      RECT 146.425 47.855 146.595 48.025 ;
      RECT 146.425 50.575 146.595 50.745 ;
      RECT 146.425 53.295 146.595 53.465 ;
      RECT 146.425 56.015 146.595 56.185 ;
      RECT 146.425 58.735 146.595 58.905 ;
      RECT 145.965 9.775 146.135 9.945 ;
      RECT 145.965 12.495 146.135 12.665 ;
      RECT 145.965 15.215 146.135 15.385 ;
      RECT 145.965 17.935 146.135 18.105 ;
      RECT 145.965 20.655 146.135 20.825 ;
      RECT 145.965 23.375 146.135 23.545 ;
      RECT 145.965 26.095 146.135 26.265 ;
      RECT 145.965 28.815 146.135 28.985 ;
      RECT 145.965 31.535 146.135 31.705 ;
      RECT 145.965 34.255 146.135 34.425 ;
      RECT 145.965 36.975 146.135 37.145 ;
      RECT 145.965 39.695 146.135 39.865 ;
      RECT 145.965 42.415 146.135 42.585 ;
      RECT 145.965 45.135 146.135 45.305 ;
      RECT 145.965 47.855 146.135 48.025 ;
      RECT 145.965 50.575 146.135 50.745 ;
      RECT 145.965 53.295 146.135 53.465 ;
      RECT 145.965 56.015 146.135 56.185 ;
      RECT 145.965 58.735 146.135 58.905 ;
      RECT 145.505 9.775 145.675 9.945 ;
      RECT 145.505 12.495 145.675 12.665 ;
      RECT 145.505 15.215 145.675 15.385 ;
      RECT 145.505 17.935 145.675 18.105 ;
      RECT 145.505 20.655 145.675 20.825 ;
      RECT 145.505 23.375 145.675 23.545 ;
      RECT 145.505 26.095 145.675 26.265 ;
      RECT 145.505 26.605 145.675 26.775 ;
      RECT 145.505 28.305 145.675 28.475 ;
      RECT 145.505 28.815 145.675 28.985 ;
      RECT 145.505 31.535 145.675 31.705 ;
      RECT 145.505 34.255 145.675 34.425 ;
      RECT 145.505 36.975 145.675 37.145 ;
      RECT 145.505 39.695 145.675 39.865 ;
      RECT 145.505 42.415 145.675 42.585 ;
      RECT 145.505 45.135 145.675 45.305 ;
      RECT 145.505 47.855 145.675 48.025 ;
      RECT 145.505 50.575 145.675 50.745 ;
      RECT 145.505 53.295 145.675 53.465 ;
      RECT 145.505 56.015 145.675 56.185 ;
      RECT 145.505 58.735 145.675 58.905 ;
      RECT 145.045 9.775 145.215 9.945 ;
      RECT 145.045 12.495 145.215 12.665 ;
      RECT 145.045 15.215 145.215 15.385 ;
      RECT 145.045 17.935 145.215 18.105 ;
      RECT 145.045 20.655 145.215 20.825 ;
      RECT 145.045 22.865 145.215 23.035 ;
      RECT 145.045 23.375 145.215 23.545 ;
      RECT 145.045 26.095 145.215 26.265 ;
      RECT 145.045 28.815 145.215 28.985 ;
      RECT 145.045 31.535 145.215 31.705 ;
      RECT 145.045 34.255 145.215 34.425 ;
      RECT 145.045 36.975 145.215 37.145 ;
      RECT 145.045 39.695 145.215 39.865 ;
      RECT 145.045 42.415 145.215 42.585 ;
      RECT 145.045 45.135 145.215 45.305 ;
      RECT 145.045 47.855 145.215 48.025 ;
      RECT 145.045 50.575 145.215 50.745 ;
      RECT 145.045 53.295 145.215 53.465 ;
      RECT 145.045 56.015 145.215 56.185 ;
      RECT 145.045 58.735 145.215 58.905 ;
      RECT 144.585 9.775 144.755 9.945 ;
      RECT 144.585 12.495 144.755 12.665 ;
      RECT 144.585 15.215 144.755 15.385 ;
      RECT 144.585 17.935 144.755 18.105 ;
      RECT 144.585 20.655 144.755 20.825 ;
      RECT 144.585 23.375 144.755 23.545 ;
      RECT 144.585 26.095 144.755 26.265 ;
      RECT 144.585 28.815 144.755 28.985 ;
      RECT 144.585 31.535 144.755 31.705 ;
      RECT 144.585 34.255 144.755 34.425 ;
      RECT 144.585 36.975 144.755 37.145 ;
      RECT 144.585 39.695 144.755 39.865 ;
      RECT 144.585 42.415 144.755 42.585 ;
      RECT 144.585 45.135 144.755 45.305 ;
      RECT 144.585 47.855 144.755 48.025 ;
      RECT 144.585 50.575 144.755 50.745 ;
      RECT 144.585 53.295 144.755 53.465 ;
      RECT 144.585 56.015 144.755 56.185 ;
      RECT 144.585 58.735 144.755 58.905 ;
      RECT 144.125 9.775 144.295 9.945 ;
      RECT 144.125 12.495 144.295 12.665 ;
      RECT 144.125 15.215 144.295 15.385 ;
      RECT 144.125 17.935 144.295 18.105 ;
      RECT 144.125 20.655 144.295 20.825 ;
      RECT 144.125 23.375 144.295 23.545 ;
      RECT 144.125 24.565 144.295 24.735 ;
      RECT 144.125 26.095 144.295 26.265 ;
      RECT 144.125 28.815 144.295 28.985 ;
      RECT 144.125 31.535 144.295 31.705 ;
      RECT 144.125 34.255 144.295 34.425 ;
      RECT 144.125 36.975 144.295 37.145 ;
      RECT 144.125 39.695 144.295 39.865 ;
      RECT 144.125 42.415 144.295 42.585 ;
      RECT 144.125 45.135 144.295 45.305 ;
      RECT 144.125 47.855 144.295 48.025 ;
      RECT 144.125 50.575 144.295 50.745 ;
      RECT 144.125 53.295 144.295 53.465 ;
      RECT 144.125 56.015 144.295 56.185 ;
      RECT 144.125 58.735 144.295 58.905 ;
      RECT 143.665 9.775 143.835 9.945 ;
      RECT 143.665 12.495 143.835 12.665 ;
      RECT 143.665 15.215 143.835 15.385 ;
      RECT 143.665 17.935 143.835 18.105 ;
      RECT 143.665 20.655 143.835 20.825 ;
      RECT 143.665 23.375 143.835 23.545 ;
      RECT 143.665 26.095 143.835 26.265 ;
      RECT 143.665 28.815 143.835 28.985 ;
      RECT 143.665 31.535 143.835 31.705 ;
      RECT 143.665 34.255 143.835 34.425 ;
      RECT 143.665 36.975 143.835 37.145 ;
      RECT 143.665 39.695 143.835 39.865 ;
      RECT 143.665 42.415 143.835 42.585 ;
      RECT 143.665 45.135 143.835 45.305 ;
      RECT 143.665 47.855 143.835 48.025 ;
      RECT 143.665 50.575 143.835 50.745 ;
      RECT 143.665 53.295 143.835 53.465 ;
      RECT 143.665 56.015 143.835 56.185 ;
      RECT 143.665 58.735 143.835 58.905 ;
      RECT 143.52 24.565 143.69 24.735 ;
      RECT 143.205 9.775 143.375 9.945 ;
      RECT 143.205 12.495 143.375 12.665 ;
      RECT 143.205 15.215 143.375 15.385 ;
      RECT 143.205 17.935 143.375 18.105 ;
      RECT 143.205 20.655 143.375 20.825 ;
      RECT 143.205 21.505 143.375 21.675 ;
      RECT 143.205 23.375 143.375 23.545 ;
      RECT 143.205 26.095 143.375 26.265 ;
      RECT 143.205 28.815 143.375 28.985 ;
      RECT 143.205 31.535 143.375 31.705 ;
      RECT 143.205 34.255 143.375 34.425 ;
      RECT 143.205 36.975 143.375 37.145 ;
      RECT 143.205 39.695 143.375 39.865 ;
      RECT 143.205 42.415 143.375 42.585 ;
      RECT 143.205 45.135 143.375 45.305 ;
      RECT 143.205 47.855 143.375 48.025 ;
      RECT 143.205 50.575 143.375 50.745 ;
      RECT 143.205 53.295 143.375 53.465 ;
      RECT 143.205 56.015 143.375 56.185 ;
      RECT 143.205 58.735 143.375 58.905 ;
      RECT 143.195 27.285 143.365 27.455 ;
      RECT 142.76 26.945 142.93 27.115 ;
      RECT 142.745 9.775 142.915 9.945 ;
      RECT 142.745 12.495 142.915 12.665 ;
      RECT 142.745 15.215 142.915 15.385 ;
      RECT 142.745 17.935 142.915 18.105 ;
      RECT 142.745 20.655 142.915 20.825 ;
      RECT 142.745 23.375 142.915 23.545 ;
      RECT 142.745 24.565 142.915 24.735 ;
      RECT 142.745 26.095 142.915 26.265 ;
      RECT 142.745 28.815 142.915 28.985 ;
      RECT 142.745 31.535 142.915 31.705 ;
      RECT 142.745 34.255 142.915 34.425 ;
      RECT 142.745 36.975 142.915 37.145 ;
      RECT 142.745 39.695 142.915 39.865 ;
      RECT 142.745 42.415 142.915 42.585 ;
      RECT 142.745 45.135 142.915 45.305 ;
      RECT 142.745 47.855 142.915 48.025 ;
      RECT 142.745 50.575 142.915 50.745 ;
      RECT 142.745 53.295 142.915 53.465 ;
      RECT 142.745 56.015 142.915 56.185 ;
      RECT 142.745 58.735 142.915 58.905 ;
      RECT 142.285 9.775 142.455 9.945 ;
      RECT 142.285 12.495 142.455 12.665 ;
      RECT 142.285 15.215 142.455 15.385 ;
      RECT 142.285 17.935 142.455 18.105 ;
      RECT 142.285 20.655 142.455 20.825 ;
      RECT 142.285 23.375 142.455 23.545 ;
      RECT 142.285 24.225 142.455 24.395 ;
      RECT 142.285 26.095 142.455 26.265 ;
      RECT 142.285 28.815 142.455 28.985 ;
      RECT 142.285 31.535 142.455 31.705 ;
      RECT 142.285 34.255 142.455 34.425 ;
      RECT 142.285 36.975 142.455 37.145 ;
      RECT 142.285 39.695 142.455 39.865 ;
      RECT 142.285 42.415 142.455 42.585 ;
      RECT 142.285 45.135 142.455 45.305 ;
      RECT 142.285 47.855 142.455 48.025 ;
      RECT 142.285 50.575 142.455 50.745 ;
      RECT 142.285 53.295 142.455 53.465 ;
      RECT 142.285 56.015 142.455 56.185 ;
      RECT 142.285 58.735 142.455 58.905 ;
      RECT 141.825 9.775 141.995 9.945 ;
      RECT 141.825 12.495 141.995 12.665 ;
      RECT 141.825 15.215 141.995 15.385 ;
      RECT 141.825 17.935 141.995 18.105 ;
      RECT 141.825 20.655 141.995 20.825 ;
      RECT 141.825 23.375 141.995 23.545 ;
      RECT 141.825 26.095 141.995 26.265 ;
      RECT 141.825 28.815 141.995 28.985 ;
      RECT 141.825 31.535 141.995 31.705 ;
      RECT 141.825 34.255 141.995 34.425 ;
      RECT 141.825 36.975 141.995 37.145 ;
      RECT 141.825 39.695 141.995 39.865 ;
      RECT 141.825 42.415 141.995 42.585 ;
      RECT 141.825 45.135 141.995 45.305 ;
      RECT 141.825 47.855 141.995 48.025 ;
      RECT 141.825 50.575 141.995 50.745 ;
      RECT 141.825 53.295 141.995 53.465 ;
      RECT 141.825 56.015 141.995 56.185 ;
      RECT 141.825 58.735 141.995 58.905 ;
      RECT 141.595 24.565 141.765 24.735 ;
      RECT 141.365 9.775 141.535 9.945 ;
      RECT 141.365 12.495 141.535 12.665 ;
      RECT 141.365 15.215 141.535 15.385 ;
      RECT 141.365 17.935 141.535 18.105 ;
      RECT 141.365 20.655 141.535 20.825 ;
      RECT 141.365 23.375 141.535 23.545 ;
      RECT 141.365 26.095 141.535 26.265 ;
      RECT 141.365 28.815 141.535 28.985 ;
      RECT 141.365 31.535 141.535 31.705 ;
      RECT 141.365 34.255 141.535 34.425 ;
      RECT 141.365 36.975 141.535 37.145 ;
      RECT 141.365 39.695 141.535 39.865 ;
      RECT 141.365 42.415 141.535 42.585 ;
      RECT 141.365 45.135 141.535 45.305 ;
      RECT 141.365 47.855 141.535 48.025 ;
      RECT 141.365 50.575 141.535 50.745 ;
      RECT 141.365 53.295 141.535 53.465 ;
      RECT 141.365 56.015 141.535 56.185 ;
      RECT 141.365 58.735 141.535 58.905 ;
      RECT 141.19 26.945 141.36 27.115 ;
      RECT 140.905 9.775 141.075 9.945 ;
      RECT 140.905 12.495 141.075 12.665 ;
      RECT 140.905 15.215 141.075 15.385 ;
      RECT 140.905 17.935 141.075 18.105 ;
      RECT 140.905 20.655 141.075 20.825 ;
      RECT 140.905 23.375 141.075 23.545 ;
      RECT 140.905 25.585 141.075 25.755 ;
      RECT 140.905 26.095 141.075 26.265 ;
      RECT 140.905 28.815 141.075 28.985 ;
      RECT 140.905 31.535 141.075 31.705 ;
      RECT 140.905 34.255 141.075 34.425 ;
      RECT 140.905 36.975 141.075 37.145 ;
      RECT 140.905 39.695 141.075 39.865 ;
      RECT 140.905 42.415 141.075 42.585 ;
      RECT 140.905 45.135 141.075 45.305 ;
      RECT 140.905 47.855 141.075 48.025 ;
      RECT 140.905 50.575 141.075 50.745 ;
      RECT 140.905 53.295 141.075 53.465 ;
      RECT 140.905 56.015 141.075 56.185 ;
      RECT 140.905 58.735 141.075 58.905 ;
      RECT 140.675 27.285 140.845 27.455 ;
      RECT 140.445 9.775 140.615 9.945 ;
      RECT 140.445 12.495 140.615 12.665 ;
      RECT 140.445 15.215 140.615 15.385 ;
      RECT 140.445 17.935 140.615 18.105 ;
      RECT 140.445 20.655 140.615 20.825 ;
      RECT 140.445 23.375 140.615 23.545 ;
      RECT 140.445 26.095 140.615 26.265 ;
      RECT 140.445 28.815 140.615 28.985 ;
      RECT 140.445 31.535 140.615 31.705 ;
      RECT 140.445 34.255 140.615 34.425 ;
      RECT 140.445 36.975 140.615 37.145 ;
      RECT 140.445 39.695 140.615 39.865 ;
      RECT 140.445 42.415 140.615 42.585 ;
      RECT 140.445 45.135 140.615 45.305 ;
      RECT 140.445 47.855 140.615 48.025 ;
      RECT 140.445 50.575 140.615 50.745 ;
      RECT 140.445 53.295 140.615 53.465 ;
      RECT 140.445 56.015 140.615 56.185 ;
      RECT 140.445 58.735 140.615 58.905 ;
      RECT 139.985 9.775 140.155 9.945 ;
      RECT 139.985 12.495 140.155 12.665 ;
      RECT 139.985 15.215 140.155 15.385 ;
      RECT 139.985 15.725 140.155 15.895 ;
      RECT 139.985 17.425 140.155 17.595 ;
      RECT 139.985 17.935 140.155 18.105 ;
      RECT 139.985 20.145 140.155 20.315 ;
      RECT 139.985 20.655 140.155 20.825 ;
      RECT 139.985 23.375 140.155 23.545 ;
      RECT 139.985 26.095 140.155 26.265 ;
      RECT 139.985 28.815 140.155 28.985 ;
      RECT 139.985 31.535 140.155 31.705 ;
      RECT 139.985 34.255 140.155 34.425 ;
      RECT 139.985 36.975 140.155 37.145 ;
      RECT 139.985 39.695 140.155 39.865 ;
      RECT 139.985 42.415 140.155 42.585 ;
      RECT 139.985 45.135 140.155 45.305 ;
      RECT 139.985 47.855 140.155 48.025 ;
      RECT 139.985 50.575 140.155 50.745 ;
      RECT 139.985 53.295 140.155 53.465 ;
      RECT 139.985 56.015 140.155 56.185 ;
      RECT 139.985 58.735 140.155 58.905 ;
      RECT 139.91 27.965 140.08 28.135 ;
      RECT 139.525 9.775 139.695 9.945 ;
      RECT 139.525 12.495 139.695 12.665 ;
      RECT 139.525 15.215 139.695 15.385 ;
      RECT 139.525 17.935 139.695 18.105 ;
      RECT 139.525 20.655 139.695 20.825 ;
      RECT 139.525 23.375 139.695 23.545 ;
      RECT 139.525 26.095 139.695 26.265 ;
      RECT 139.525 28.815 139.695 28.985 ;
      RECT 139.525 31.535 139.695 31.705 ;
      RECT 139.525 34.255 139.695 34.425 ;
      RECT 139.525 36.975 139.695 37.145 ;
      RECT 139.525 39.695 139.695 39.865 ;
      RECT 139.525 42.415 139.695 42.585 ;
      RECT 139.525 45.135 139.695 45.305 ;
      RECT 139.525 47.855 139.695 48.025 ;
      RECT 139.525 50.575 139.695 50.745 ;
      RECT 139.525 53.295 139.695 53.465 ;
      RECT 139.525 56.015 139.695 56.185 ;
      RECT 139.525 58.735 139.695 58.905 ;
      RECT 139.485 27.285 139.655 27.455 ;
      RECT 139.09 26.945 139.26 27.115 ;
      RECT 139.065 9.775 139.235 9.945 ;
      RECT 139.065 12.495 139.235 12.665 ;
      RECT 139.065 15.215 139.235 15.385 ;
      RECT 139.065 17.935 139.235 18.105 ;
      RECT 139.065 20.655 139.235 20.825 ;
      RECT 139.065 23.375 139.235 23.545 ;
      RECT 139.065 26.095 139.235 26.265 ;
      RECT 139.065 28.815 139.235 28.985 ;
      RECT 139.065 31.535 139.235 31.705 ;
      RECT 139.065 34.255 139.235 34.425 ;
      RECT 139.065 36.975 139.235 37.145 ;
      RECT 139.065 39.695 139.235 39.865 ;
      RECT 139.065 42.415 139.235 42.585 ;
      RECT 139.065 45.135 139.235 45.305 ;
      RECT 139.065 47.855 139.235 48.025 ;
      RECT 139.065 50.575 139.235 50.745 ;
      RECT 139.065 53.295 139.235 53.465 ;
      RECT 139.065 56.015 139.235 56.185 ;
      RECT 139.065 58.735 139.235 58.905 ;
      RECT 138.605 9.775 138.775 9.945 ;
      RECT 138.605 12.495 138.775 12.665 ;
      RECT 138.605 13.685 138.775 13.855 ;
      RECT 138.605 15.215 138.775 15.385 ;
      RECT 138.605 17.935 138.775 18.105 ;
      RECT 138.605 20.655 138.775 20.825 ;
      RECT 138.605 23.375 138.775 23.545 ;
      RECT 138.605 26.095 138.775 26.265 ;
      RECT 138.605 27.285 138.775 27.455 ;
      RECT 138.605 28.815 138.775 28.985 ;
      RECT 138.605 31.535 138.775 31.705 ;
      RECT 138.605 34.255 138.775 34.425 ;
      RECT 138.605 36.975 138.775 37.145 ;
      RECT 138.605 39.695 138.775 39.865 ;
      RECT 138.605 42.415 138.775 42.585 ;
      RECT 138.605 45.135 138.775 45.305 ;
      RECT 138.605 47.855 138.775 48.025 ;
      RECT 138.605 50.575 138.775 50.745 ;
      RECT 138.605 53.295 138.775 53.465 ;
      RECT 138.605 56.015 138.775 56.185 ;
      RECT 138.605 58.735 138.775 58.905 ;
      RECT 138.145 9.775 138.315 9.945 ;
      RECT 138.145 12.495 138.315 12.665 ;
      RECT 138.145 15.215 138.315 15.385 ;
      RECT 138.145 17.935 138.315 18.105 ;
      RECT 138.145 20.655 138.315 20.825 ;
      RECT 138.145 22.185 138.315 22.355 ;
      RECT 138.145 23.375 138.315 23.545 ;
      RECT 138.145 26.095 138.315 26.265 ;
      RECT 138.145 28.815 138.315 28.985 ;
      RECT 138.145 31.535 138.315 31.705 ;
      RECT 138.145 34.255 138.315 34.425 ;
      RECT 138.145 36.975 138.315 37.145 ;
      RECT 138.145 39.695 138.315 39.865 ;
      RECT 138.145 42.415 138.315 42.585 ;
      RECT 138.145 45.135 138.315 45.305 ;
      RECT 138.145 47.855 138.315 48.025 ;
      RECT 138.145 50.575 138.315 50.745 ;
      RECT 138.145 53.295 138.315 53.465 ;
      RECT 138.145 56.015 138.315 56.185 ;
      RECT 138.145 58.735 138.315 58.905 ;
      RECT 137.685 9.775 137.855 9.945 ;
      RECT 137.685 12.495 137.855 12.665 ;
      RECT 137.685 15.215 137.855 15.385 ;
      RECT 137.685 17.935 137.855 18.105 ;
      RECT 137.685 20.655 137.855 20.825 ;
      RECT 137.685 23.375 137.855 23.545 ;
      RECT 137.685 24.565 137.855 24.735 ;
      RECT 137.685 26.095 137.855 26.265 ;
      RECT 137.685 28.815 137.855 28.985 ;
      RECT 137.685 31.535 137.855 31.705 ;
      RECT 137.685 34.255 137.855 34.425 ;
      RECT 137.685 36.975 137.855 37.145 ;
      RECT 137.685 39.695 137.855 39.865 ;
      RECT 137.685 42.415 137.855 42.585 ;
      RECT 137.685 45.135 137.855 45.305 ;
      RECT 137.685 47.855 137.855 48.025 ;
      RECT 137.685 50.575 137.855 50.745 ;
      RECT 137.685 53.295 137.855 53.465 ;
      RECT 137.685 56.015 137.855 56.185 ;
      RECT 137.685 58.735 137.855 58.905 ;
      RECT 137.675 16.405 137.845 16.575 ;
      RECT 137.675 19.465 137.845 19.635 ;
      RECT 137.455 22.185 137.625 22.355 ;
      RECT 137.24 16.065 137.41 16.235 ;
      RECT 137.24 19.805 137.41 19.975 ;
      RECT 137.225 9.775 137.395 9.945 ;
      RECT 137.225 12.495 137.395 12.665 ;
      RECT 137.225 15.215 137.395 15.385 ;
      RECT 137.225 17.935 137.395 18.105 ;
      RECT 137.225 20.655 137.395 20.825 ;
      RECT 137.225 23.375 137.395 23.545 ;
      RECT 137.225 26.095 137.395 26.265 ;
      RECT 137.225 28.815 137.395 28.985 ;
      RECT 137.225 31.535 137.395 31.705 ;
      RECT 137.225 34.255 137.395 34.425 ;
      RECT 137.225 36.975 137.395 37.145 ;
      RECT 137.225 39.695 137.395 39.865 ;
      RECT 137.225 42.415 137.395 42.585 ;
      RECT 137.225 45.135 137.395 45.305 ;
      RECT 137.225 47.855 137.395 48.025 ;
      RECT 137.225 50.575 137.395 50.745 ;
      RECT 137.225 53.295 137.395 53.465 ;
      RECT 137.225 56.015 137.395 56.185 ;
      RECT 137.225 58.735 137.395 58.905 ;
      RECT 136.995 24.565 137.165 24.735 ;
      RECT 136.765 9.775 136.935 9.945 ;
      RECT 136.765 12.495 136.935 12.665 ;
      RECT 136.765 15.215 136.935 15.385 ;
      RECT 136.765 17.935 136.935 18.105 ;
      RECT 136.765 20.655 136.935 20.825 ;
      RECT 136.765 22.525 136.935 22.695 ;
      RECT 136.765 23.375 136.935 23.545 ;
      RECT 136.765 26.095 136.935 26.265 ;
      RECT 136.765 28.815 136.935 28.985 ;
      RECT 136.765 31.535 136.935 31.705 ;
      RECT 136.765 34.255 136.935 34.425 ;
      RECT 136.765 36.975 136.935 37.145 ;
      RECT 136.765 39.695 136.935 39.865 ;
      RECT 136.765 42.415 136.935 42.585 ;
      RECT 136.765 45.135 136.935 45.305 ;
      RECT 136.765 47.855 136.935 48.025 ;
      RECT 136.765 50.575 136.935 50.745 ;
      RECT 136.765 53.295 136.935 53.465 ;
      RECT 136.765 56.015 136.935 56.185 ;
      RECT 136.765 58.735 136.935 58.905 ;
      RECT 136.305 9.775 136.475 9.945 ;
      RECT 136.305 12.495 136.475 12.665 ;
      RECT 136.305 15.215 136.475 15.385 ;
      RECT 136.305 17.935 136.475 18.105 ;
      RECT 136.305 20.655 136.475 20.825 ;
      RECT 136.305 22.185 136.475 22.355 ;
      RECT 136.305 23.375 136.475 23.545 ;
      RECT 136.305 24.565 136.475 24.735 ;
      RECT 136.305 26.095 136.475 26.265 ;
      RECT 136.305 28.815 136.475 28.985 ;
      RECT 136.305 31.535 136.475 31.705 ;
      RECT 136.305 34.255 136.475 34.425 ;
      RECT 136.305 36.975 136.475 37.145 ;
      RECT 136.305 39.695 136.475 39.865 ;
      RECT 136.305 42.415 136.475 42.585 ;
      RECT 136.305 45.135 136.475 45.305 ;
      RECT 136.305 47.855 136.475 48.025 ;
      RECT 136.305 50.575 136.475 50.745 ;
      RECT 136.305 53.295 136.475 53.465 ;
      RECT 136.305 56.015 136.475 56.185 ;
      RECT 136.305 58.735 136.475 58.905 ;
      RECT 135.845 9.775 136.015 9.945 ;
      RECT 135.845 12.495 136.015 12.665 ;
      RECT 135.845 15.215 136.015 15.385 ;
      RECT 135.845 17.935 136.015 18.105 ;
      RECT 135.845 20.655 136.015 20.825 ;
      RECT 135.845 23.375 136.015 23.545 ;
      RECT 135.845 24.565 136.015 24.735 ;
      RECT 135.845 26.095 136.015 26.265 ;
      RECT 135.845 28.815 136.015 28.985 ;
      RECT 135.845 31.535 136.015 31.705 ;
      RECT 135.845 34.255 136.015 34.425 ;
      RECT 135.845 36.975 136.015 37.145 ;
      RECT 135.845 39.695 136.015 39.865 ;
      RECT 135.845 42.415 136.015 42.585 ;
      RECT 135.845 45.135 136.015 45.305 ;
      RECT 135.845 47.855 136.015 48.025 ;
      RECT 135.845 50.575 136.015 50.745 ;
      RECT 135.845 53.295 136.015 53.465 ;
      RECT 135.845 56.015 136.015 56.185 ;
      RECT 135.845 58.735 136.015 58.905 ;
      RECT 135.67 16.065 135.84 16.235 ;
      RECT 135.67 19.805 135.84 19.975 ;
      RECT 135.615 22.185 135.785 22.355 ;
      RECT 135.385 9.775 135.555 9.945 ;
      RECT 135.385 12.495 135.555 12.665 ;
      RECT 135.385 15.215 135.555 15.385 ;
      RECT 135.385 17.935 135.555 18.105 ;
      RECT 135.385 20.655 135.555 20.825 ;
      RECT 135.385 23.375 135.555 23.545 ;
      RECT 135.385 26.095 135.555 26.265 ;
      RECT 135.385 28.815 135.555 28.985 ;
      RECT 135.385 31.535 135.555 31.705 ;
      RECT 135.385 34.255 135.555 34.425 ;
      RECT 135.385 36.975 135.555 37.145 ;
      RECT 135.385 39.695 135.555 39.865 ;
      RECT 135.385 42.415 135.555 42.585 ;
      RECT 135.385 45.135 135.555 45.305 ;
      RECT 135.385 47.855 135.555 48.025 ;
      RECT 135.385 50.575 135.555 50.745 ;
      RECT 135.385 53.295 135.555 53.465 ;
      RECT 135.385 56.015 135.555 56.185 ;
      RECT 135.385 58.735 135.555 58.905 ;
      RECT 135.155 16.405 135.325 16.575 ;
      RECT 135.155 19.465 135.325 19.635 ;
      RECT 135.155 24.565 135.325 24.735 ;
      RECT 134.925 9.775 135.095 9.945 ;
      RECT 134.925 12.495 135.095 12.665 ;
      RECT 134.925 15.215 135.095 15.385 ;
      RECT 134.925 17.935 135.095 18.105 ;
      RECT 134.925 20.655 135.095 20.825 ;
      RECT 134.925 21.505 135.095 21.675 ;
      RECT 134.925 23.375 135.095 23.545 ;
      RECT 134.925 26.095 135.095 26.265 ;
      RECT 134.925 28.815 135.095 28.985 ;
      RECT 134.925 31.535 135.095 31.705 ;
      RECT 134.925 34.255 135.095 34.425 ;
      RECT 134.925 36.975 135.095 37.145 ;
      RECT 134.925 39.695 135.095 39.865 ;
      RECT 134.925 42.415 135.095 42.585 ;
      RECT 134.925 45.135 135.095 45.305 ;
      RECT 134.925 47.855 135.095 48.025 ;
      RECT 134.925 50.575 135.095 50.745 ;
      RECT 134.925 53.295 135.095 53.465 ;
      RECT 134.925 56.015 135.095 56.185 ;
      RECT 134.925 58.735 135.095 58.905 ;
      RECT 134.465 9.775 134.635 9.945 ;
      RECT 134.465 12.495 134.635 12.665 ;
      RECT 134.465 15.215 134.635 15.385 ;
      RECT 134.465 17.935 134.635 18.105 ;
      RECT 134.465 20.655 134.635 20.825 ;
      RECT 134.465 23.375 134.635 23.545 ;
      RECT 134.465 23.885 134.635 24.055 ;
      RECT 134.465 26.095 134.635 26.265 ;
      RECT 134.465 28.815 134.635 28.985 ;
      RECT 134.465 31.535 134.635 31.705 ;
      RECT 134.465 34.255 134.635 34.425 ;
      RECT 134.465 36.975 134.635 37.145 ;
      RECT 134.465 39.695 134.635 39.865 ;
      RECT 134.465 42.415 134.635 42.585 ;
      RECT 134.465 45.135 134.635 45.305 ;
      RECT 134.465 47.855 134.635 48.025 ;
      RECT 134.465 50.575 134.635 50.745 ;
      RECT 134.465 53.295 134.635 53.465 ;
      RECT 134.465 56.015 134.635 56.185 ;
      RECT 134.465 58.735 134.635 58.905 ;
      RECT 134.39 16.745 134.56 16.915 ;
      RECT 134.39 18.785 134.56 18.955 ;
      RECT 134.005 9.775 134.175 9.945 ;
      RECT 134.005 12.495 134.175 12.665 ;
      RECT 134.005 15.215 134.175 15.385 ;
      RECT 134.005 17.935 134.175 18.105 ;
      RECT 134.005 20.655 134.175 20.825 ;
      RECT 134.005 23.375 134.175 23.545 ;
      RECT 134.005 26.095 134.175 26.265 ;
      RECT 134.005 28.815 134.175 28.985 ;
      RECT 134.005 31.535 134.175 31.705 ;
      RECT 134.005 34.255 134.175 34.425 ;
      RECT 134.005 36.975 134.175 37.145 ;
      RECT 134.005 39.695 134.175 39.865 ;
      RECT 134.005 42.415 134.175 42.585 ;
      RECT 134.005 45.135 134.175 45.305 ;
      RECT 134.005 47.855 134.175 48.025 ;
      RECT 134.005 50.575 134.175 50.745 ;
      RECT 134.005 53.295 134.175 53.465 ;
      RECT 134.005 56.015 134.175 56.185 ;
      RECT 134.005 58.735 134.175 58.905 ;
      RECT 133.965 16.405 134.135 16.575 ;
      RECT 133.965 19.465 134.135 19.635 ;
      RECT 133.57 16.065 133.74 16.235 ;
      RECT 133.57 19.805 133.74 19.975 ;
      RECT 133.545 9.775 133.715 9.945 ;
      RECT 133.545 12.495 133.715 12.665 ;
      RECT 133.545 15.215 133.715 15.385 ;
      RECT 133.545 17.935 133.715 18.105 ;
      RECT 133.545 20.655 133.715 20.825 ;
      RECT 133.545 23.375 133.715 23.545 ;
      RECT 133.545 26.095 133.715 26.265 ;
      RECT 133.545 28.815 133.715 28.985 ;
      RECT 133.545 31.535 133.715 31.705 ;
      RECT 133.545 34.255 133.715 34.425 ;
      RECT 133.545 36.975 133.715 37.145 ;
      RECT 133.545 39.695 133.715 39.865 ;
      RECT 133.545 42.415 133.715 42.585 ;
      RECT 133.545 45.135 133.715 45.305 ;
      RECT 133.545 47.855 133.715 48.025 ;
      RECT 133.545 50.575 133.715 50.745 ;
      RECT 133.545 53.295 133.715 53.465 ;
      RECT 133.545 56.015 133.715 56.185 ;
      RECT 133.545 58.735 133.715 58.905 ;
      RECT 133.085 9.775 133.255 9.945 ;
      RECT 133.085 11.305 133.255 11.475 ;
      RECT 133.085 12.495 133.255 12.665 ;
      RECT 133.085 15.215 133.255 15.385 ;
      RECT 133.085 16.745 133.255 16.915 ;
      RECT 133.085 17.935 133.255 18.105 ;
      RECT 133.085 19.125 133.255 19.295 ;
      RECT 133.085 20.655 133.255 20.825 ;
      RECT 133.085 23.375 133.255 23.545 ;
      RECT 133.085 26.095 133.255 26.265 ;
      RECT 133.085 28.815 133.255 28.985 ;
      RECT 133.085 31.535 133.255 31.705 ;
      RECT 133.085 34.255 133.255 34.425 ;
      RECT 133.085 36.975 133.255 37.145 ;
      RECT 133.085 39.695 133.255 39.865 ;
      RECT 133.085 42.415 133.255 42.585 ;
      RECT 133.085 45.135 133.255 45.305 ;
      RECT 133.085 47.855 133.255 48.025 ;
      RECT 133.085 50.575 133.255 50.745 ;
      RECT 133.085 53.295 133.255 53.465 ;
      RECT 133.085 56.015 133.255 56.185 ;
      RECT 133.085 58.735 133.255 58.905 ;
      RECT 132.625 9.775 132.795 9.945 ;
      RECT 132.625 12.495 132.795 12.665 ;
      RECT 132.625 15.215 132.795 15.385 ;
      RECT 132.625 17.935 132.795 18.105 ;
      RECT 132.625 20.655 132.795 20.825 ;
      RECT 132.625 23.375 132.795 23.545 ;
      RECT 132.625 26.095 132.795 26.265 ;
      RECT 132.625 28.815 132.795 28.985 ;
      RECT 132.625 31.535 132.795 31.705 ;
      RECT 132.625 34.255 132.795 34.425 ;
      RECT 132.625 36.975 132.795 37.145 ;
      RECT 132.625 39.695 132.795 39.865 ;
      RECT 132.625 42.415 132.795 42.585 ;
      RECT 132.625 45.135 132.795 45.305 ;
      RECT 132.625 47.855 132.795 48.025 ;
      RECT 132.625 50.575 132.795 50.745 ;
      RECT 132.625 53.295 132.795 53.465 ;
      RECT 132.625 56.015 132.795 56.185 ;
      RECT 132.625 58.735 132.795 58.905 ;
      RECT 132.165 9.775 132.335 9.945 ;
      RECT 132.165 12.495 132.335 12.665 ;
      RECT 132.165 15.215 132.335 15.385 ;
      RECT 132.165 17.935 132.335 18.105 ;
      RECT 132.165 20.655 132.335 20.825 ;
      RECT 132.165 21.165 132.335 21.335 ;
      RECT 132.165 22.865 132.335 23.035 ;
      RECT 132.165 23.375 132.335 23.545 ;
      RECT 132.165 26.095 132.335 26.265 ;
      RECT 132.165 28.815 132.335 28.985 ;
      RECT 132.165 31.535 132.335 31.705 ;
      RECT 132.165 34.255 132.335 34.425 ;
      RECT 132.165 36.975 132.335 37.145 ;
      RECT 132.165 39.695 132.335 39.865 ;
      RECT 132.165 42.415 132.335 42.585 ;
      RECT 132.165 45.135 132.335 45.305 ;
      RECT 132.165 47.855 132.335 48.025 ;
      RECT 132.165 50.575 132.335 50.745 ;
      RECT 132.165 53.295 132.335 53.465 ;
      RECT 132.165 56.015 132.335 56.185 ;
      RECT 132.165 58.735 132.335 58.905 ;
      RECT 131.705 9.775 131.875 9.945 ;
      RECT 131.705 12.495 131.875 12.665 ;
      RECT 131.705 15.215 131.875 15.385 ;
      RECT 131.705 17.935 131.875 18.105 ;
      RECT 131.705 20.655 131.875 20.825 ;
      RECT 131.705 22.865 131.875 23.035 ;
      RECT 131.705 23.375 131.875 23.545 ;
      RECT 131.705 26.095 131.875 26.265 ;
      RECT 131.705 28.815 131.875 28.985 ;
      RECT 131.705 31.535 131.875 31.705 ;
      RECT 131.705 34.255 131.875 34.425 ;
      RECT 131.705 36.975 131.875 37.145 ;
      RECT 131.705 39.695 131.875 39.865 ;
      RECT 131.705 42.415 131.875 42.585 ;
      RECT 131.705 45.135 131.875 45.305 ;
      RECT 131.705 47.855 131.875 48.025 ;
      RECT 131.705 50.575 131.875 50.745 ;
      RECT 131.705 53.295 131.875 53.465 ;
      RECT 131.705 56.015 131.875 56.185 ;
      RECT 131.705 58.735 131.875 58.905 ;
      RECT 131.245 9.775 131.415 9.945 ;
      RECT 131.245 12.495 131.415 12.665 ;
      RECT 131.245 15.215 131.415 15.385 ;
      RECT 131.245 17.935 131.415 18.105 ;
      RECT 131.245 20.655 131.415 20.825 ;
      RECT 131.245 23.375 131.415 23.545 ;
      RECT 131.245 26.095 131.415 26.265 ;
      RECT 131.245 28.815 131.415 28.985 ;
      RECT 131.245 31.535 131.415 31.705 ;
      RECT 131.245 34.255 131.415 34.425 ;
      RECT 131.245 34.765 131.415 34.935 ;
      RECT 131.245 36.975 131.415 37.145 ;
      RECT 131.245 39.695 131.415 39.865 ;
      RECT 131.245 42.415 131.415 42.585 ;
      RECT 131.245 45.135 131.415 45.305 ;
      RECT 131.245 47.855 131.415 48.025 ;
      RECT 131.245 50.575 131.415 50.745 ;
      RECT 131.245 53.295 131.415 53.465 ;
      RECT 131.245 56.015 131.415 56.185 ;
      RECT 131.245 58.735 131.415 58.905 ;
      RECT 131.015 22.185 131.185 22.355 ;
      RECT 130.785 9.775 130.955 9.945 ;
      RECT 130.785 12.495 130.955 12.665 ;
      RECT 130.785 15.215 130.955 15.385 ;
      RECT 130.785 17.935 130.955 18.105 ;
      RECT 130.785 20.655 130.955 20.825 ;
      RECT 130.785 23.375 130.955 23.545 ;
      RECT 130.785 26.095 130.955 26.265 ;
      RECT 130.785 28.815 130.955 28.985 ;
      RECT 130.785 31.535 130.955 31.705 ;
      RECT 130.785 34.255 130.955 34.425 ;
      RECT 130.785 36.975 130.955 37.145 ;
      RECT 130.785 39.695 130.955 39.865 ;
      RECT 130.785 42.415 130.955 42.585 ;
      RECT 130.785 45.135 130.955 45.305 ;
      RECT 130.785 47.855 130.955 48.025 ;
      RECT 130.785 50.575 130.955 50.745 ;
      RECT 130.785 53.295 130.955 53.465 ;
      RECT 130.785 56.015 130.955 56.185 ;
      RECT 130.785 58.735 130.955 58.905 ;
      RECT 130.325 9.775 130.495 9.945 ;
      RECT 130.325 12.495 130.495 12.665 ;
      RECT 130.325 15.215 130.495 15.385 ;
      RECT 130.325 17.935 130.495 18.105 ;
      RECT 130.325 20.655 130.495 20.825 ;
      RECT 130.325 22.185 130.495 22.355 ;
      RECT 130.325 23.375 130.495 23.545 ;
      RECT 130.325 26.095 130.495 26.265 ;
      RECT 130.325 27.625 130.495 27.795 ;
      RECT 130.325 28.815 130.495 28.985 ;
      RECT 130.325 31.535 130.495 31.705 ;
      RECT 130.325 34.255 130.495 34.425 ;
      RECT 130.325 36.975 130.495 37.145 ;
      RECT 130.325 39.695 130.495 39.865 ;
      RECT 130.325 42.415 130.495 42.585 ;
      RECT 130.325 45.135 130.495 45.305 ;
      RECT 130.325 47.855 130.495 48.025 ;
      RECT 130.325 50.575 130.495 50.745 ;
      RECT 130.325 53.295 130.495 53.465 ;
      RECT 130.325 56.015 130.495 56.185 ;
      RECT 130.325 58.735 130.495 58.905 ;
      RECT 129.865 9.775 130.035 9.945 ;
      RECT 129.865 12.495 130.035 12.665 ;
      RECT 129.865 15.215 130.035 15.385 ;
      RECT 129.865 17.935 130.035 18.105 ;
      RECT 129.865 20.655 130.035 20.825 ;
      RECT 129.865 22.525 130.035 22.695 ;
      RECT 129.865 23.375 130.035 23.545 ;
      RECT 129.865 26.095 130.035 26.265 ;
      RECT 129.865 28.815 130.035 28.985 ;
      RECT 129.865 31.535 130.035 31.705 ;
      RECT 129.865 34.255 130.035 34.425 ;
      RECT 129.865 36.975 130.035 37.145 ;
      RECT 129.865 39.695 130.035 39.865 ;
      RECT 129.865 42.415 130.035 42.585 ;
      RECT 129.865 45.135 130.035 45.305 ;
      RECT 129.865 47.855 130.035 48.025 ;
      RECT 129.865 50.575 130.035 50.745 ;
      RECT 129.865 53.295 130.035 53.465 ;
      RECT 129.865 56.015 130.035 56.185 ;
      RECT 129.865 58.735 130.035 58.905 ;
      RECT 129.635 27.625 129.805 27.795 ;
      RECT 129.405 9.775 129.575 9.945 ;
      RECT 129.405 12.495 129.575 12.665 ;
      RECT 129.405 15.215 129.575 15.385 ;
      RECT 129.405 17.935 129.575 18.105 ;
      RECT 129.405 20.655 129.575 20.825 ;
      RECT 129.405 23.375 129.575 23.545 ;
      RECT 129.405 26.095 129.575 26.265 ;
      RECT 129.405 28.815 129.575 28.985 ;
      RECT 129.405 31.535 129.575 31.705 ;
      RECT 129.405 34.255 129.575 34.425 ;
      RECT 129.405 36.975 129.575 37.145 ;
      RECT 129.405 39.695 129.575 39.865 ;
      RECT 129.405 42.415 129.575 42.585 ;
      RECT 129.405 45.135 129.575 45.305 ;
      RECT 129.405 47.855 129.575 48.025 ;
      RECT 129.405 50.575 129.575 50.745 ;
      RECT 129.405 53.295 129.575 53.465 ;
      RECT 129.405 56.015 129.575 56.185 ;
      RECT 129.405 58.735 129.575 58.905 ;
      RECT 129.175 22.185 129.345 22.355 ;
      RECT 128.945 9.775 129.115 9.945 ;
      RECT 128.945 12.495 129.115 12.665 ;
      RECT 128.945 15.215 129.115 15.385 ;
      RECT 128.945 17.935 129.115 18.105 ;
      RECT 128.945 20.655 129.115 20.825 ;
      RECT 128.945 23.375 129.115 23.545 ;
      RECT 128.945 26.095 129.115 26.265 ;
      RECT 128.945 27.965 129.115 28.135 ;
      RECT 128.945 28.815 129.115 28.985 ;
      RECT 128.945 31.535 129.115 31.705 ;
      RECT 128.945 34.255 129.115 34.425 ;
      RECT 128.945 36.975 129.115 37.145 ;
      RECT 128.945 39.695 129.115 39.865 ;
      RECT 128.945 42.415 129.115 42.585 ;
      RECT 128.945 45.135 129.115 45.305 ;
      RECT 128.945 47.855 129.115 48.025 ;
      RECT 128.945 50.575 129.115 50.745 ;
      RECT 128.945 53.295 129.115 53.465 ;
      RECT 128.945 56.015 129.115 56.185 ;
      RECT 128.945 58.735 129.115 58.905 ;
      RECT 128.935 35.785 129.105 35.955 ;
      RECT 128.5 36.125 128.67 36.295 ;
      RECT 128.485 9.775 128.655 9.945 ;
      RECT 128.485 12.495 128.655 12.665 ;
      RECT 128.485 15.215 128.655 15.385 ;
      RECT 128.485 17.935 128.655 18.105 ;
      RECT 128.485 20.655 128.655 20.825 ;
      RECT 128.485 22.185 128.655 22.355 ;
      RECT 128.485 23.375 128.655 23.545 ;
      RECT 128.485 26.095 128.655 26.265 ;
      RECT 128.485 27.625 128.655 27.795 ;
      RECT 128.485 28.815 128.655 28.985 ;
      RECT 128.485 31.535 128.655 31.705 ;
      RECT 128.485 34.255 128.655 34.425 ;
      RECT 128.485 36.975 128.655 37.145 ;
      RECT 128.485 39.695 128.655 39.865 ;
      RECT 128.485 42.415 128.655 42.585 ;
      RECT 128.485 45.135 128.655 45.305 ;
      RECT 128.485 47.855 128.655 48.025 ;
      RECT 128.485 50.575 128.655 50.745 ;
      RECT 128.485 53.295 128.655 53.465 ;
      RECT 128.485 56.015 128.655 56.185 ;
      RECT 128.485 58.735 128.655 58.905 ;
      RECT 128.025 9.775 128.195 9.945 ;
      RECT 128.025 12.495 128.195 12.665 ;
      RECT 128.025 15.215 128.195 15.385 ;
      RECT 128.025 17.935 128.195 18.105 ;
      RECT 128.025 20.655 128.195 20.825 ;
      RECT 128.025 21.165 128.195 21.335 ;
      RECT 128.025 23.375 128.195 23.545 ;
      RECT 128.025 26.095 128.195 26.265 ;
      RECT 128.025 28.815 128.195 28.985 ;
      RECT 128.025 31.535 128.195 31.705 ;
      RECT 128.025 34.255 128.195 34.425 ;
      RECT 128.025 36.975 128.195 37.145 ;
      RECT 128.025 39.695 128.195 39.865 ;
      RECT 128.025 42.415 128.195 42.585 ;
      RECT 128.025 45.135 128.195 45.305 ;
      RECT 128.025 47.855 128.195 48.025 ;
      RECT 128.025 50.575 128.195 50.745 ;
      RECT 128.025 53.295 128.195 53.465 ;
      RECT 128.025 56.015 128.195 56.185 ;
      RECT 128.025 58.735 128.195 58.905 ;
      RECT 127.795 27.625 127.965 27.795 ;
      RECT 127.565 9.775 127.735 9.945 ;
      RECT 127.565 12.495 127.735 12.665 ;
      RECT 127.565 15.215 127.735 15.385 ;
      RECT 127.565 17.935 127.735 18.105 ;
      RECT 127.565 20.655 127.735 20.825 ;
      RECT 127.565 23.375 127.735 23.545 ;
      RECT 127.565 26.095 127.735 26.265 ;
      RECT 127.565 28.815 127.735 28.985 ;
      RECT 127.565 31.535 127.735 31.705 ;
      RECT 127.565 34.255 127.735 34.425 ;
      RECT 127.565 36.975 127.735 37.145 ;
      RECT 127.565 39.695 127.735 39.865 ;
      RECT 127.565 42.415 127.735 42.585 ;
      RECT 127.565 45.135 127.735 45.305 ;
      RECT 127.565 47.855 127.735 48.025 ;
      RECT 127.565 50.575 127.735 50.745 ;
      RECT 127.565 53.295 127.735 53.465 ;
      RECT 127.565 56.015 127.735 56.185 ;
      RECT 127.565 58.735 127.735 58.905 ;
      RECT 127.105 9.775 127.275 9.945 ;
      RECT 127.105 12.495 127.275 12.665 ;
      RECT 127.105 15.215 127.275 15.385 ;
      RECT 127.105 17.935 127.275 18.105 ;
      RECT 127.105 20.655 127.275 20.825 ;
      RECT 127.105 23.375 127.275 23.545 ;
      RECT 127.105 26.095 127.275 26.265 ;
      RECT 127.105 28.305 127.275 28.475 ;
      RECT 127.105 28.815 127.275 28.985 ;
      RECT 127.105 31.535 127.275 31.705 ;
      RECT 127.105 34.255 127.275 34.425 ;
      RECT 127.105 36.975 127.275 37.145 ;
      RECT 127.105 39.695 127.275 39.865 ;
      RECT 127.105 42.415 127.275 42.585 ;
      RECT 127.105 45.135 127.275 45.305 ;
      RECT 127.105 47.855 127.275 48.025 ;
      RECT 127.105 50.575 127.275 50.745 ;
      RECT 127.105 53.295 127.275 53.465 ;
      RECT 127.105 56.015 127.275 56.185 ;
      RECT 127.105 58.735 127.275 58.905 ;
      RECT 126.93 36.125 127.1 36.295 ;
      RECT 126.645 9.775 126.815 9.945 ;
      RECT 126.645 12.495 126.815 12.665 ;
      RECT 126.645 15.215 126.815 15.385 ;
      RECT 126.645 17.935 126.815 18.105 ;
      RECT 126.645 20.655 126.815 20.825 ;
      RECT 126.645 23.375 126.815 23.545 ;
      RECT 126.645 26.095 126.815 26.265 ;
      RECT 126.645 28.815 126.815 28.985 ;
      RECT 126.645 31.535 126.815 31.705 ;
      RECT 126.645 34.255 126.815 34.425 ;
      RECT 126.645 36.975 126.815 37.145 ;
      RECT 126.645 39.695 126.815 39.865 ;
      RECT 126.645 42.415 126.815 42.585 ;
      RECT 126.645 45.135 126.815 45.305 ;
      RECT 126.645 47.855 126.815 48.025 ;
      RECT 126.645 50.575 126.815 50.745 ;
      RECT 126.645 53.295 126.815 53.465 ;
      RECT 126.645 56.015 126.815 56.185 ;
      RECT 126.645 58.735 126.815 58.905 ;
      RECT 126.415 35.785 126.585 35.955 ;
      RECT 126.185 9.775 126.355 9.945 ;
      RECT 126.185 12.495 126.355 12.665 ;
      RECT 126.185 15.215 126.355 15.385 ;
      RECT 126.185 17.935 126.355 18.105 ;
      RECT 126.185 20.655 126.355 20.825 ;
      RECT 126.185 23.375 126.355 23.545 ;
      RECT 126.185 26.095 126.355 26.265 ;
      RECT 126.185 28.815 126.355 28.985 ;
      RECT 126.185 31.535 126.355 31.705 ;
      RECT 126.185 34.255 126.355 34.425 ;
      RECT 126.185 36.975 126.355 37.145 ;
      RECT 126.185 39.695 126.355 39.865 ;
      RECT 126.185 42.415 126.355 42.585 ;
      RECT 126.185 45.135 126.355 45.305 ;
      RECT 126.185 47.855 126.355 48.025 ;
      RECT 126.185 50.575 126.355 50.745 ;
      RECT 126.185 53.295 126.355 53.465 ;
      RECT 126.185 56.015 126.355 56.185 ;
      RECT 126.185 58.735 126.355 58.905 ;
      RECT 125.725 9.775 125.895 9.945 ;
      RECT 125.725 12.495 125.895 12.665 ;
      RECT 125.725 15.215 125.895 15.385 ;
      RECT 125.725 17.935 125.895 18.105 ;
      RECT 125.725 20.655 125.895 20.825 ;
      RECT 125.725 23.375 125.895 23.545 ;
      RECT 125.725 26.095 125.895 26.265 ;
      RECT 125.725 28.815 125.895 28.985 ;
      RECT 125.725 31.535 125.895 31.705 ;
      RECT 125.725 34.255 125.895 34.425 ;
      RECT 125.725 36.975 125.895 37.145 ;
      RECT 125.725 39.695 125.895 39.865 ;
      RECT 125.725 42.415 125.895 42.585 ;
      RECT 125.725 45.135 125.895 45.305 ;
      RECT 125.725 47.855 125.895 48.025 ;
      RECT 125.725 50.575 125.895 50.745 ;
      RECT 125.725 53.295 125.895 53.465 ;
      RECT 125.725 56.015 125.895 56.185 ;
      RECT 125.725 58.735 125.895 58.905 ;
      RECT 125.715 21.845 125.885 22.015 ;
      RECT 125.65 35.105 125.82 35.275 ;
      RECT 125.28 21.505 125.45 21.675 ;
      RECT 125.265 9.775 125.435 9.945 ;
      RECT 125.265 12.495 125.435 12.665 ;
      RECT 125.265 15.215 125.435 15.385 ;
      RECT 125.265 15.725 125.435 15.895 ;
      RECT 125.265 17.425 125.435 17.595 ;
      RECT 125.265 17.935 125.435 18.105 ;
      RECT 125.265 20.655 125.435 20.825 ;
      RECT 125.265 23.375 125.435 23.545 ;
      RECT 125.265 26.095 125.435 26.265 ;
      RECT 125.265 28.815 125.435 28.985 ;
      RECT 125.265 31.535 125.435 31.705 ;
      RECT 125.265 34.255 125.435 34.425 ;
      RECT 125.265 36.975 125.435 37.145 ;
      RECT 125.265 39.695 125.435 39.865 ;
      RECT 125.265 42.415 125.435 42.585 ;
      RECT 125.265 45.135 125.435 45.305 ;
      RECT 125.265 47.855 125.435 48.025 ;
      RECT 125.265 50.575 125.435 50.745 ;
      RECT 125.265 53.295 125.435 53.465 ;
      RECT 125.265 56.015 125.435 56.185 ;
      RECT 125.265 58.735 125.435 58.905 ;
      RECT 125.225 35.785 125.395 35.955 ;
      RECT 124.83 36.125 125 36.295 ;
      RECT 124.805 9.775 124.975 9.945 ;
      RECT 124.805 11.305 124.975 11.475 ;
      RECT 124.805 12.495 124.975 12.665 ;
      RECT 124.805 15.215 124.975 15.385 ;
      RECT 124.805 17.935 124.975 18.105 ;
      RECT 124.805 19.125 124.975 19.295 ;
      RECT 124.805 20.145 124.975 20.315 ;
      RECT 124.805 20.655 124.975 20.825 ;
      RECT 124.805 23.375 124.975 23.545 ;
      RECT 124.805 26.095 124.975 26.265 ;
      RECT 124.805 28.815 124.975 28.985 ;
      RECT 124.805 31.535 124.975 31.705 ;
      RECT 124.805 34.255 124.975 34.425 ;
      RECT 124.805 36.975 124.975 37.145 ;
      RECT 124.805 39.695 124.975 39.865 ;
      RECT 124.805 42.415 124.975 42.585 ;
      RECT 124.805 45.135 124.975 45.305 ;
      RECT 124.805 47.855 124.975 48.025 ;
      RECT 124.805 50.575 124.975 50.745 ;
      RECT 124.805 53.295 124.975 53.465 ;
      RECT 124.805 56.015 124.975 56.185 ;
      RECT 124.805 58.735 124.975 58.905 ;
      RECT 124.345 9.775 124.515 9.945 ;
      RECT 124.345 12.495 124.515 12.665 ;
      RECT 124.345 15.215 124.515 15.385 ;
      RECT 124.345 17.935 124.515 18.105 ;
      RECT 124.345 20.655 124.515 20.825 ;
      RECT 124.345 23.375 124.515 23.545 ;
      RECT 124.345 26.095 124.515 26.265 ;
      RECT 124.345 28.815 124.515 28.985 ;
      RECT 124.345 31.535 124.515 31.705 ;
      RECT 124.345 34.255 124.515 34.425 ;
      RECT 124.345 35.445 124.515 35.615 ;
      RECT 124.345 36.975 124.515 37.145 ;
      RECT 124.345 39.695 124.515 39.865 ;
      RECT 124.345 42.415 124.515 42.585 ;
      RECT 124.345 45.135 124.515 45.305 ;
      RECT 124.345 47.855 124.515 48.025 ;
      RECT 124.345 50.575 124.515 50.745 ;
      RECT 124.345 53.295 124.515 53.465 ;
      RECT 124.345 56.015 124.515 56.185 ;
      RECT 124.345 58.735 124.515 58.905 ;
      RECT 123.885 9.775 124.055 9.945 ;
      RECT 123.885 12.495 124.055 12.665 ;
      RECT 123.885 15.215 124.055 15.385 ;
      RECT 123.885 17.935 124.055 18.105 ;
      RECT 123.885 20.655 124.055 20.825 ;
      RECT 123.885 23.375 124.055 23.545 ;
      RECT 123.885 26.095 124.055 26.265 ;
      RECT 123.885 28.815 124.055 28.985 ;
      RECT 123.885 31.535 124.055 31.705 ;
      RECT 123.885 34.255 124.055 34.425 ;
      RECT 123.885 36.975 124.055 37.145 ;
      RECT 123.885 39.695 124.055 39.865 ;
      RECT 123.885 42.415 124.055 42.585 ;
      RECT 123.885 45.135 124.055 45.305 ;
      RECT 123.885 47.855 124.055 48.025 ;
      RECT 123.885 50.575 124.055 50.745 ;
      RECT 123.885 53.295 124.055 53.465 ;
      RECT 123.885 56.015 124.055 56.185 ;
      RECT 123.885 58.735 124.055 58.905 ;
      RECT 123.71 21.505 123.88 21.675 ;
      RECT 123.425 9.775 123.595 9.945 ;
      RECT 123.425 12.495 123.595 12.665 ;
      RECT 123.425 15.215 123.595 15.385 ;
      RECT 123.425 17.935 123.595 18.105 ;
      RECT 123.425 20.655 123.595 20.825 ;
      RECT 123.425 23.375 123.595 23.545 ;
      RECT 123.425 26.095 123.595 26.265 ;
      RECT 123.425 28.815 123.595 28.985 ;
      RECT 123.425 31.535 123.595 31.705 ;
      RECT 123.425 34.255 123.595 34.425 ;
      RECT 123.425 36.975 123.595 37.145 ;
      RECT 123.425 39.695 123.595 39.865 ;
      RECT 123.425 42.415 123.595 42.585 ;
      RECT 123.425 45.135 123.595 45.305 ;
      RECT 123.425 47.855 123.595 48.025 ;
      RECT 123.425 50.575 123.595 50.745 ;
      RECT 123.425 53.295 123.595 53.465 ;
      RECT 123.425 56.015 123.595 56.185 ;
      RECT 123.425 58.735 123.595 58.905 ;
      RECT 123.195 21.845 123.365 22.015 ;
      RECT 122.965 9.775 123.135 9.945 ;
      RECT 122.965 12.495 123.135 12.665 ;
      RECT 122.965 15.215 123.135 15.385 ;
      RECT 122.965 17.935 123.135 18.105 ;
      RECT 122.965 20.655 123.135 20.825 ;
      RECT 122.965 23.375 123.135 23.545 ;
      RECT 122.965 26.095 123.135 26.265 ;
      RECT 122.965 28.815 123.135 28.985 ;
      RECT 122.965 31.535 123.135 31.705 ;
      RECT 122.965 34.255 123.135 34.425 ;
      RECT 122.965 36.975 123.135 37.145 ;
      RECT 122.965 39.695 123.135 39.865 ;
      RECT 122.965 42.415 123.135 42.585 ;
      RECT 122.965 45.135 123.135 45.305 ;
      RECT 122.965 47.855 123.135 48.025 ;
      RECT 122.965 50.575 123.135 50.745 ;
      RECT 122.965 53.295 123.135 53.465 ;
      RECT 122.965 56.015 123.135 56.185 ;
      RECT 122.965 58.735 123.135 58.905 ;
      RECT 122.955 16.405 123.125 16.575 ;
      RECT 122.52 16.065 122.69 16.235 ;
      RECT 122.505 9.775 122.675 9.945 ;
      RECT 122.505 12.495 122.675 12.665 ;
      RECT 122.505 15.215 122.675 15.385 ;
      RECT 122.505 17.935 122.675 18.105 ;
      RECT 122.505 20.655 122.675 20.825 ;
      RECT 122.505 23.375 122.675 23.545 ;
      RECT 122.505 26.095 122.675 26.265 ;
      RECT 122.505 28.815 122.675 28.985 ;
      RECT 122.505 31.535 122.675 31.705 ;
      RECT 122.505 34.255 122.675 34.425 ;
      RECT 122.505 36.975 122.675 37.145 ;
      RECT 122.505 39.695 122.675 39.865 ;
      RECT 122.505 42.415 122.675 42.585 ;
      RECT 122.505 45.135 122.675 45.305 ;
      RECT 122.505 47.855 122.675 48.025 ;
      RECT 122.505 50.575 122.675 50.745 ;
      RECT 122.505 53.295 122.675 53.465 ;
      RECT 122.505 56.015 122.675 56.185 ;
      RECT 122.505 58.735 122.675 58.905 ;
      RECT 122.43 22.525 122.6 22.695 ;
      RECT 122.045 9.775 122.215 9.945 ;
      RECT 122.045 12.495 122.215 12.665 ;
      RECT 122.045 14.705 122.215 14.875 ;
      RECT 122.045 15.215 122.215 15.385 ;
      RECT 122.045 17.935 122.215 18.105 ;
      RECT 122.045 20.655 122.215 20.825 ;
      RECT 122.045 23.375 122.215 23.545 ;
      RECT 122.045 26.095 122.215 26.265 ;
      RECT 122.045 28.815 122.215 28.985 ;
      RECT 122.045 31.535 122.215 31.705 ;
      RECT 122.045 34.255 122.215 34.425 ;
      RECT 122.045 36.975 122.215 37.145 ;
      RECT 122.045 39.695 122.215 39.865 ;
      RECT 122.045 42.415 122.215 42.585 ;
      RECT 122.045 45.135 122.215 45.305 ;
      RECT 122.045 47.855 122.215 48.025 ;
      RECT 122.045 50.575 122.215 50.745 ;
      RECT 122.045 53.295 122.215 53.465 ;
      RECT 122.045 56.015 122.215 56.185 ;
      RECT 122.045 58.735 122.215 58.905 ;
      RECT 122.005 21.845 122.175 22.015 ;
      RECT 121.61 21.505 121.78 21.675 ;
      RECT 121.585 9.775 121.755 9.945 ;
      RECT 121.585 12.495 121.755 12.665 ;
      RECT 121.585 15.215 121.755 15.385 ;
      RECT 121.585 17.935 121.755 18.105 ;
      RECT 121.585 20.655 121.755 20.825 ;
      RECT 121.585 23.375 121.755 23.545 ;
      RECT 121.585 26.095 121.755 26.265 ;
      RECT 121.585 28.815 121.755 28.985 ;
      RECT 121.585 31.535 121.755 31.705 ;
      RECT 121.585 34.255 121.755 34.425 ;
      RECT 121.585 36.975 121.755 37.145 ;
      RECT 121.585 39.695 121.755 39.865 ;
      RECT 121.585 42.415 121.755 42.585 ;
      RECT 121.585 45.135 121.755 45.305 ;
      RECT 121.585 47.855 121.755 48.025 ;
      RECT 121.585 50.575 121.755 50.745 ;
      RECT 121.585 53.295 121.755 53.465 ;
      RECT 121.585 56.015 121.755 56.185 ;
      RECT 121.585 58.735 121.755 58.905 ;
      RECT 121.125 9.775 121.295 9.945 ;
      RECT 121.125 12.495 121.295 12.665 ;
      RECT 121.125 15.215 121.295 15.385 ;
      RECT 121.125 17.935 121.295 18.105 ;
      RECT 121.125 20.655 121.295 20.825 ;
      RECT 121.125 22.185 121.295 22.355 ;
      RECT 121.125 23.375 121.295 23.545 ;
      RECT 121.125 26.095 121.295 26.265 ;
      RECT 121.125 28.815 121.295 28.985 ;
      RECT 121.125 31.535 121.295 31.705 ;
      RECT 121.125 34.255 121.295 34.425 ;
      RECT 121.125 36.975 121.295 37.145 ;
      RECT 121.125 39.695 121.295 39.865 ;
      RECT 121.125 42.415 121.295 42.585 ;
      RECT 121.125 45.135 121.295 45.305 ;
      RECT 121.125 47.855 121.295 48.025 ;
      RECT 121.125 50.575 121.295 50.745 ;
      RECT 121.125 53.295 121.295 53.465 ;
      RECT 121.125 56.015 121.295 56.185 ;
      RECT 121.125 58.735 121.295 58.905 ;
      RECT 120.95 16.065 121.12 16.235 ;
      RECT 120.665 9.775 120.835 9.945 ;
      RECT 120.665 12.495 120.835 12.665 ;
      RECT 120.665 15.215 120.835 15.385 ;
      RECT 120.665 17.935 120.835 18.105 ;
      RECT 120.665 19.125 120.835 19.295 ;
      RECT 120.665 20.655 120.835 20.825 ;
      RECT 120.665 23.375 120.835 23.545 ;
      RECT 120.665 26.095 120.835 26.265 ;
      RECT 120.665 28.815 120.835 28.985 ;
      RECT 120.665 31.535 120.835 31.705 ;
      RECT 120.665 34.255 120.835 34.425 ;
      RECT 120.665 36.975 120.835 37.145 ;
      RECT 120.665 39.695 120.835 39.865 ;
      RECT 120.665 42.415 120.835 42.585 ;
      RECT 120.665 45.135 120.835 45.305 ;
      RECT 120.665 47.855 120.835 48.025 ;
      RECT 120.665 50.575 120.835 50.745 ;
      RECT 120.665 53.295 120.835 53.465 ;
      RECT 120.665 56.015 120.835 56.185 ;
      RECT 120.665 58.735 120.835 58.905 ;
      RECT 120.435 16.405 120.605 16.575 ;
      RECT 120.205 9.775 120.375 9.945 ;
      RECT 120.205 12.495 120.375 12.665 ;
      RECT 120.205 15.215 120.375 15.385 ;
      RECT 120.205 17.935 120.375 18.105 ;
      RECT 120.205 20.655 120.375 20.825 ;
      RECT 120.205 23.375 120.375 23.545 ;
      RECT 120.205 26.095 120.375 26.265 ;
      RECT 120.205 28.815 120.375 28.985 ;
      RECT 120.205 31.535 120.375 31.705 ;
      RECT 120.205 34.255 120.375 34.425 ;
      RECT 120.205 36.975 120.375 37.145 ;
      RECT 120.205 39.695 120.375 39.865 ;
      RECT 120.205 42.415 120.375 42.585 ;
      RECT 120.205 45.135 120.375 45.305 ;
      RECT 120.205 47.855 120.375 48.025 ;
      RECT 120.205 50.575 120.375 50.745 ;
      RECT 120.205 53.295 120.375 53.465 ;
      RECT 120.205 56.015 120.375 56.185 ;
      RECT 120.205 58.735 120.375 58.905 ;
      RECT 119.745 9.775 119.915 9.945 ;
      RECT 119.745 12.495 119.915 12.665 ;
      RECT 119.745 15.215 119.915 15.385 ;
      RECT 119.745 17.935 119.915 18.105 ;
      RECT 119.745 20.655 119.915 20.825 ;
      RECT 119.745 23.375 119.915 23.545 ;
      RECT 119.745 26.095 119.915 26.265 ;
      RECT 119.745 28.815 119.915 28.985 ;
      RECT 119.745 31.535 119.915 31.705 ;
      RECT 119.745 34.255 119.915 34.425 ;
      RECT 119.745 36.975 119.915 37.145 ;
      RECT 119.745 39.695 119.915 39.865 ;
      RECT 119.745 42.415 119.915 42.585 ;
      RECT 119.745 45.135 119.915 45.305 ;
      RECT 119.745 47.855 119.915 48.025 ;
      RECT 119.745 50.575 119.915 50.745 ;
      RECT 119.745 53.295 119.915 53.465 ;
      RECT 119.745 56.015 119.915 56.185 ;
      RECT 119.745 58.735 119.915 58.905 ;
      RECT 119.7 16.745 119.87 16.915 ;
      RECT 119.285 9.775 119.455 9.945 ;
      RECT 119.285 11.305 119.455 11.475 ;
      RECT 119.285 12.495 119.455 12.665 ;
      RECT 119.285 15.215 119.455 15.385 ;
      RECT 119.285 17.935 119.455 18.105 ;
      RECT 119.285 18.445 119.455 18.615 ;
      RECT 119.285 20.655 119.455 20.825 ;
      RECT 119.285 23.375 119.455 23.545 ;
      RECT 119.285 26.095 119.455 26.265 ;
      RECT 119.285 28.815 119.455 28.985 ;
      RECT 119.285 31.535 119.455 31.705 ;
      RECT 119.285 34.255 119.455 34.425 ;
      RECT 119.285 36.975 119.455 37.145 ;
      RECT 119.285 39.695 119.455 39.865 ;
      RECT 119.285 42.415 119.455 42.585 ;
      RECT 119.285 45.135 119.455 45.305 ;
      RECT 119.285 47.855 119.455 48.025 ;
      RECT 119.285 50.575 119.455 50.745 ;
      RECT 119.285 53.295 119.455 53.465 ;
      RECT 119.285 56.015 119.455 56.185 ;
      RECT 119.285 58.735 119.455 58.905 ;
      RECT 119.245 16.405 119.415 16.575 ;
      RECT 118.85 16.065 119.02 16.235 ;
      RECT 118.825 9.775 118.995 9.945 ;
      RECT 118.825 12.495 118.995 12.665 ;
      RECT 118.825 15.215 118.995 15.385 ;
      RECT 118.825 17.935 118.995 18.105 ;
      RECT 118.825 20.655 118.995 20.825 ;
      RECT 118.825 23.375 118.995 23.545 ;
      RECT 118.825 26.095 118.995 26.265 ;
      RECT 118.825 28.815 118.995 28.985 ;
      RECT 118.825 31.535 118.995 31.705 ;
      RECT 118.825 34.255 118.995 34.425 ;
      RECT 118.825 36.975 118.995 37.145 ;
      RECT 118.825 39.695 118.995 39.865 ;
      RECT 118.825 42.415 118.995 42.585 ;
      RECT 118.825 45.135 118.995 45.305 ;
      RECT 118.825 47.855 118.995 48.025 ;
      RECT 118.825 50.575 118.995 50.745 ;
      RECT 118.825 53.295 118.995 53.465 ;
      RECT 118.825 56.015 118.995 56.185 ;
      RECT 118.825 58.735 118.995 58.905 ;
      RECT 118.365 9.775 118.535 9.945 ;
      RECT 118.365 12.495 118.535 12.665 ;
      RECT 118.365 15.215 118.535 15.385 ;
      RECT 118.365 16.745 118.535 16.915 ;
      RECT 118.365 17.935 118.535 18.105 ;
      RECT 118.365 20.655 118.535 20.825 ;
      RECT 118.365 23.375 118.535 23.545 ;
      RECT 118.365 26.095 118.535 26.265 ;
      RECT 118.365 28.815 118.535 28.985 ;
      RECT 118.365 31.535 118.535 31.705 ;
      RECT 118.365 34.255 118.535 34.425 ;
      RECT 118.365 36.975 118.535 37.145 ;
      RECT 118.365 39.695 118.535 39.865 ;
      RECT 118.365 42.415 118.535 42.585 ;
      RECT 118.365 45.135 118.535 45.305 ;
      RECT 118.365 47.855 118.535 48.025 ;
      RECT 118.365 50.575 118.535 50.745 ;
      RECT 118.365 53.295 118.535 53.465 ;
      RECT 118.365 56.015 118.535 56.185 ;
      RECT 118.365 58.735 118.535 58.905 ;
      RECT 117.905 9.775 118.075 9.945 ;
      RECT 117.905 12.495 118.075 12.665 ;
      RECT 117.905 15.215 118.075 15.385 ;
      RECT 117.905 17.935 118.075 18.105 ;
      RECT 117.905 20.655 118.075 20.825 ;
      RECT 117.905 23.375 118.075 23.545 ;
      RECT 117.905 26.095 118.075 26.265 ;
      RECT 117.905 28.815 118.075 28.985 ;
      RECT 117.905 31.535 118.075 31.705 ;
      RECT 117.905 34.255 118.075 34.425 ;
      RECT 117.905 36.975 118.075 37.145 ;
      RECT 117.905 39.695 118.075 39.865 ;
      RECT 117.905 42.415 118.075 42.585 ;
      RECT 117.905 45.135 118.075 45.305 ;
      RECT 117.905 47.855 118.075 48.025 ;
      RECT 117.905 50.575 118.075 50.745 ;
      RECT 117.905 53.295 118.075 53.465 ;
      RECT 117.905 56.015 118.075 56.185 ;
      RECT 117.905 58.735 118.075 58.905 ;
      RECT 117.445 9.775 117.615 9.945 ;
      RECT 117.445 12.495 117.615 12.665 ;
      RECT 117.445 14.705 117.615 14.875 ;
      RECT 117.445 15.215 117.615 15.385 ;
      RECT 117.445 17.935 117.615 18.105 ;
      RECT 117.445 20.655 117.615 20.825 ;
      RECT 117.445 22.865 117.615 23.035 ;
      RECT 117.445 23.375 117.615 23.545 ;
      RECT 117.445 26.095 117.615 26.265 ;
      RECT 117.445 26.605 117.615 26.775 ;
      RECT 117.445 28.815 117.615 28.985 ;
      RECT 117.445 31.535 117.615 31.705 ;
      RECT 117.445 34.255 117.615 34.425 ;
      RECT 117.445 36.975 117.615 37.145 ;
      RECT 117.445 39.695 117.615 39.865 ;
      RECT 117.445 42.415 117.615 42.585 ;
      RECT 117.445 45.135 117.615 45.305 ;
      RECT 117.445 47.855 117.615 48.025 ;
      RECT 117.445 50.575 117.615 50.745 ;
      RECT 117.445 53.295 117.615 53.465 ;
      RECT 117.445 56.015 117.615 56.185 ;
      RECT 117.445 58.735 117.615 58.905 ;
      RECT 116.985 9.775 117.155 9.945 ;
      RECT 116.985 12.495 117.155 12.665 ;
      RECT 116.985 15.215 117.155 15.385 ;
      RECT 116.985 17.935 117.155 18.105 ;
      RECT 116.985 20.145 117.155 20.315 ;
      RECT 116.985 20.655 117.155 20.825 ;
      RECT 116.985 23.375 117.155 23.545 ;
      RECT 116.985 26.095 117.155 26.265 ;
      RECT 116.985 28.815 117.155 28.985 ;
      RECT 116.985 31.535 117.155 31.705 ;
      RECT 116.985 34.255 117.155 34.425 ;
      RECT 116.985 36.975 117.155 37.145 ;
      RECT 116.985 39.695 117.155 39.865 ;
      RECT 116.985 42.415 117.155 42.585 ;
      RECT 116.985 45.135 117.155 45.305 ;
      RECT 116.985 47.855 117.155 48.025 ;
      RECT 116.985 50.575 117.155 50.745 ;
      RECT 116.985 53.295 117.155 53.465 ;
      RECT 116.985 56.015 117.155 56.185 ;
      RECT 116.985 58.735 117.155 58.905 ;
      RECT 116.755 13.685 116.925 13.855 ;
      RECT 116.755 22.185 116.925 22.355 ;
      RECT 116.525 9.775 116.695 9.945 ;
      RECT 116.525 12.495 116.695 12.665 ;
      RECT 116.525 15.215 116.695 15.385 ;
      RECT 116.525 17.935 116.695 18.105 ;
      RECT 116.525 20.655 116.695 20.825 ;
      RECT 116.525 23.375 116.695 23.545 ;
      RECT 116.525 26.095 116.695 26.265 ;
      RECT 116.525 28.815 116.695 28.985 ;
      RECT 116.525 31.535 116.695 31.705 ;
      RECT 116.525 34.255 116.695 34.425 ;
      RECT 116.525 36.975 116.695 37.145 ;
      RECT 116.525 39.695 116.695 39.865 ;
      RECT 116.525 42.415 116.695 42.585 ;
      RECT 116.525 45.135 116.695 45.305 ;
      RECT 116.525 47.855 116.695 48.025 ;
      RECT 116.525 50.575 116.695 50.745 ;
      RECT 116.525 53.295 116.695 53.465 ;
      RECT 116.525 56.015 116.695 56.185 ;
      RECT 116.525 58.735 116.695 58.905 ;
      RECT 116.065 9.775 116.235 9.945 ;
      RECT 116.065 12.495 116.235 12.665 ;
      RECT 116.065 13.345 116.235 13.515 ;
      RECT 116.065 15.215 116.235 15.385 ;
      RECT 116.065 17.425 116.235 17.595 ;
      RECT 116.065 17.935 116.235 18.105 ;
      RECT 116.065 20.655 116.235 20.825 ;
      RECT 116.065 22.185 116.235 22.355 ;
      RECT 116.065 23.375 116.235 23.545 ;
      RECT 116.065 26.095 116.235 26.265 ;
      RECT 116.065 28.815 116.235 28.985 ;
      RECT 116.065 31.535 116.235 31.705 ;
      RECT 116.065 34.255 116.235 34.425 ;
      RECT 116.065 36.975 116.235 37.145 ;
      RECT 116.065 39.695 116.235 39.865 ;
      RECT 116.065 42.415 116.235 42.585 ;
      RECT 116.065 45.135 116.235 45.305 ;
      RECT 116.065 47.855 116.235 48.025 ;
      RECT 116.065 50.575 116.235 50.745 ;
      RECT 116.065 53.295 116.235 53.465 ;
      RECT 116.065 56.015 116.235 56.185 ;
      RECT 116.065 58.735 116.235 58.905 ;
      RECT 115.605 9.775 115.775 9.945 ;
      RECT 115.605 12.495 115.775 12.665 ;
      RECT 115.605 13.345 115.775 13.515 ;
      RECT 115.605 15.215 115.775 15.385 ;
      RECT 115.605 17.935 115.775 18.105 ;
      RECT 115.605 20.655 115.775 20.825 ;
      RECT 115.605 22.185 115.775 22.355 ;
      RECT 115.605 23.375 115.775 23.545 ;
      RECT 115.605 26.095 115.775 26.265 ;
      RECT 115.605 28.815 115.775 28.985 ;
      RECT 115.605 31.535 115.775 31.705 ;
      RECT 115.605 34.255 115.775 34.425 ;
      RECT 115.605 36.975 115.775 37.145 ;
      RECT 115.605 39.695 115.775 39.865 ;
      RECT 115.605 42.415 115.775 42.585 ;
      RECT 115.605 45.135 115.775 45.305 ;
      RECT 115.605 47.855 115.775 48.025 ;
      RECT 115.605 50.575 115.775 50.745 ;
      RECT 115.605 53.295 115.775 53.465 ;
      RECT 115.605 56.015 115.775 56.185 ;
      RECT 115.605 58.735 115.775 58.905 ;
      RECT 115.375 16.745 115.545 16.915 ;
      RECT 115.145 9.775 115.315 9.945 ;
      RECT 115.145 11.305 115.315 11.475 ;
      RECT 115.145 12.495 115.315 12.665 ;
      RECT 115.145 15.215 115.315 15.385 ;
      RECT 115.145 17.935 115.315 18.105 ;
      RECT 115.145 20.655 115.315 20.825 ;
      RECT 115.145 23.375 115.315 23.545 ;
      RECT 115.145 26.095 115.315 26.265 ;
      RECT 115.145 28.815 115.315 28.985 ;
      RECT 115.145 31.535 115.315 31.705 ;
      RECT 115.145 34.255 115.315 34.425 ;
      RECT 115.145 36.975 115.315 37.145 ;
      RECT 115.145 39.695 115.315 39.865 ;
      RECT 115.145 42.415 115.315 42.585 ;
      RECT 115.145 45.135 115.315 45.305 ;
      RECT 115.145 47.855 115.315 48.025 ;
      RECT 115.145 50.575 115.315 50.745 ;
      RECT 115.145 53.295 115.315 53.465 ;
      RECT 115.145 56.015 115.315 56.185 ;
      RECT 115.145 58.735 115.315 58.905 ;
      RECT 115.135 27.285 115.305 27.455 ;
      RECT 114.915 13.685 115.085 13.855 ;
      RECT 114.915 22.185 115.085 22.355 ;
      RECT 114.7 26.945 114.87 27.115 ;
      RECT 114.685 9.775 114.855 9.945 ;
      RECT 114.685 12.495 114.855 12.665 ;
      RECT 114.685 15.215 114.855 15.385 ;
      RECT 114.685 17.085 114.855 17.255 ;
      RECT 114.685 17.935 114.855 18.105 ;
      RECT 114.685 20.655 114.855 20.825 ;
      RECT 114.685 23.375 114.855 23.545 ;
      RECT 114.685 26.095 114.855 26.265 ;
      RECT 114.685 28.815 114.855 28.985 ;
      RECT 114.685 31.535 114.855 31.705 ;
      RECT 114.685 34.255 114.855 34.425 ;
      RECT 114.685 36.975 114.855 37.145 ;
      RECT 114.685 39.695 114.855 39.865 ;
      RECT 114.685 42.415 114.855 42.585 ;
      RECT 114.685 45.135 114.855 45.305 ;
      RECT 114.685 47.855 114.855 48.025 ;
      RECT 114.685 50.575 114.855 50.745 ;
      RECT 114.685 53.295 114.855 53.465 ;
      RECT 114.685 56.015 114.855 56.185 ;
      RECT 114.685 58.735 114.855 58.905 ;
      RECT 114.675 19.465 114.845 19.635 ;
      RECT 114.24 19.805 114.41 19.975 ;
      RECT 114.225 9.775 114.395 9.945 ;
      RECT 114.225 12.495 114.395 12.665 ;
      RECT 114.225 13.685 114.395 13.855 ;
      RECT 114.225 15.215 114.395 15.385 ;
      RECT 114.225 16.745 114.395 16.915 ;
      RECT 114.225 17.935 114.395 18.105 ;
      RECT 114.225 20.655 114.395 20.825 ;
      RECT 114.225 22.185 114.395 22.355 ;
      RECT 114.225 23.375 114.395 23.545 ;
      RECT 114.225 26.095 114.395 26.265 ;
      RECT 114.225 28.815 114.395 28.985 ;
      RECT 114.225 29.325 114.395 29.495 ;
      RECT 114.225 31.535 114.395 31.705 ;
      RECT 114.225 34.255 114.395 34.425 ;
      RECT 114.225 36.975 114.395 37.145 ;
      RECT 114.225 39.695 114.395 39.865 ;
      RECT 114.225 42.415 114.395 42.585 ;
      RECT 114.225 45.135 114.395 45.305 ;
      RECT 114.225 47.855 114.395 48.025 ;
      RECT 114.225 50.575 114.395 50.745 ;
      RECT 114.225 53.295 114.395 53.465 ;
      RECT 114.225 56.015 114.395 56.185 ;
      RECT 114.225 58.735 114.395 58.905 ;
      RECT 113.765 9.775 113.935 9.945 ;
      RECT 113.765 12.495 113.935 12.665 ;
      RECT 113.765 15.215 113.935 15.385 ;
      RECT 113.765 17.935 113.935 18.105 ;
      RECT 113.765 20.655 113.935 20.825 ;
      RECT 113.765 23.375 113.935 23.545 ;
      RECT 113.765 26.095 113.935 26.265 ;
      RECT 113.765 28.815 113.935 28.985 ;
      RECT 113.765 31.535 113.935 31.705 ;
      RECT 113.765 34.255 113.935 34.425 ;
      RECT 113.765 36.975 113.935 37.145 ;
      RECT 113.765 39.695 113.935 39.865 ;
      RECT 113.765 42.415 113.935 42.585 ;
      RECT 113.765 45.135 113.935 45.305 ;
      RECT 113.765 47.855 113.935 48.025 ;
      RECT 113.765 50.575 113.935 50.745 ;
      RECT 113.765 53.295 113.935 53.465 ;
      RECT 113.765 56.015 113.935 56.185 ;
      RECT 113.765 58.735 113.935 58.905 ;
      RECT 113.535 16.745 113.705 16.915 ;
      RECT 113.305 9.775 113.475 9.945 ;
      RECT 113.305 12.495 113.475 12.665 ;
      RECT 113.305 15.215 113.475 15.385 ;
      RECT 113.305 17.935 113.475 18.105 ;
      RECT 113.305 20.655 113.475 20.825 ;
      RECT 113.305 23.375 113.475 23.545 ;
      RECT 113.305 24.565 113.475 24.735 ;
      RECT 113.305 26.095 113.475 26.265 ;
      RECT 113.305 28.815 113.475 28.985 ;
      RECT 113.305 31.535 113.475 31.705 ;
      RECT 113.305 34.255 113.475 34.425 ;
      RECT 113.305 36.975 113.475 37.145 ;
      RECT 113.305 39.695 113.475 39.865 ;
      RECT 113.305 42.415 113.475 42.585 ;
      RECT 113.305 45.135 113.475 45.305 ;
      RECT 113.305 47.855 113.475 48.025 ;
      RECT 113.305 50.575 113.475 50.745 ;
      RECT 113.305 53.295 113.475 53.465 ;
      RECT 113.305 56.015 113.475 56.185 ;
      RECT 113.305 58.735 113.475 58.905 ;
      RECT 113.13 26.945 113.3 27.115 ;
      RECT 112.845 9.775 113.015 9.945 ;
      RECT 112.845 12.495 113.015 12.665 ;
      RECT 112.845 15.215 113.015 15.385 ;
      RECT 112.845 16.745 113.015 16.915 ;
      RECT 112.845 17.935 113.015 18.105 ;
      RECT 112.845 20.655 113.015 20.825 ;
      RECT 112.845 23.375 113.015 23.545 ;
      RECT 112.845 26.095 113.015 26.265 ;
      RECT 112.845 28.815 113.015 28.985 ;
      RECT 112.845 31.535 113.015 31.705 ;
      RECT 112.845 34.255 113.015 34.425 ;
      RECT 112.845 36.975 113.015 37.145 ;
      RECT 112.845 39.695 113.015 39.865 ;
      RECT 112.845 42.415 113.015 42.585 ;
      RECT 112.845 45.135 113.015 45.305 ;
      RECT 112.845 47.855 113.015 48.025 ;
      RECT 112.845 50.575 113.015 50.745 ;
      RECT 112.845 53.295 113.015 53.465 ;
      RECT 112.845 56.015 113.015 56.185 ;
      RECT 112.845 58.735 113.015 58.905 ;
      RECT 112.67 19.805 112.84 19.975 ;
      RECT 112.615 27.285 112.785 27.455 ;
      RECT 112.385 9.775 112.555 9.945 ;
      RECT 112.385 12.495 112.555 12.665 ;
      RECT 112.385 15.215 112.555 15.385 ;
      RECT 112.385 17.935 112.555 18.105 ;
      RECT 112.385 20.655 112.555 20.825 ;
      RECT 112.385 23.375 112.555 23.545 ;
      RECT 112.385 26.095 112.555 26.265 ;
      RECT 112.385 28.815 112.555 28.985 ;
      RECT 112.385 31.535 112.555 31.705 ;
      RECT 112.385 34.255 112.555 34.425 ;
      RECT 112.385 36.975 112.555 37.145 ;
      RECT 112.385 39.695 112.555 39.865 ;
      RECT 112.385 42.415 112.555 42.585 ;
      RECT 112.385 45.135 112.555 45.305 ;
      RECT 112.385 47.855 112.555 48.025 ;
      RECT 112.385 50.575 112.555 50.745 ;
      RECT 112.385 53.295 112.555 53.465 ;
      RECT 112.385 56.015 112.555 56.185 ;
      RECT 112.385 58.735 112.555 58.905 ;
      RECT 112.155 19.465 112.325 19.635 ;
      RECT 111.925 9.775 112.095 9.945 ;
      RECT 111.925 12.495 112.095 12.665 ;
      RECT 111.925 15.215 112.095 15.385 ;
      RECT 111.925 17.935 112.095 18.105 ;
      RECT 111.925 20.655 112.095 20.825 ;
      RECT 111.925 22.185 112.095 22.355 ;
      RECT 111.925 23.375 112.095 23.545 ;
      RECT 111.925 26.095 112.095 26.265 ;
      RECT 111.925 28.815 112.095 28.985 ;
      RECT 111.925 31.535 112.095 31.705 ;
      RECT 111.925 34.255 112.095 34.425 ;
      RECT 111.925 36.975 112.095 37.145 ;
      RECT 111.925 39.695 112.095 39.865 ;
      RECT 111.925 42.415 112.095 42.585 ;
      RECT 111.925 45.135 112.095 45.305 ;
      RECT 111.925 47.855 112.095 48.025 ;
      RECT 111.925 50.575 112.095 50.745 ;
      RECT 111.925 53.295 112.095 53.465 ;
      RECT 111.925 56.015 112.095 56.185 ;
      RECT 111.925 58.735 112.095 58.905 ;
      RECT 111.915 30.345 112.085 30.515 ;
      RECT 111.85 27.625 112.02 27.795 ;
      RECT 111.48 30.685 111.65 30.855 ;
      RECT 111.465 9.775 111.635 9.945 ;
      RECT 111.465 12.495 111.635 12.665 ;
      RECT 111.465 15.215 111.635 15.385 ;
      RECT 111.465 17.935 111.635 18.105 ;
      RECT 111.465 20.655 111.635 20.825 ;
      RECT 111.465 23.375 111.635 23.545 ;
      RECT 111.465 26.095 111.635 26.265 ;
      RECT 111.465 28.815 111.635 28.985 ;
      RECT 111.465 31.535 111.635 31.705 ;
      RECT 111.465 34.255 111.635 34.425 ;
      RECT 111.465 36.975 111.635 37.145 ;
      RECT 111.465 39.695 111.635 39.865 ;
      RECT 111.465 42.415 111.635 42.585 ;
      RECT 111.465 45.135 111.635 45.305 ;
      RECT 111.465 47.855 111.635 48.025 ;
      RECT 111.465 50.575 111.635 50.745 ;
      RECT 111.465 53.295 111.635 53.465 ;
      RECT 111.465 56.015 111.635 56.185 ;
      RECT 111.465 58.735 111.635 58.905 ;
      RECT 111.425 27.285 111.595 27.455 ;
      RECT 111.42 19.125 111.59 19.295 ;
      RECT 111.39 22.185 111.56 22.355 ;
      RECT 111.03 26.945 111.2 27.115 ;
      RECT 111.005 9.775 111.175 9.945 ;
      RECT 111.005 12.495 111.175 12.665 ;
      RECT 111.005 15.215 111.175 15.385 ;
      RECT 111.005 17.935 111.175 18.105 ;
      RECT 111.005 20.655 111.175 20.825 ;
      RECT 111.005 23.375 111.175 23.545 ;
      RECT 111.005 26.095 111.175 26.265 ;
      RECT 111.005 28.815 111.175 28.985 ;
      RECT 111.005 31.535 111.175 31.705 ;
      RECT 111.005 34.255 111.175 34.425 ;
      RECT 111.005 36.975 111.175 37.145 ;
      RECT 111.005 39.695 111.175 39.865 ;
      RECT 111.005 42.415 111.175 42.585 ;
      RECT 111.005 45.135 111.175 45.305 ;
      RECT 111.005 47.855 111.175 48.025 ;
      RECT 111.005 50.575 111.175 50.745 ;
      RECT 111.005 53.295 111.175 53.465 ;
      RECT 111.005 56.015 111.175 56.185 ;
      RECT 111.005 58.735 111.175 58.905 ;
      RECT 110.965 19.465 111.135 19.635 ;
      RECT 110.57 19.805 110.74 19.975 ;
      RECT 110.545 9.775 110.715 9.945 ;
      RECT 110.545 12.495 110.715 12.665 ;
      RECT 110.545 15.215 110.715 15.385 ;
      RECT 110.545 15.725 110.715 15.895 ;
      RECT 110.545 17.935 110.715 18.105 ;
      RECT 110.545 20.655 110.715 20.825 ;
      RECT 110.545 22.185 110.715 22.355 ;
      RECT 110.545 23.375 110.715 23.545 ;
      RECT 110.545 26.095 110.715 26.265 ;
      RECT 110.545 27.625 110.715 27.795 ;
      RECT 110.545 28.815 110.715 28.985 ;
      RECT 110.545 31.535 110.715 31.705 ;
      RECT 110.545 34.255 110.715 34.425 ;
      RECT 110.545 36.975 110.715 37.145 ;
      RECT 110.545 39.695 110.715 39.865 ;
      RECT 110.545 42.415 110.715 42.585 ;
      RECT 110.545 45.135 110.715 45.305 ;
      RECT 110.545 47.855 110.715 48.025 ;
      RECT 110.545 50.575 110.715 50.745 ;
      RECT 110.545 53.295 110.715 53.465 ;
      RECT 110.545 56.015 110.715 56.185 ;
      RECT 110.545 58.735 110.715 58.905 ;
      RECT 110.085 9.775 110.255 9.945 ;
      RECT 110.085 12.495 110.255 12.665 ;
      RECT 110.085 15.215 110.255 15.385 ;
      RECT 110.085 17.935 110.255 18.105 ;
      RECT 110.085 19.125 110.255 19.295 ;
      RECT 110.085 20.655 110.255 20.825 ;
      RECT 110.085 22.525 110.255 22.695 ;
      RECT 110.085 23.375 110.255 23.545 ;
      RECT 110.085 26.095 110.255 26.265 ;
      RECT 110.085 28.815 110.255 28.985 ;
      RECT 110.085 31.535 110.255 31.705 ;
      RECT 110.085 34.255 110.255 34.425 ;
      RECT 110.085 36.975 110.255 37.145 ;
      RECT 110.085 39.695 110.255 39.865 ;
      RECT 110.085 42.415 110.255 42.585 ;
      RECT 110.085 45.135 110.255 45.305 ;
      RECT 110.085 47.855 110.255 48.025 ;
      RECT 110.085 50.575 110.255 50.745 ;
      RECT 110.085 53.295 110.255 53.465 ;
      RECT 110.085 56.015 110.255 56.185 ;
      RECT 110.085 58.735 110.255 58.905 ;
      RECT 109.91 30.685 110.08 30.855 ;
      RECT 109.625 9.775 109.795 9.945 ;
      RECT 109.625 12.495 109.795 12.665 ;
      RECT 109.625 15.215 109.795 15.385 ;
      RECT 109.625 17.935 109.795 18.105 ;
      RECT 109.625 20.655 109.795 20.825 ;
      RECT 109.625 23.375 109.795 23.545 ;
      RECT 109.625 26.095 109.795 26.265 ;
      RECT 109.625 28.815 109.795 28.985 ;
      RECT 109.625 31.535 109.795 31.705 ;
      RECT 109.625 34.255 109.795 34.425 ;
      RECT 109.625 36.975 109.795 37.145 ;
      RECT 109.625 39.695 109.795 39.865 ;
      RECT 109.625 42.415 109.795 42.585 ;
      RECT 109.625 45.135 109.795 45.305 ;
      RECT 109.625 47.855 109.795 48.025 ;
      RECT 109.625 50.575 109.795 50.745 ;
      RECT 109.625 53.295 109.795 53.465 ;
      RECT 109.625 56.015 109.795 56.185 ;
      RECT 109.625 58.735 109.795 58.905 ;
      RECT 109.395 22.185 109.565 22.355 ;
      RECT 109.395 30.345 109.565 30.515 ;
      RECT 109.165 9.775 109.335 9.945 ;
      RECT 109.165 12.495 109.335 12.665 ;
      RECT 109.165 15.215 109.335 15.385 ;
      RECT 109.165 17.935 109.335 18.105 ;
      RECT 109.165 20.655 109.335 20.825 ;
      RECT 109.165 23.375 109.335 23.545 ;
      RECT 109.165 26.095 109.335 26.265 ;
      RECT 109.165 28.815 109.335 28.985 ;
      RECT 109.165 31.535 109.335 31.705 ;
      RECT 109.165 34.255 109.335 34.425 ;
      RECT 109.165 36.975 109.335 37.145 ;
      RECT 109.165 39.695 109.335 39.865 ;
      RECT 109.165 42.415 109.335 42.585 ;
      RECT 109.165 45.135 109.335 45.305 ;
      RECT 109.165 47.855 109.335 48.025 ;
      RECT 109.165 50.575 109.335 50.745 ;
      RECT 109.165 53.295 109.335 53.465 ;
      RECT 109.165 56.015 109.335 56.185 ;
      RECT 109.165 58.735 109.335 58.905 ;
      RECT 108.705 9.775 108.875 9.945 ;
      RECT 108.705 12.495 108.875 12.665 ;
      RECT 108.705 15.215 108.875 15.385 ;
      RECT 108.705 17.935 108.875 18.105 ;
      RECT 108.705 20.655 108.875 20.825 ;
      RECT 108.705 22.865 108.875 23.035 ;
      RECT 108.705 23.375 108.875 23.545 ;
      RECT 108.705 26.095 108.875 26.265 ;
      RECT 108.705 28.815 108.875 28.985 ;
      RECT 108.705 31.535 108.875 31.705 ;
      RECT 108.705 34.255 108.875 34.425 ;
      RECT 108.705 36.975 108.875 37.145 ;
      RECT 108.705 39.695 108.875 39.865 ;
      RECT 108.705 42.415 108.875 42.585 ;
      RECT 108.705 45.135 108.875 45.305 ;
      RECT 108.705 47.855 108.875 48.025 ;
      RECT 108.705 50.575 108.875 50.745 ;
      RECT 108.705 53.295 108.875 53.465 ;
      RECT 108.705 56.015 108.875 56.185 ;
      RECT 108.705 58.735 108.875 58.905 ;
      RECT 108.63 29.665 108.8 29.835 ;
      RECT 108.245 9.775 108.415 9.945 ;
      RECT 108.245 12.495 108.415 12.665 ;
      RECT 108.245 15.215 108.415 15.385 ;
      RECT 108.245 17.935 108.415 18.105 ;
      RECT 108.245 19.125 108.415 19.295 ;
      RECT 108.245 20.655 108.415 20.825 ;
      RECT 108.245 23.375 108.415 23.545 ;
      RECT 108.245 26.095 108.415 26.265 ;
      RECT 108.245 28.815 108.415 28.985 ;
      RECT 108.245 31.535 108.415 31.705 ;
      RECT 108.245 34.255 108.415 34.425 ;
      RECT 108.245 36.975 108.415 37.145 ;
      RECT 108.245 39.695 108.415 39.865 ;
      RECT 108.245 42.415 108.415 42.585 ;
      RECT 108.245 45.135 108.415 45.305 ;
      RECT 108.245 47.855 108.415 48.025 ;
      RECT 108.245 50.575 108.415 50.745 ;
      RECT 108.245 53.295 108.415 53.465 ;
      RECT 108.245 56.015 108.415 56.185 ;
      RECT 108.245 58.735 108.415 58.905 ;
      RECT 108.235 16.405 108.405 16.575 ;
      RECT 108.205 30.345 108.375 30.515 ;
      RECT 107.81 30.685 107.98 30.855 ;
      RECT 107.8 16.065 107.97 16.235 ;
      RECT 107.785 9.775 107.955 9.945 ;
      RECT 107.785 12.495 107.955 12.665 ;
      RECT 107.785 15.215 107.955 15.385 ;
      RECT 107.785 17.935 107.955 18.105 ;
      RECT 107.785 20.655 107.955 20.825 ;
      RECT 107.785 23.375 107.955 23.545 ;
      RECT 107.785 26.095 107.955 26.265 ;
      RECT 107.785 28.815 107.955 28.985 ;
      RECT 107.785 31.535 107.955 31.705 ;
      RECT 107.785 34.255 107.955 34.425 ;
      RECT 107.785 36.975 107.955 37.145 ;
      RECT 107.785 39.695 107.955 39.865 ;
      RECT 107.785 42.415 107.955 42.585 ;
      RECT 107.785 45.135 107.955 45.305 ;
      RECT 107.785 47.855 107.955 48.025 ;
      RECT 107.785 50.575 107.955 50.745 ;
      RECT 107.785 53.295 107.955 53.465 ;
      RECT 107.785 56.015 107.955 56.185 ;
      RECT 107.785 58.735 107.955 58.905 ;
      RECT 107.555 19.125 107.725 19.295 ;
      RECT 107.325 9.775 107.495 9.945 ;
      RECT 107.325 12.495 107.495 12.665 ;
      RECT 107.325 15.215 107.495 15.385 ;
      RECT 107.325 17.935 107.495 18.105 ;
      RECT 107.325 20.655 107.495 20.825 ;
      RECT 107.325 23.375 107.495 23.545 ;
      RECT 107.325 26.095 107.495 26.265 ;
      RECT 107.325 28.815 107.495 28.985 ;
      RECT 107.325 30.005 107.495 30.175 ;
      RECT 107.325 31.535 107.495 31.705 ;
      RECT 107.325 34.255 107.495 34.425 ;
      RECT 107.325 36.975 107.495 37.145 ;
      RECT 107.325 39.695 107.495 39.865 ;
      RECT 107.325 42.415 107.495 42.585 ;
      RECT 107.325 45.135 107.495 45.305 ;
      RECT 107.325 47.855 107.495 48.025 ;
      RECT 107.325 50.575 107.495 50.745 ;
      RECT 107.325 53.295 107.495 53.465 ;
      RECT 107.325 56.015 107.495 56.185 ;
      RECT 107.325 58.735 107.495 58.905 ;
      RECT 106.865 9.775 107.035 9.945 ;
      RECT 106.865 12.495 107.035 12.665 ;
      RECT 106.865 15.215 107.035 15.385 ;
      RECT 106.865 17.935 107.035 18.105 ;
      RECT 106.865 18.785 107.035 18.955 ;
      RECT 106.865 20.655 107.035 20.825 ;
      RECT 106.865 23.375 107.035 23.545 ;
      RECT 106.865 26.095 107.035 26.265 ;
      RECT 106.865 28.815 107.035 28.985 ;
      RECT 106.865 31.535 107.035 31.705 ;
      RECT 106.865 34.255 107.035 34.425 ;
      RECT 106.865 36.975 107.035 37.145 ;
      RECT 106.865 39.695 107.035 39.865 ;
      RECT 106.865 42.415 107.035 42.585 ;
      RECT 106.865 45.135 107.035 45.305 ;
      RECT 106.865 47.855 107.035 48.025 ;
      RECT 106.865 50.575 107.035 50.745 ;
      RECT 106.865 53.295 107.035 53.465 ;
      RECT 106.865 56.015 107.035 56.185 ;
      RECT 106.865 58.735 107.035 58.905 ;
      RECT 106.405 9.775 106.575 9.945 ;
      RECT 106.405 12.495 106.575 12.665 ;
      RECT 106.405 15.215 106.575 15.385 ;
      RECT 106.405 17.935 106.575 18.105 ;
      RECT 106.405 19.125 106.575 19.295 ;
      RECT 106.405 20.655 106.575 20.825 ;
      RECT 106.405 23.375 106.575 23.545 ;
      RECT 106.405 26.095 106.575 26.265 ;
      RECT 106.405 28.815 106.575 28.985 ;
      RECT 106.405 31.535 106.575 31.705 ;
      RECT 106.405 34.255 106.575 34.425 ;
      RECT 106.405 36.975 106.575 37.145 ;
      RECT 106.405 39.695 106.575 39.865 ;
      RECT 106.405 42.415 106.575 42.585 ;
      RECT 106.405 45.135 106.575 45.305 ;
      RECT 106.405 47.855 106.575 48.025 ;
      RECT 106.405 50.575 106.575 50.745 ;
      RECT 106.405 53.295 106.575 53.465 ;
      RECT 106.405 56.015 106.575 56.185 ;
      RECT 106.405 58.735 106.575 58.905 ;
      RECT 106.23 16.065 106.4 16.235 ;
      RECT 105.945 9.775 106.115 9.945 ;
      RECT 105.945 12.495 106.115 12.665 ;
      RECT 105.945 15.215 106.115 15.385 ;
      RECT 105.945 17.935 106.115 18.105 ;
      RECT 105.945 20.655 106.115 20.825 ;
      RECT 105.945 23.375 106.115 23.545 ;
      RECT 105.945 26.095 106.115 26.265 ;
      RECT 105.945 28.815 106.115 28.985 ;
      RECT 105.945 31.535 106.115 31.705 ;
      RECT 105.945 34.255 106.115 34.425 ;
      RECT 105.945 36.975 106.115 37.145 ;
      RECT 105.945 39.695 106.115 39.865 ;
      RECT 105.945 42.415 106.115 42.585 ;
      RECT 105.945 45.135 106.115 45.305 ;
      RECT 105.945 47.855 106.115 48.025 ;
      RECT 105.945 50.575 106.115 50.745 ;
      RECT 105.945 53.295 106.115 53.465 ;
      RECT 105.945 56.015 106.115 56.185 ;
      RECT 105.945 58.735 106.115 58.905 ;
      RECT 105.715 16.405 105.885 16.575 ;
      RECT 105.715 19.125 105.885 19.295 ;
      RECT 105.485 9.775 105.655 9.945 ;
      RECT 105.485 12.495 105.655 12.665 ;
      RECT 105.485 15.215 105.655 15.385 ;
      RECT 105.485 17.935 105.655 18.105 ;
      RECT 105.485 20.655 105.655 20.825 ;
      RECT 105.485 23.375 105.655 23.545 ;
      RECT 105.485 26.095 105.655 26.265 ;
      RECT 105.485 28.815 105.655 28.985 ;
      RECT 105.485 31.535 105.655 31.705 ;
      RECT 105.485 34.255 105.655 34.425 ;
      RECT 105.485 36.975 105.655 37.145 ;
      RECT 105.485 39.695 105.655 39.865 ;
      RECT 105.485 42.415 105.655 42.585 ;
      RECT 105.485 45.135 105.655 45.305 ;
      RECT 105.485 47.855 105.655 48.025 ;
      RECT 105.485 50.575 105.655 50.745 ;
      RECT 105.485 53.295 105.655 53.465 ;
      RECT 105.485 56.015 105.655 56.185 ;
      RECT 105.485 58.735 105.655 58.905 ;
      RECT 105.025 9.775 105.195 9.945 ;
      RECT 105.025 12.495 105.195 12.665 ;
      RECT 105.025 15.215 105.195 15.385 ;
      RECT 105.025 17.935 105.195 18.105 ;
      RECT 105.025 18.445 105.195 18.615 ;
      RECT 105.025 20.655 105.195 20.825 ;
      RECT 105.025 23.375 105.195 23.545 ;
      RECT 105.025 26.095 105.195 26.265 ;
      RECT 105.025 28.815 105.195 28.985 ;
      RECT 105.025 31.535 105.195 31.705 ;
      RECT 105.025 34.255 105.195 34.425 ;
      RECT 105.025 36.975 105.195 37.145 ;
      RECT 105.025 39.695 105.195 39.865 ;
      RECT 105.025 42.415 105.195 42.585 ;
      RECT 105.025 45.135 105.195 45.305 ;
      RECT 105.025 47.855 105.195 48.025 ;
      RECT 105.025 50.575 105.195 50.745 ;
      RECT 105.025 53.295 105.195 53.465 ;
      RECT 105.025 56.015 105.195 56.185 ;
      RECT 105.025 58.735 105.195 58.905 ;
      RECT 104.95 16.745 105.12 16.915 ;
      RECT 104.565 9.775 104.735 9.945 ;
      RECT 104.565 12.495 104.735 12.665 ;
      RECT 104.565 15.215 104.735 15.385 ;
      RECT 104.565 17.935 104.735 18.105 ;
      RECT 104.565 20.655 104.735 20.825 ;
      RECT 104.565 23.375 104.735 23.545 ;
      RECT 104.565 26.095 104.735 26.265 ;
      RECT 104.565 28.815 104.735 28.985 ;
      RECT 104.565 31.535 104.735 31.705 ;
      RECT 104.565 34.255 104.735 34.425 ;
      RECT 104.565 36.975 104.735 37.145 ;
      RECT 104.565 39.695 104.735 39.865 ;
      RECT 104.565 42.415 104.735 42.585 ;
      RECT 104.565 45.135 104.735 45.305 ;
      RECT 104.565 47.855 104.735 48.025 ;
      RECT 104.565 50.575 104.735 50.745 ;
      RECT 104.565 53.295 104.735 53.465 ;
      RECT 104.565 56.015 104.735 56.185 ;
      RECT 104.565 58.735 104.735 58.905 ;
      RECT 104.525 16.405 104.695 16.575 ;
      RECT 104.13 16.065 104.3 16.235 ;
      RECT 104.105 9.775 104.275 9.945 ;
      RECT 104.105 12.495 104.275 12.665 ;
      RECT 104.105 15.215 104.275 15.385 ;
      RECT 104.105 17.935 104.275 18.105 ;
      RECT 104.105 20.655 104.275 20.825 ;
      RECT 104.105 23.375 104.275 23.545 ;
      RECT 104.105 26.095 104.275 26.265 ;
      RECT 104.105 28.815 104.275 28.985 ;
      RECT 104.105 31.535 104.275 31.705 ;
      RECT 104.105 34.255 104.275 34.425 ;
      RECT 104.105 36.975 104.275 37.145 ;
      RECT 104.105 39.695 104.275 39.865 ;
      RECT 104.105 42.415 104.275 42.585 ;
      RECT 104.105 45.135 104.275 45.305 ;
      RECT 104.105 47.855 104.275 48.025 ;
      RECT 104.105 50.575 104.275 50.745 ;
      RECT 104.105 53.295 104.275 53.465 ;
      RECT 104.105 56.015 104.275 56.185 ;
      RECT 104.105 58.735 104.275 58.905 ;
      RECT 103.645 9.775 103.815 9.945 ;
      RECT 103.645 11.305 103.815 11.475 ;
      RECT 103.645 12.495 103.815 12.665 ;
      RECT 103.645 15.215 103.815 15.385 ;
      RECT 103.645 16.745 103.815 16.915 ;
      RECT 103.645 17.935 103.815 18.105 ;
      RECT 103.645 20.655 103.815 20.825 ;
      RECT 103.645 23.375 103.815 23.545 ;
      RECT 103.645 26.095 103.815 26.265 ;
      RECT 103.645 28.815 103.815 28.985 ;
      RECT 103.645 31.535 103.815 31.705 ;
      RECT 103.645 34.255 103.815 34.425 ;
      RECT 103.645 36.975 103.815 37.145 ;
      RECT 103.645 39.695 103.815 39.865 ;
      RECT 103.645 42.415 103.815 42.585 ;
      RECT 103.645 45.135 103.815 45.305 ;
      RECT 103.645 47.855 103.815 48.025 ;
      RECT 103.645 50.575 103.815 50.745 ;
      RECT 103.645 53.295 103.815 53.465 ;
      RECT 103.645 56.015 103.815 56.185 ;
      RECT 103.645 58.735 103.815 58.905 ;
      RECT 103.185 9.775 103.355 9.945 ;
      RECT 103.185 12.495 103.355 12.665 ;
      RECT 103.185 15.215 103.355 15.385 ;
      RECT 103.185 17.935 103.355 18.105 ;
      RECT 103.185 20.655 103.355 20.825 ;
      RECT 103.185 23.375 103.355 23.545 ;
      RECT 103.185 26.095 103.355 26.265 ;
      RECT 103.185 28.815 103.355 28.985 ;
      RECT 103.185 31.535 103.355 31.705 ;
      RECT 103.185 34.255 103.355 34.425 ;
      RECT 103.185 36.975 103.355 37.145 ;
      RECT 103.185 39.695 103.355 39.865 ;
      RECT 103.185 42.415 103.355 42.585 ;
      RECT 103.185 45.135 103.355 45.305 ;
      RECT 103.185 47.855 103.355 48.025 ;
      RECT 103.185 50.575 103.355 50.745 ;
      RECT 103.185 53.295 103.355 53.465 ;
      RECT 103.185 56.015 103.355 56.185 ;
      RECT 103.185 58.735 103.355 58.905 ;
      RECT 102.725 9.775 102.895 9.945 ;
      RECT 102.725 12.495 102.895 12.665 ;
      RECT 102.725 15.215 102.895 15.385 ;
      RECT 102.725 17.935 102.895 18.105 ;
      RECT 102.725 20.655 102.895 20.825 ;
      RECT 102.725 23.375 102.895 23.545 ;
      RECT 102.725 26.095 102.895 26.265 ;
      RECT 102.725 28.815 102.895 28.985 ;
      RECT 102.725 31.535 102.895 31.705 ;
      RECT 102.725 34.255 102.895 34.425 ;
      RECT 102.725 36.975 102.895 37.145 ;
      RECT 102.725 39.695 102.895 39.865 ;
      RECT 102.725 42.415 102.895 42.585 ;
      RECT 102.725 45.135 102.895 45.305 ;
      RECT 102.725 47.855 102.895 48.025 ;
      RECT 102.725 50.575 102.895 50.745 ;
      RECT 102.725 53.295 102.895 53.465 ;
      RECT 102.725 56.015 102.895 56.185 ;
      RECT 102.725 58.735 102.895 58.905 ;
      RECT 102.265 9.775 102.435 9.945 ;
      RECT 102.265 12.495 102.435 12.665 ;
      RECT 102.265 15.215 102.435 15.385 ;
      RECT 102.265 17.935 102.435 18.105 ;
      RECT 102.265 20.655 102.435 20.825 ;
      RECT 102.265 23.375 102.435 23.545 ;
      RECT 102.265 26.095 102.435 26.265 ;
      RECT 102.265 28.815 102.435 28.985 ;
      RECT 102.265 31.535 102.435 31.705 ;
      RECT 102.265 34.255 102.435 34.425 ;
      RECT 102.265 36.975 102.435 37.145 ;
      RECT 102.265 39.695 102.435 39.865 ;
      RECT 102.265 42.415 102.435 42.585 ;
      RECT 102.265 45.135 102.435 45.305 ;
      RECT 102.265 47.855 102.435 48.025 ;
      RECT 102.265 50.575 102.435 50.745 ;
      RECT 102.265 53.295 102.435 53.465 ;
      RECT 102.265 56.015 102.435 56.185 ;
      RECT 102.265 58.735 102.435 58.905 ;
      RECT 101.805 9.775 101.975 9.945 ;
      RECT 101.805 12.495 101.975 12.665 ;
      RECT 101.805 15.215 101.975 15.385 ;
      RECT 101.805 17.935 101.975 18.105 ;
      RECT 101.805 20.655 101.975 20.825 ;
      RECT 101.805 23.375 101.975 23.545 ;
      RECT 101.805 26.095 101.975 26.265 ;
      RECT 101.805 28.815 101.975 28.985 ;
      RECT 101.805 31.535 101.975 31.705 ;
      RECT 101.805 34.255 101.975 34.425 ;
      RECT 101.805 36.975 101.975 37.145 ;
      RECT 101.805 39.695 101.975 39.865 ;
      RECT 101.805 42.415 101.975 42.585 ;
      RECT 101.805 45.135 101.975 45.305 ;
      RECT 101.805 47.855 101.975 48.025 ;
      RECT 101.805 50.575 101.975 50.745 ;
      RECT 101.805 53.295 101.975 53.465 ;
      RECT 101.805 56.015 101.975 56.185 ;
      RECT 101.805 58.735 101.975 58.905 ;
      RECT 101.345 9.775 101.515 9.945 ;
      RECT 101.345 12.495 101.515 12.665 ;
      RECT 101.345 15.215 101.515 15.385 ;
      RECT 101.345 17.935 101.515 18.105 ;
      RECT 101.345 20.655 101.515 20.825 ;
      RECT 101.345 23.375 101.515 23.545 ;
      RECT 101.345 26.095 101.515 26.265 ;
      RECT 101.345 28.815 101.515 28.985 ;
      RECT 101.345 31.535 101.515 31.705 ;
      RECT 101.345 34.255 101.515 34.425 ;
      RECT 101.345 36.975 101.515 37.145 ;
      RECT 101.345 39.695 101.515 39.865 ;
      RECT 101.345 42.415 101.515 42.585 ;
      RECT 101.345 45.135 101.515 45.305 ;
      RECT 101.345 47.855 101.515 48.025 ;
      RECT 101.345 50.575 101.515 50.745 ;
      RECT 101.345 53.295 101.515 53.465 ;
      RECT 101.345 56.015 101.515 56.185 ;
      RECT 101.345 58.735 101.515 58.905 ;
      RECT 100.885 9.775 101.055 9.945 ;
      RECT 100.885 12.495 101.055 12.665 ;
      RECT 100.885 15.215 101.055 15.385 ;
      RECT 100.885 17.425 101.055 17.595 ;
      RECT 100.885 17.935 101.055 18.105 ;
      RECT 100.885 20.655 101.055 20.825 ;
      RECT 100.885 23.375 101.055 23.545 ;
      RECT 100.885 26.095 101.055 26.265 ;
      RECT 100.885 28.815 101.055 28.985 ;
      RECT 100.885 31.535 101.055 31.705 ;
      RECT 100.885 34.255 101.055 34.425 ;
      RECT 100.885 36.975 101.055 37.145 ;
      RECT 100.885 39.695 101.055 39.865 ;
      RECT 100.885 42.415 101.055 42.585 ;
      RECT 100.885 45.135 101.055 45.305 ;
      RECT 100.885 47.855 101.055 48.025 ;
      RECT 100.885 50.575 101.055 50.745 ;
      RECT 100.885 53.295 101.055 53.465 ;
      RECT 100.885 56.015 101.055 56.185 ;
      RECT 100.885 58.735 101.055 58.905 ;
      RECT 100.425 9.775 100.595 9.945 ;
      RECT 100.425 12.495 100.595 12.665 ;
      RECT 100.425 15.215 100.595 15.385 ;
      RECT 100.425 17.935 100.595 18.105 ;
      RECT 100.425 20.655 100.595 20.825 ;
      RECT 100.425 21.165 100.595 21.335 ;
      RECT 100.425 23.375 100.595 23.545 ;
      RECT 100.425 26.095 100.595 26.265 ;
      RECT 100.425 28.815 100.595 28.985 ;
      RECT 100.425 31.535 100.595 31.705 ;
      RECT 100.425 34.255 100.595 34.425 ;
      RECT 100.425 36.975 100.595 37.145 ;
      RECT 100.425 39.695 100.595 39.865 ;
      RECT 100.425 42.415 100.595 42.585 ;
      RECT 100.425 45.135 100.595 45.305 ;
      RECT 100.425 47.855 100.595 48.025 ;
      RECT 100.425 50.575 100.595 50.745 ;
      RECT 100.425 53.295 100.595 53.465 ;
      RECT 100.425 56.015 100.595 56.185 ;
      RECT 100.425 58.735 100.595 58.905 ;
      RECT 99.965 9.775 100.135 9.945 ;
      RECT 99.965 12.495 100.135 12.665 ;
      RECT 99.965 15.215 100.135 15.385 ;
      RECT 99.965 17.935 100.135 18.105 ;
      RECT 99.965 20.655 100.135 20.825 ;
      RECT 99.965 23.375 100.135 23.545 ;
      RECT 99.965 26.095 100.135 26.265 ;
      RECT 99.965 28.815 100.135 28.985 ;
      RECT 99.965 31.535 100.135 31.705 ;
      RECT 99.965 34.255 100.135 34.425 ;
      RECT 99.965 34.765 100.135 34.935 ;
      RECT 99.965 36.975 100.135 37.145 ;
      RECT 99.965 39.695 100.135 39.865 ;
      RECT 99.965 42.415 100.135 42.585 ;
      RECT 99.965 45.135 100.135 45.305 ;
      RECT 99.965 47.855 100.135 48.025 ;
      RECT 99.965 50.575 100.135 50.745 ;
      RECT 99.965 53.295 100.135 53.465 ;
      RECT 99.965 56.015 100.135 56.185 ;
      RECT 99.965 58.735 100.135 58.905 ;
      RECT 99.505 9.775 99.675 9.945 ;
      RECT 99.505 12.495 99.675 12.665 ;
      RECT 99.505 15.215 99.675 15.385 ;
      RECT 99.505 17.935 99.675 18.105 ;
      RECT 99.505 20.655 99.675 20.825 ;
      RECT 99.505 23.375 99.675 23.545 ;
      RECT 99.505 26.095 99.675 26.265 ;
      RECT 99.505 28.815 99.675 28.985 ;
      RECT 99.505 31.535 99.675 31.705 ;
      RECT 99.505 34.255 99.675 34.425 ;
      RECT 99.505 36.975 99.675 37.145 ;
      RECT 99.505 39.695 99.675 39.865 ;
      RECT 99.505 42.415 99.675 42.585 ;
      RECT 99.505 45.135 99.675 45.305 ;
      RECT 99.505 47.855 99.675 48.025 ;
      RECT 99.505 50.575 99.675 50.745 ;
      RECT 99.505 53.295 99.675 53.465 ;
      RECT 99.505 56.015 99.675 56.185 ;
      RECT 99.505 58.735 99.675 58.905 ;
      RECT 99.045 9.775 99.215 9.945 ;
      RECT 99.045 12.495 99.215 12.665 ;
      RECT 99.045 15.215 99.215 15.385 ;
      RECT 99.045 17.935 99.215 18.105 ;
      RECT 99.045 20.655 99.215 20.825 ;
      RECT 99.045 23.375 99.215 23.545 ;
      RECT 99.045 26.095 99.215 26.265 ;
      RECT 99.045 28.815 99.215 28.985 ;
      RECT 99.045 31.535 99.215 31.705 ;
      RECT 99.045 34.255 99.215 34.425 ;
      RECT 99.045 36.975 99.215 37.145 ;
      RECT 99.045 39.695 99.215 39.865 ;
      RECT 99.045 42.415 99.215 42.585 ;
      RECT 99.045 45.135 99.215 45.305 ;
      RECT 99.045 47.855 99.215 48.025 ;
      RECT 99.045 50.575 99.215 50.745 ;
      RECT 99.045 53.295 99.215 53.465 ;
      RECT 99.045 56.015 99.215 56.185 ;
      RECT 99.045 58.735 99.215 58.905 ;
      RECT 98.585 9.775 98.755 9.945 ;
      RECT 98.585 12.495 98.755 12.665 ;
      RECT 98.585 15.215 98.755 15.385 ;
      RECT 98.585 17.935 98.755 18.105 ;
      RECT 98.585 20.655 98.755 20.825 ;
      RECT 98.585 23.375 98.755 23.545 ;
      RECT 98.585 26.095 98.755 26.265 ;
      RECT 98.585 28.815 98.755 28.985 ;
      RECT 98.585 31.535 98.755 31.705 ;
      RECT 98.585 34.255 98.755 34.425 ;
      RECT 98.585 36.975 98.755 37.145 ;
      RECT 98.585 39.695 98.755 39.865 ;
      RECT 98.585 42.415 98.755 42.585 ;
      RECT 98.585 45.135 98.755 45.305 ;
      RECT 98.585 47.855 98.755 48.025 ;
      RECT 98.585 50.575 98.755 50.745 ;
      RECT 98.585 53.295 98.755 53.465 ;
      RECT 98.585 56.015 98.755 56.185 ;
      RECT 98.585 58.735 98.755 58.905 ;
      RECT 98.575 16.405 98.745 16.575 ;
      RECT 98.14 16.065 98.31 16.235 ;
      RECT 98.125 9.775 98.295 9.945 ;
      RECT 98.125 12.495 98.295 12.665 ;
      RECT 98.125 15.215 98.295 15.385 ;
      RECT 98.125 17.935 98.295 18.105 ;
      RECT 98.125 18.445 98.295 18.615 ;
      RECT 98.125 20.655 98.295 20.825 ;
      RECT 98.125 23.375 98.295 23.545 ;
      RECT 98.125 23.885 98.295 24.055 ;
      RECT 98.125 26.095 98.295 26.265 ;
      RECT 98.125 28.815 98.295 28.985 ;
      RECT 98.125 31.535 98.295 31.705 ;
      RECT 98.125 33.745 98.295 33.915 ;
      RECT 98.125 34.255 98.295 34.425 ;
      RECT 98.125 36.975 98.295 37.145 ;
      RECT 98.125 39.695 98.295 39.865 ;
      RECT 98.125 42.415 98.295 42.585 ;
      RECT 98.125 45.135 98.295 45.305 ;
      RECT 98.125 47.855 98.295 48.025 ;
      RECT 98.125 50.575 98.295 50.745 ;
      RECT 98.125 53.295 98.295 53.465 ;
      RECT 98.125 56.015 98.295 56.185 ;
      RECT 98.125 58.735 98.295 58.905 ;
      RECT 98.115 21.845 98.285 22.015 ;
      RECT 97.68 21.505 97.85 21.675 ;
      RECT 97.665 9.775 97.835 9.945 ;
      RECT 97.665 12.495 97.835 12.665 ;
      RECT 97.665 15.215 97.835 15.385 ;
      RECT 97.665 17.935 97.835 18.105 ;
      RECT 97.665 20.655 97.835 20.825 ;
      RECT 97.665 23.375 97.835 23.545 ;
      RECT 97.665 26.095 97.835 26.265 ;
      RECT 97.665 28.815 97.835 28.985 ;
      RECT 97.665 31.535 97.835 31.705 ;
      RECT 97.665 34.255 97.835 34.425 ;
      RECT 97.665 36.975 97.835 37.145 ;
      RECT 97.665 39.695 97.835 39.865 ;
      RECT 97.665 42.415 97.835 42.585 ;
      RECT 97.665 45.135 97.835 45.305 ;
      RECT 97.665 47.855 97.835 48.025 ;
      RECT 97.665 50.575 97.835 50.745 ;
      RECT 97.665 53.295 97.835 53.465 ;
      RECT 97.665 56.015 97.835 56.185 ;
      RECT 97.665 58.735 97.835 58.905 ;
      RECT 97.655 35.785 97.825 35.955 ;
      RECT 97.435 19.125 97.605 19.295 ;
      RECT 97.435 24.565 97.605 24.735 ;
      RECT 97.435 33.065 97.605 33.235 ;
      RECT 97.22 36.125 97.39 36.295 ;
      RECT 97.205 9.775 97.375 9.945 ;
      RECT 97.205 11.305 97.375 11.475 ;
      RECT 97.205 12.495 97.375 12.665 ;
      RECT 97.205 15.215 97.375 15.385 ;
      RECT 97.205 17.935 97.375 18.105 ;
      RECT 97.205 20.655 97.375 20.825 ;
      RECT 97.205 23.375 97.375 23.545 ;
      RECT 97.205 26.095 97.375 26.265 ;
      RECT 97.205 28.815 97.375 28.985 ;
      RECT 97.205 31.535 97.375 31.705 ;
      RECT 97.205 34.255 97.375 34.425 ;
      RECT 97.205 36.975 97.375 37.145 ;
      RECT 97.205 39.695 97.375 39.865 ;
      RECT 97.205 42.415 97.375 42.585 ;
      RECT 97.205 45.135 97.375 45.305 ;
      RECT 97.205 47.855 97.375 48.025 ;
      RECT 97.205 50.575 97.375 50.745 ;
      RECT 97.205 53.295 97.375 53.465 ;
      RECT 97.205 56.015 97.375 56.185 ;
      RECT 97.205 58.735 97.375 58.905 ;
      RECT 96.745 9.775 96.915 9.945 ;
      RECT 96.745 12.495 96.915 12.665 ;
      RECT 96.745 15.215 96.915 15.385 ;
      RECT 96.745 17.935 96.915 18.105 ;
      RECT 96.745 19.125 96.915 19.295 ;
      RECT 96.745 20.655 96.915 20.825 ;
      RECT 96.745 23.375 96.915 23.545 ;
      RECT 96.745 24.565 96.915 24.735 ;
      RECT 96.745 26.095 96.915 26.265 ;
      RECT 96.745 28.815 96.915 28.985 ;
      RECT 96.745 31.535 96.915 31.705 ;
      RECT 96.745 33.065 96.915 33.235 ;
      RECT 96.745 34.255 96.915 34.425 ;
      RECT 96.745 36.975 96.915 37.145 ;
      RECT 96.745 39.695 96.915 39.865 ;
      RECT 96.745 42.415 96.915 42.585 ;
      RECT 96.745 45.135 96.915 45.305 ;
      RECT 96.745 47.855 96.915 48.025 ;
      RECT 96.745 50.575 96.915 50.745 ;
      RECT 96.745 53.295 96.915 53.465 ;
      RECT 96.745 56.015 96.915 56.185 ;
      RECT 96.745 58.735 96.915 58.905 ;
      RECT 96.57 16.065 96.74 16.235 ;
      RECT 96.285 9.775 96.455 9.945 ;
      RECT 96.285 12.495 96.455 12.665 ;
      RECT 96.285 15.215 96.455 15.385 ;
      RECT 96.285 17.935 96.455 18.105 ;
      RECT 96.285 18.785 96.455 18.955 ;
      RECT 96.285 20.655 96.455 20.825 ;
      RECT 96.285 23.375 96.455 23.545 ;
      RECT 96.285 24.225 96.455 24.395 ;
      RECT 96.285 26.095 96.455 26.265 ;
      RECT 96.285 28.815 96.455 28.985 ;
      RECT 96.285 31.535 96.455 31.705 ;
      RECT 96.285 33.405 96.455 33.575 ;
      RECT 96.285 34.255 96.455 34.425 ;
      RECT 96.285 36.975 96.455 37.145 ;
      RECT 96.285 39.695 96.455 39.865 ;
      RECT 96.285 42.415 96.455 42.585 ;
      RECT 96.285 45.135 96.455 45.305 ;
      RECT 96.285 47.855 96.455 48.025 ;
      RECT 96.285 50.575 96.455 50.745 ;
      RECT 96.285 53.295 96.455 53.465 ;
      RECT 96.285 56.015 96.455 56.185 ;
      RECT 96.285 58.735 96.455 58.905 ;
      RECT 96.11 21.505 96.28 21.675 ;
      RECT 96.055 16.405 96.225 16.575 ;
      RECT 95.825 9.775 95.995 9.945 ;
      RECT 95.825 12.495 95.995 12.665 ;
      RECT 95.825 15.215 95.995 15.385 ;
      RECT 95.825 17.935 95.995 18.105 ;
      RECT 95.825 20.655 95.995 20.825 ;
      RECT 95.825 23.375 95.995 23.545 ;
      RECT 95.825 26.095 95.995 26.265 ;
      RECT 95.825 28.815 95.995 28.985 ;
      RECT 95.825 31.535 95.995 31.705 ;
      RECT 95.825 34.255 95.995 34.425 ;
      RECT 95.825 36.975 95.995 37.145 ;
      RECT 95.825 39.695 95.995 39.865 ;
      RECT 95.825 42.415 95.995 42.585 ;
      RECT 95.825 45.135 95.995 45.305 ;
      RECT 95.825 47.855 95.995 48.025 ;
      RECT 95.825 50.575 95.995 50.745 ;
      RECT 95.825 53.295 95.995 53.465 ;
      RECT 95.825 56.015 95.995 56.185 ;
      RECT 95.825 58.735 95.995 58.905 ;
      RECT 95.65 36.125 95.82 36.295 ;
      RECT 95.595 19.125 95.765 19.295 ;
      RECT 95.595 21.845 95.765 22.015 ;
      RECT 95.595 24.565 95.765 24.735 ;
      RECT 95.595 33.065 95.765 33.235 ;
      RECT 95.365 9.775 95.535 9.945 ;
      RECT 95.365 12.495 95.535 12.665 ;
      RECT 95.365 15.215 95.535 15.385 ;
      RECT 95.365 17.935 95.535 18.105 ;
      RECT 95.365 20.655 95.535 20.825 ;
      RECT 95.365 23.375 95.535 23.545 ;
      RECT 95.365 26.095 95.535 26.265 ;
      RECT 95.365 28.815 95.535 28.985 ;
      RECT 95.365 31.535 95.535 31.705 ;
      RECT 95.365 34.255 95.535 34.425 ;
      RECT 95.365 36.975 95.535 37.145 ;
      RECT 95.365 39.695 95.535 39.865 ;
      RECT 95.365 42.415 95.535 42.585 ;
      RECT 95.365 45.135 95.535 45.305 ;
      RECT 95.365 47.855 95.535 48.025 ;
      RECT 95.365 50.575 95.535 50.745 ;
      RECT 95.365 53.295 95.535 53.465 ;
      RECT 95.365 56.015 95.535 56.185 ;
      RECT 95.365 58.735 95.535 58.905 ;
      RECT 95.29 16.745 95.46 16.915 ;
      RECT 95.135 35.785 95.305 35.955 ;
      RECT 94.905 9.775 95.075 9.945 ;
      RECT 94.905 12.495 95.075 12.665 ;
      RECT 94.905 15.215 95.075 15.385 ;
      RECT 94.905 17.935 95.075 18.105 ;
      RECT 94.905 19.125 95.075 19.295 ;
      RECT 94.905 20.655 95.075 20.825 ;
      RECT 94.905 23.375 95.075 23.545 ;
      RECT 94.905 24.565 95.075 24.735 ;
      RECT 94.905 26.095 95.075 26.265 ;
      RECT 94.905 28.815 95.075 28.985 ;
      RECT 94.905 31.535 95.075 31.705 ;
      RECT 94.905 33.065 95.075 33.235 ;
      RECT 94.905 34.255 95.075 34.425 ;
      RECT 94.905 36.975 95.075 37.145 ;
      RECT 94.905 39.695 95.075 39.865 ;
      RECT 94.905 42.415 95.075 42.585 ;
      RECT 94.905 45.135 95.075 45.305 ;
      RECT 94.905 47.855 95.075 48.025 ;
      RECT 94.905 50.575 95.075 50.745 ;
      RECT 94.905 53.295 95.075 53.465 ;
      RECT 94.905 56.015 95.075 56.185 ;
      RECT 94.905 58.735 95.075 58.905 ;
      RECT 94.865 16.405 95.035 16.575 ;
      RECT 94.86 22.185 95.03 22.355 ;
      RECT 94.47 16.065 94.64 16.235 ;
      RECT 94.445 9.775 94.615 9.945 ;
      RECT 94.445 12.495 94.615 12.665 ;
      RECT 94.445 15.215 94.615 15.385 ;
      RECT 94.445 17.935 94.615 18.105 ;
      RECT 94.445 20.655 94.615 20.825 ;
      RECT 94.445 23.375 94.615 23.545 ;
      RECT 94.445 26.095 94.615 26.265 ;
      RECT 94.445 28.815 94.615 28.985 ;
      RECT 94.445 31.535 94.615 31.705 ;
      RECT 94.445 34.255 94.615 34.425 ;
      RECT 94.445 36.975 94.615 37.145 ;
      RECT 94.445 39.695 94.615 39.865 ;
      RECT 94.445 42.415 94.615 42.585 ;
      RECT 94.445 45.135 94.615 45.305 ;
      RECT 94.445 47.855 94.615 48.025 ;
      RECT 94.445 50.575 94.615 50.745 ;
      RECT 94.445 53.295 94.615 53.465 ;
      RECT 94.445 56.015 94.615 56.185 ;
      RECT 94.445 58.735 94.615 58.905 ;
      RECT 94.405 21.845 94.575 22.015 ;
      RECT 94.4 35.105 94.57 35.275 ;
      RECT 94.01 21.505 94.18 21.675 ;
      RECT 93.985 9.775 94.155 9.945 ;
      RECT 93.985 12.495 94.155 12.665 ;
      RECT 93.985 15.215 94.155 15.385 ;
      RECT 93.985 16.745 94.155 16.915 ;
      RECT 93.985 17.935 94.155 18.105 ;
      RECT 93.985 20.655 94.155 20.825 ;
      RECT 93.985 23.375 94.155 23.545 ;
      RECT 93.985 26.095 94.155 26.265 ;
      RECT 93.985 28.815 94.155 28.985 ;
      RECT 93.985 31.535 94.155 31.705 ;
      RECT 93.985 34.255 94.155 34.425 ;
      RECT 93.985 36.975 94.155 37.145 ;
      RECT 93.985 39.695 94.155 39.865 ;
      RECT 93.985 42.415 94.155 42.585 ;
      RECT 93.985 45.135 94.155 45.305 ;
      RECT 93.985 47.855 94.155 48.025 ;
      RECT 93.985 50.575 94.155 50.745 ;
      RECT 93.985 53.295 94.155 53.465 ;
      RECT 93.985 56.015 94.155 56.185 ;
      RECT 93.985 58.735 94.155 58.905 ;
      RECT 93.945 35.785 94.115 35.955 ;
      RECT 93.55 36.125 93.72 36.295 ;
      RECT 93.525 9.775 93.695 9.945 ;
      RECT 93.525 12.495 93.695 12.665 ;
      RECT 93.525 15.215 93.695 15.385 ;
      RECT 93.525 17.935 93.695 18.105 ;
      RECT 93.525 20.655 93.695 20.825 ;
      RECT 93.525 22.185 93.695 22.355 ;
      RECT 93.525 23.375 93.695 23.545 ;
      RECT 93.525 26.095 93.695 26.265 ;
      RECT 93.525 28.815 93.695 28.985 ;
      RECT 93.525 31.535 93.695 31.705 ;
      RECT 93.525 34.255 93.695 34.425 ;
      RECT 93.525 36.975 93.695 37.145 ;
      RECT 93.525 39.695 93.695 39.865 ;
      RECT 93.525 42.415 93.695 42.585 ;
      RECT 93.525 45.135 93.695 45.305 ;
      RECT 93.525 47.855 93.695 48.025 ;
      RECT 93.525 50.575 93.695 50.745 ;
      RECT 93.525 53.295 93.695 53.465 ;
      RECT 93.525 56.015 93.695 56.185 ;
      RECT 93.525 58.735 93.695 58.905 ;
      RECT 93.065 9.775 93.235 9.945 ;
      RECT 93.065 12.495 93.235 12.665 ;
      RECT 93.065 15.215 93.235 15.385 ;
      RECT 93.065 17.935 93.235 18.105 ;
      RECT 93.065 20.655 93.235 20.825 ;
      RECT 93.065 23.375 93.235 23.545 ;
      RECT 93.065 26.095 93.235 26.265 ;
      RECT 93.065 28.815 93.235 28.985 ;
      RECT 93.065 31.535 93.235 31.705 ;
      RECT 93.065 34.255 93.235 34.425 ;
      RECT 93.065 35.445 93.235 35.615 ;
      RECT 93.065 36.975 93.235 37.145 ;
      RECT 93.065 39.695 93.235 39.865 ;
      RECT 93.065 42.415 93.235 42.585 ;
      RECT 93.065 45.135 93.235 45.305 ;
      RECT 93.065 47.855 93.235 48.025 ;
      RECT 93.065 50.575 93.235 50.745 ;
      RECT 93.065 53.295 93.235 53.465 ;
      RECT 93.065 56.015 93.235 56.185 ;
      RECT 93.065 58.735 93.235 58.905 ;
      RECT 92.605 9.775 92.775 9.945 ;
      RECT 92.605 12.495 92.775 12.665 ;
      RECT 92.605 15.215 92.775 15.385 ;
      RECT 92.605 17.935 92.775 18.105 ;
      RECT 92.605 20.655 92.775 20.825 ;
      RECT 92.605 23.375 92.775 23.545 ;
      RECT 92.605 26.095 92.775 26.265 ;
      RECT 92.605 28.815 92.775 28.985 ;
      RECT 92.605 31.535 92.775 31.705 ;
      RECT 92.605 34.255 92.775 34.425 ;
      RECT 92.605 36.975 92.775 37.145 ;
      RECT 92.605 39.695 92.775 39.865 ;
      RECT 92.605 42.415 92.775 42.585 ;
      RECT 92.605 45.135 92.775 45.305 ;
      RECT 92.605 47.855 92.775 48.025 ;
      RECT 92.605 50.575 92.775 50.745 ;
      RECT 92.605 53.295 92.775 53.465 ;
      RECT 92.605 56.015 92.775 56.185 ;
      RECT 92.605 58.735 92.775 58.905 ;
      RECT 92.145 9.775 92.315 9.945 ;
      RECT 92.145 12.495 92.315 12.665 ;
      RECT 92.145 15.215 92.315 15.385 ;
      RECT 92.145 17.935 92.315 18.105 ;
      RECT 92.145 20.655 92.315 20.825 ;
      RECT 92.145 23.375 92.315 23.545 ;
      RECT 92.145 26.095 92.315 26.265 ;
      RECT 92.145 28.815 92.315 28.985 ;
      RECT 92.145 31.535 92.315 31.705 ;
      RECT 92.145 34.255 92.315 34.425 ;
      RECT 92.145 36.975 92.315 37.145 ;
      RECT 92.145 39.695 92.315 39.865 ;
      RECT 92.145 42.415 92.315 42.585 ;
      RECT 92.145 45.135 92.315 45.305 ;
      RECT 92.145 47.855 92.315 48.025 ;
      RECT 92.145 50.575 92.315 50.745 ;
      RECT 92.145 53.295 92.315 53.465 ;
      RECT 92.145 56.015 92.315 56.185 ;
      RECT 92.145 58.735 92.315 58.905 ;
      RECT 91.685 9.775 91.855 9.945 ;
      RECT 91.685 11.305 91.855 11.475 ;
      RECT 91.685 12.495 91.855 12.665 ;
      RECT 91.685 15.215 91.855 15.385 ;
      RECT 91.685 17.935 91.855 18.105 ;
      RECT 91.685 20.655 91.855 20.825 ;
      RECT 91.685 23.375 91.855 23.545 ;
      RECT 91.685 26.095 91.855 26.265 ;
      RECT 91.685 28.815 91.855 28.985 ;
      RECT 91.685 31.535 91.855 31.705 ;
      RECT 91.685 34.255 91.855 34.425 ;
      RECT 91.685 36.975 91.855 37.145 ;
      RECT 91.685 39.695 91.855 39.865 ;
      RECT 91.685 42.415 91.855 42.585 ;
      RECT 91.685 45.135 91.855 45.305 ;
      RECT 91.685 47.855 91.855 48.025 ;
      RECT 91.685 50.575 91.855 50.745 ;
      RECT 91.685 53.295 91.855 53.465 ;
      RECT 91.685 56.015 91.855 56.185 ;
      RECT 91.685 58.735 91.855 58.905 ;
      RECT 91.225 9.775 91.395 9.945 ;
      RECT 91.225 12.495 91.395 12.665 ;
      RECT 91.225 15.215 91.395 15.385 ;
      RECT 91.225 17.935 91.395 18.105 ;
      RECT 91.225 20.655 91.395 20.825 ;
      RECT 91.225 23.375 91.395 23.545 ;
      RECT 91.225 26.095 91.395 26.265 ;
      RECT 91.225 28.815 91.395 28.985 ;
      RECT 91.225 31.535 91.395 31.705 ;
      RECT 91.225 34.255 91.395 34.425 ;
      RECT 91.225 36.975 91.395 37.145 ;
      RECT 91.225 39.695 91.395 39.865 ;
      RECT 91.225 42.415 91.395 42.585 ;
      RECT 91.225 45.135 91.395 45.305 ;
      RECT 91.225 47.855 91.395 48.025 ;
      RECT 91.225 50.575 91.395 50.745 ;
      RECT 91.225 53.295 91.395 53.465 ;
      RECT 91.225 56.015 91.395 56.185 ;
      RECT 91.225 58.735 91.395 58.905 ;
      RECT 90.765 9.775 90.935 9.945 ;
      RECT 90.765 12.495 90.935 12.665 ;
      RECT 90.765 15.215 90.935 15.385 ;
      RECT 90.765 17.935 90.935 18.105 ;
      RECT 90.765 20.655 90.935 20.825 ;
      RECT 90.765 23.375 90.935 23.545 ;
      RECT 90.765 26.095 90.935 26.265 ;
      RECT 90.765 28.815 90.935 28.985 ;
      RECT 90.765 31.535 90.935 31.705 ;
      RECT 90.765 34.255 90.935 34.425 ;
      RECT 90.765 36.975 90.935 37.145 ;
      RECT 90.765 39.695 90.935 39.865 ;
      RECT 90.765 42.415 90.935 42.585 ;
      RECT 90.765 45.135 90.935 45.305 ;
      RECT 90.765 47.855 90.935 48.025 ;
      RECT 90.765 50.575 90.935 50.745 ;
      RECT 90.765 53.295 90.935 53.465 ;
      RECT 90.765 56.015 90.935 56.185 ;
      RECT 90.765 58.735 90.935 58.905 ;
      RECT 90.305 9.775 90.475 9.945 ;
      RECT 90.305 12.495 90.475 12.665 ;
      RECT 90.305 15.215 90.475 15.385 ;
      RECT 90.305 17.935 90.475 18.105 ;
      RECT 90.305 20.655 90.475 20.825 ;
      RECT 90.305 23.375 90.475 23.545 ;
      RECT 90.305 26.095 90.475 26.265 ;
      RECT 90.305 28.815 90.475 28.985 ;
      RECT 90.305 31.535 90.475 31.705 ;
      RECT 90.305 34.255 90.475 34.425 ;
      RECT 90.305 36.975 90.475 37.145 ;
      RECT 90.305 39.695 90.475 39.865 ;
      RECT 90.305 42.415 90.475 42.585 ;
      RECT 90.305 45.135 90.475 45.305 ;
      RECT 90.305 47.855 90.475 48.025 ;
      RECT 90.305 50.575 90.475 50.745 ;
      RECT 90.305 53.295 90.475 53.465 ;
      RECT 90.305 56.015 90.475 56.185 ;
      RECT 90.305 58.735 90.475 58.905 ;
      RECT 89.845 9.775 90.015 9.945 ;
      RECT 89.845 12.495 90.015 12.665 ;
      RECT 89.845 15.215 90.015 15.385 ;
      RECT 89.845 17.935 90.015 18.105 ;
      RECT 89.845 20.655 90.015 20.825 ;
      RECT 89.845 23.375 90.015 23.545 ;
      RECT 89.845 26.095 90.015 26.265 ;
      RECT 89.845 28.815 90.015 28.985 ;
      RECT 89.845 31.535 90.015 31.705 ;
      RECT 89.845 34.255 90.015 34.425 ;
      RECT 89.845 36.975 90.015 37.145 ;
      RECT 89.845 39.695 90.015 39.865 ;
      RECT 89.845 42.415 90.015 42.585 ;
      RECT 89.845 45.135 90.015 45.305 ;
      RECT 89.845 47.855 90.015 48.025 ;
      RECT 89.845 50.575 90.015 50.745 ;
      RECT 89.845 53.295 90.015 53.465 ;
      RECT 89.845 56.015 90.015 56.185 ;
      RECT 89.845 58.735 90.015 58.905 ;
      RECT 89.385 9.775 89.555 9.945 ;
      RECT 89.385 12.495 89.555 12.665 ;
      RECT 89.385 15.215 89.555 15.385 ;
      RECT 89.385 17.935 89.555 18.105 ;
      RECT 89.385 20.655 89.555 20.825 ;
      RECT 89.385 23.375 89.555 23.545 ;
      RECT 89.385 26.095 89.555 26.265 ;
      RECT 89.385 28.815 89.555 28.985 ;
      RECT 89.385 31.535 89.555 31.705 ;
      RECT 89.385 34.255 89.555 34.425 ;
      RECT 89.385 36.975 89.555 37.145 ;
      RECT 89.385 39.695 89.555 39.865 ;
      RECT 89.385 42.415 89.555 42.585 ;
      RECT 89.385 45.135 89.555 45.305 ;
      RECT 89.385 47.855 89.555 48.025 ;
      RECT 89.385 50.575 89.555 50.745 ;
      RECT 89.385 53.295 89.555 53.465 ;
      RECT 89.385 56.015 89.555 56.185 ;
      RECT 89.385 58.735 89.555 58.905 ;
      RECT 88.925 9.775 89.095 9.945 ;
      RECT 88.925 12.495 89.095 12.665 ;
      RECT 88.925 15.215 89.095 15.385 ;
      RECT 88.925 17.935 89.095 18.105 ;
      RECT 88.925 20.655 89.095 20.825 ;
      RECT 88.925 23.375 89.095 23.545 ;
      RECT 88.925 26.095 89.095 26.265 ;
      RECT 88.925 28.815 89.095 28.985 ;
      RECT 88.925 31.535 89.095 31.705 ;
      RECT 88.925 34.255 89.095 34.425 ;
      RECT 88.925 36.975 89.095 37.145 ;
      RECT 88.925 39.695 89.095 39.865 ;
      RECT 88.925 42.415 89.095 42.585 ;
      RECT 88.925 45.135 89.095 45.305 ;
      RECT 88.925 47.855 89.095 48.025 ;
      RECT 88.925 50.575 89.095 50.745 ;
      RECT 88.925 53.295 89.095 53.465 ;
      RECT 88.925 56.015 89.095 56.185 ;
      RECT 88.925 58.735 89.095 58.905 ;
      RECT 88.465 9.775 88.635 9.945 ;
      RECT 88.465 12.495 88.635 12.665 ;
      RECT 88.465 15.215 88.635 15.385 ;
      RECT 88.465 17.935 88.635 18.105 ;
      RECT 88.465 20.655 88.635 20.825 ;
      RECT 88.465 23.375 88.635 23.545 ;
      RECT 88.465 26.095 88.635 26.265 ;
      RECT 88.465 28.815 88.635 28.985 ;
      RECT 88.465 31.535 88.635 31.705 ;
      RECT 88.465 34.255 88.635 34.425 ;
      RECT 88.465 36.975 88.635 37.145 ;
      RECT 88.465 39.695 88.635 39.865 ;
      RECT 88.465 42.415 88.635 42.585 ;
      RECT 88.465 45.135 88.635 45.305 ;
      RECT 88.465 47.855 88.635 48.025 ;
      RECT 88.465 50.575 88.635 50.745 ;
      RECT 88.465 53.295 88.635 53.465 ;
      RECT 88.465 56.015 88.635 56.185 ;
      RECT 88.465 58.735 88.635 58.905 ;
      RECT 88.005 9.775 88.175 9.945 ;
      RECT 88.005 12.495 88.175 12.665 ;
      RECT 88.005 15.215 88.175 15.385 ;
      RECT 88.005 15.725 88.175 15.895 ;
      RECT 88.005 17.935 88.175 18.105 ;
      RECT 88.005 20.655 88.175 20.825 ;
      RECT 88.005 23.375 88.175 23.545 ;
      RECT 88.005 26.095 88.175 26.265 ;
      RECT 88.005 28.815 88.175 28.985 ;
      RECT 88.005 31.535 88.175 31.705 ;
      RECT 88.005 34.255 88.175 34.425 ;
      RECT 88.005 36.975 88.175 37.145 ;
      RECT 88.005 39.695 88.175 39.865 ;
      RECT 88.005 42.415 88.175 42.585 ;
      RECT 88.005 45.135 88.175 45.305 ;
      RECT 88.005 47.855 88.175 48.025 ;
      RECT 88.005 50.575 88.175 50.745 ;
      RECT 88.005 53.295 88.175 53.465 ;
      RECT 88.005 56.015 88.175 56.185 ;
      RECT 88.005 58.735 88.175 58.905 ;
      RECT 87.545 9.775 87.715 9.945 ;
      RECT 87.545 12.495 87.715 12.665 ;
      RECT 87.545 15.215 87.715 15.385 ;
      RECT 87.545 17.935 87.715 18.105 ;
      RECT 87.545 20.655 87.715 20.825 ;
      RECT 87.545 23.375 87.715 23.545 ;
      RECT 87.545 26.095 87.715 26.265 ;
      RECT 87.545 28.815 87.715 28.985 ;
      RECT 87.545 31.535 87.715 31.705 ;
      RECT 87.545 34.255 87.715 34.425 ;
      RECT 87.545 36.975 87.715 37.145 ;
      RECT 87.545 39.695 87.715 39.865 ;
      RECT 87.545 42.415 87.715 42.585 ;
      RECT 87.545 45.135 87.715 45.305 ;
      RECT 87.545 47.855 87.715 48.025 ;
      RECT 87.545 50.575 87.715 50.745 ;
      RECT 87.545 53.295 87.715 53.465 ;
      RECT 87.545 56.015 87.715 56.185 ;
      RECT 87.545 58.735 87.715 58.905 ;
      RECT 87.085 9.775 87.255 9.945 ;
      RECT 87.085 12.495 87.255 12.665 ;
      RECT 87.085 15.215 87.255 15.385 ;
      RECT 87.085 17.935 87.255 18.105 ;
      RECT 87.085 20.655 87.255 20.825 ;
      RECT 87.085 23.375 87.255 23.545 ;
      RECT 87.085 26.095 87.255 26.265 ;
      RECT 87.085 28.815 87.255 28.985 ;
      RECT 87.085 31.535 87.255 31.705 ;
      RECT 87.085 34.255 87.255 34.425 ;
      RECT 87.085 36.975 87.255 37.145 ;
      RECT 87.085 39.695 87.255 39.865 ;
      RECT 87.085 42.415 87.255 42.585 ;
      RECT 87.085 45.135 87.255 45.305 ;
      RECT 87.085 47.855 87.255 48.025 ;
      RECT 87.085 50.575 87.255 50.745 ;
      RECT 87.085 53.295 87.255 53.465 ;
      RECT 87.085 56.015 87.255 56.185 ;
      RECT 87.085 58.735 87.255 58.905 ;
      RECT 86.625 9.775 86.795 9.945 ;
      RECT 86.625 12.495 86.795 12.665 ;
      RECT 86.625 15.215 86.795 15.385 ;
      RECT 86.625 17.935 86.795 18.105 ;
      RECT 86.625 19.125 86.795 19.295 ;
      RECT 86.625 20.655 86.795 20.825 ;
      RECT 86.625 22.185 86.795 22.355 ;
      RECT 86.625 23.375 86.795 23.545 ;
      RECT 86.625 26.095 86.795 26.265 ;
      RECT 86.625 28.815 86.795 28.985 ;
      RECT 86.625 31.535 86.795 31.705 ;
      RECT 86.625 34.255 86.795 34.425 ;
      RECT 86.625 36.975 86.795 37.145 ;
      RECT 86.625 39.695 86.795 39.865 ;
      RECT 86.625 42.415 86.795 42.585 ;
      RECT 86.625 45.135 86.795 45.305 ;
      RECT 86.625 47.855 86.795 48.025 ;
      RECT 86.625 50.575 86.795 50.745 ;
      RECT 86.625 53.295 86.795 53.465 ;
      RECT 86.625 56.015 86.795 56.185 ;
      RECT 86.625 58.735 86.795 58.905 ;
      RECT 86.165 9.775 86.335 9.945 ;
      RECT 86.165 12.495 86.335 12.665 ;
      RECT 86.165 15.215 86.335 15.385 ;
      RECT 86.165 17.935 86.335 18.105 ;
      RECT 86.165 20.655 86.335 20.825 ;
      RECT 86.165 23.375 86.335 23.545 ;
      RECT 86.165 26.095 86.335 26.265 ;
      RECT 86.165 28.815 86.335 28.985 ;
      RECT 86.165 31.535 86.335 31.705 ;
      RECT 86.165 34.255 86.335 34.425 ;
      RECT 86.165 36.975 86.335 37.145 ;
      RECT 86.165 39.695 86.335 39.865 ;
      RECT 86.165 42.415 86.335 42.585 ;
      RECT 86.165 45.135 86.335 45.305 ;
      RECT 86.165 47.855 86.335 48.025 ;
      RECT 86.165 50.575 86.335 50.745 ;
      RECT 86.165 53.295 86.335 53.465 ;
      RECT 86.165 56.015 86.335 56.185 ;
      RECT 86.165 58.735 86.335 58.905 ;
      RECT 86.02 19.125 86.19 19.295 ;
      RECT 85.705 9.775 85.875 9.945 ;
      RECT 85.705 12.495 85.875 12.665 ;
      RECT 85.705 15.215 85.875 15.385 ;
      RECT 85.705 17.935 85.875 18.105 ;
      RECT 85.705 20.655 85.875 20.825 ;
      RECT 85.705 23.375 85.875 23.545 ;
      RECT 85.705 26.095 85.875 26.265 ;
      RECT 85.705 28.815 85.875 28.985 ;
      RECT 85.705 31.535 85.875 31.705 ;
      RECT 85.705 34.255 85.875 34.425 ;
      RECT 85.705 36.975 85.875 37.145 ;
      RECT 85.705 39.695 85.875 39.865 ;
      RECT 85.705 42.415 85.875 42.585 ;
      RECT 85.705 45.135 85.875 45.305 ;
      RECT 85.705 47.855 85.875 48.025 ;
      RECT 85.705 50.575 85.875 50.745 ;
      RECT 85.705 53.295 85.875 53.465 ;
      RECT 85.705 56.015 85.875 56.185 ;
      RECT 85.705 58.735 85.875 58.905 ;
      RECT 85.695 16.405 85.865 16.575 ;
      RECT 85.26 16.065 85.43 16.235 ;
      RECT 85.245 9.775 85.415 9.945 ;
      RECT 85.245 12.495 85.415 12.665 ;
      RECT 85.245 15.215 85.415 15.385 ;
      RECT 85.245 17.935 85.415 18.105 ;
      RECT 85.245 18.785 85.415 18.955 ;
      RECT 85.245 20.655 85.415 20.825 ;
      RECT 85.245 23.375 85.415 23.545 ;
      RECT 85.245 24.565 85.415 24.735 ;
      RECT 85.245 26.095 85.415 26.265 ;
      RECT 85.245 28.815 85.415 28.985 ;
      RECT 85.245 31.535 85.415 31.705 ;
      RECT 85.245 34.255 85.415 34.425 ;
      RECT 85.245 36.975 85.415 37.145 ;
      RECT 85.245 39.695 85.415 39.865 ;
      RECT 85.245 42.415 85.415 42.585 ;
      RECT 85.245 45.135 85.415 45.305 ;
      RECT 85.245 47.855 85.415 48.025 ;
      RECT 85.245 50.575 85.415 50.745 ;
      RECT 85.245 53.295 85.415 53.465 ;
      RECT 85.245 56.015 85.415 56.185 ;
      RECT 85.245 58.735 85.415 58.905 ;
      RECT 84.785 9.775 84.955 9.945 ;
      RECT 84.785 12.495 84.955 12.665 ;
      RECT 84.785 15.215 84.955 15.385 ;
      RECT 84.785 17.935 84.955 18.105 ;
      RECT 84.785 19.125 84.955 19.295 ;
      RECT 84.785 20.655 84.955 20.825 ;
      RECT 84.785 23.375 84.955 23.545 ;
      RECT 84.785 26.095 84.955 26.265 ;
      RECT 84.785 26.605 84.955 26.775 ;
      RECT 84.785 28.815 84.955 28.985 ;
      RECT 84.785 31.535 84.955 31.705 ;
      RECT 84.785 34.255 84.955 34.425 ;
      RECT 84.785 36.975 84.955 37.145 ;
      RECT 84.785 39.695 84.955 39.865 ;
      RECT 84.785 42.415 84.955 42.585 ;
      RECT 84.785 45.135 84.955 45.305 ;
      RECT 84.785 47.855 84.955 48.025 ;
      RECT 84.785 50.575 84.955 50.745 ;
      RECT 84.785 53.295 84.955 53.465 ;
      RECT 84.785 56.015 84.955 56.185 ;
      RECT 84.785 58.735 84.955 58.905 ;
      RECT 84.555 24.565 84.725 24.735 ;
      RECT 84.325 9.775 84.495 9.945 ;
      RECT 84.325 12.495 84.495 12.665 ;
      RECT 84.325 15.215 84.495 15.385 ;
      RECT 84.325 17.935 84.495 18.105 ;
      RECT 84.325 20.655 84.495 20.825 ;
      RECT 84.325 23.375 84.495 23.545 ;
      RECT 84.325 26.095 84.495 26.265 ;
      RECT 84.325 28.815 84.495 28.985 ;
      RECT 84.325 31.535 84.495 31.705 ;
      RECT 84.325 34.255 84.495 34.425 ;
      RECT 84.325 36.975 84.495 37.145 ;
      RECT 84.325 39.695 84.495 39.865 ;
      RECT 84.325 42.415 84.495 42.585 ;
      RECT 84.325 45.135 84.495 45.305 ;
      RECT 84.325 47.855 84.495 48.025 ;
      RECT 84.325 50.575 84.495 50.745 ;
      RECT 84.325 53.295 84.495 53.465 ;
      RECT 84.325 56.015 84.495 56.185 ;
      RECT 84.325 58.735 84.495 58.905 ;
      RECT 84.095 19.125 84.265 19.295 ;
      RECT 83.865 9.775 84.035 9.945 ;
      RECT 83.865 12.495 84.035 12.665 ;
      RECT 83.865 15.215 84.035 15.385 ;
      RECT 83.865 17.935 84.035 18.105 ;
      RECT 83.865 20.655 84.035 20.825 ;
      RECT 83.865 23.375 84.035 23.545 ;
      RECT 83.865 24.225 84.035 24.395 ;
      RECT 83.865 26.095 84.035 26.265 ;
      RECT 83.865 28.815 84.035 28.985 ;
      RECT 83.865 31.535 84.035 31.705 ;
      RECT 83.865 34.255 84.035 34.425 ;
      RECT 83.865 36.975 84.035 37.145 ;
      RECT 83.865 39.695 84.035 39.865 ;
      RECT 83.865 42.415 84.035 42.585 ;
      RECT 83.865 45.135 84.035 45.305 ;
      RECT 83.865 47.855 84.035 48.025 ;
      RECT 83.865 50.575 84.035 50.745 ;
      RECT 83.865 53.295 84.035 53.465 ;
      RECT 83.865 56.015 84.035 56.185 ;
      RECT 83.865 58.735 84.035 58.905 ;
      RECT 83.69 16.065 83.86 16.235 ;
      RECT 83.405 9.775 83.575 9.945 ;
      RECT 83.405 11.305 83.575 11.475 ;
      RECT 83.405 12.495 83.575 12.665 ;
      RECT 83.405 15.215 83.575 15.385 ;
      RECT 83.405 17.935 83.575 18.105 ;
      RECT 83.405 19.805 83.575 19.975 ;
      RECT 83.405 20.655 83.575 20.825 ;
      RECT 83.405 23.375 83.575 23.545 ;
      RECT 83.405 24.565 83.575 24.735 ;
      RECT 83.405 26.095 83.575 26.265 ;
      RECT 83.405 28.815 83.575 28.985 ;
      RECT 83.405 31.535 83.575 31.705 ;
      RECT 83.405 34.255 83.575 34.425 ;
      RECT 83.405 36.975 83.575 37.145 ;
      RECT 83.405 39.695 83.575 39.865 ;
      RECT 83.405 42.415 83.575 42.585 ;
      RECT 83.405 45.135 83.575 45.305 ;
      RECT 83.405 47.855 83.575 48.025 ;
      RECT 83.405 50.575 83.575 50.745 ;
      RECT 83.405 53.295 83.575 53.465 ;
      RECT 83.405 56.015 83.575 56.185 ;
      RECT 83.405 58.735 83.575 58.905 ;
      RECT 83.175 16.405 83.345 16.575 ;
      RECT 82.945 9.775 83.115 9.945 ;
      RECT 82.945 12.495 83.115 12.665 ;
      RECT 82.945 15.215 83.115 15.385 ;
      RECT 82.945 17.935 83.115 18.105 ;
      RECT 82.945 20.655 83.115 20.825 ;
      RECT 82.945 23.375 83.115 23.545 ;
      RECT 82.945 26.095 83.115 26.265 ;
      RECT 82.945 28.815 83.115 28.985 ;
      RECT 82.945 31.535 83.115 31.705 ;
      RECT 82.945 34.255 83.115 34.425 ;
      RECT 82.945 36.975 83.115 37.145 ;
      RECT 82.945 39.695 83.115 39.865 ;
      RECT 82.945 42.415 83.115 42.585 ;
      RECT 82.945 45.135 83.115 45.305 ;
      RECT 82.945 47.855 83.115 48.025 ;
      RECT 82.945 50.575 83.115 50.745 ;
      RECT 82.945 53.295 83.115 53.465 ;
      RECT 82.945 56.015 83.115 56.185 ;
      RECT 82.945 58.735 83.115 58.905 ;
      RECT 82.715 24.565 82.885 24.735 ;
      RECT 82.485 9.775 82.655 9.945 ;
      RECT 82.485 12.495 82.655 12.665 ;
      RECT 82.485 15.215 82.655 15.385 ;
      RECT 82.485 17.935 82.655 18.105 ;
      RECT 82.485 20.655 82.655 20.825 ;
      RECT 82.485 23.375 82.655 23.545 ;
      RECT 82.485 26.095 82.655 26.265 ;
      RECT 82.485 28.815 82.655 28.985 ;
      RECT 82.485 31.535 82.655 31.705 ;
      RECT 82.485 34.255 82.655 34.425 ;
      RECT 82.485 36.975 82.655 37.145 ;
      RECT 82.485 39.695 82.655 39.865 ;
      RECT 82.485 42.415 82.655 42.585 ;
      RECT 82.485 45.135 82.655 45.305 ;
      RECT 82.485 47.855 82.655 48.025 ;
      RECT 82.485 50.575 82.655 50.745 ;
      RECT 82.485 53.295 82.655 53.465 ;
      RECT 82.485 56.015 82.655 56.185 ;
      RECT 82.485 58.735 82.655 58.905 ;
      RECT 82.475 27.285 82.645 27.455 ;
      RECT 82.41 17.085 82.58 17.255 ;
      RECT 82.04 26.945 82.21 27.115 ;
      RECT 82.025 9.775 82.195 9.945 ;
      RECT 82.025 12.495 82.195 12.665 ;
      RECT 82.025 15.215 82.195 15.385 ;
      RECT 82.025 17.935 82.195 18.105 ;
      RECT 82.025 20.655 82.195 20.825 ;
      RECT 82.025 23.375 82.195 23.545 ;
      RECT 82.025 25.585 82.195 25.755 ;
      RECT 82.025 26.095 82.195 26.265 ;
      RECT 82.025 28.815 82.195 28.985 ;
      RECT 82.025 31.535 82.195 31.705 ;
      RECT 82.025 33.745 82.195 33.915 ;
      RECT 82.025 34.255 82.195 34.425 ;
      RECT 82.025 36.975 82.195 37.145 ;
      RECT 82.025 39.695 82.195 39.865 ;
      RECT 82.025 42.415 82.195 42.585 ;
      RECT 82.025 45.135 82.195 45.305 ;
      RECT 82.025 47.855 82.195 48.025 ;
      RECT 82.025 50.575 82.195 50.745 ;
      RECT 82.025 53.295 82.195 53.465 ;
      RECT 82.025 56.015 82.195 56.185 ;
      RECT 82.025 58.735 82.195 58.905 ;
      RECT 81.985 16.405 82.155 16.575 ;
      RECT 81.59 16.065 81.76 16.235 ;
      RECT 81.565 9.775 81.735 9.945 ;
      RECT 81.565 12.495 81.735 12.665 ;
      RECT 81.565 15.215 81.735 15.385 ;
      RECT 81.565 17.935 81.735 18.105 ;
      RECT 81.565 20.655 81.735 20.825 ;
      RECT 81.565 23.375 81.735 23.545 ;
      RECT 81.565 26.095 81.735 26.265 ;
      RECT 81.565 28.815 81.735 28.985 ;
      RECT 81.565 31.535 81.735 31.705 ;
      RECT 81.565 34.255 81.735 34.425 ;
      RECT 81.565 36.975 81.735 37.145 ;
      RECT 81.565 39.695 81.735 39.865 ;
      RECT 81.565 42.415 81.735 42.585 ;
      RECT 81.565 45.135 81.735 45.305 ;
      RECT 81.565 47.855 81.735 48.025 ;
      RECT 81.565 50.575 81.735 50.745 ;
      RECT 81.565 53.295 81.735 53.465 ;
      RECT 81.565 56.015 81.735 56.185 ;
      RECT 81.565 58.735 81.735 58.905 ;
      RECT 81.105 9.775 81.275 9.945 ;
      RECT 81.105 12.495 81.275 12.665 ;
      RECT 81.105 15.215 81.275 15.385 ;
      RECT 81.105 16.745 81.275 16.915 ;
      RECT 81.105 17.935 81.275 18.105 ;
      RECT 81.105 18.445 81.275 18.615 ;
      RECT 81.105 20.655 81.275 20.825 ;
      RECT 81.105 23.375 81.275 23.545 ;
      RECT 81.105 26.095 81.275 26.265 ;
      RECT 81.105 28.815 81.275 28.985 ;
      RECT 81.105 31.535 81.275 31.705 ;
      RECT 81.105 34.255 81.275 34.425 ;
      RECT 81.105 36.975 81.275 37.145 ;
      RECT 81.105 39.695 81.275 39.865 ;
      RECT 81.105 42.415 81.275 42.585 ;
      RECT 81.105 45.135 81.275 45.305 ;
      RECT 81.105 47.855 81.275 48.025 ;
      RECT 81.105 50.575 81.275 50.745 ;
      RECT 81.105 53.295 81.275 53.465 ;
      RECT 81.105 56.015 81.275 56.185 ;
      RECT 81.105 58.735 81.275 58.905 ;
      RECT 80.645 9.775 80.815 9.945 ;
      RECT 80.645 12.495 80.815 12.665 ;
      RECT 80.645 15.215 80.815 15.385 ;
      RECT 80.645 17.935 80.815 18.105 ;
      RECT 80.645 20.655 80.815 20.825 ;
      RECT 80.645 23.375 80.815 23.545 ;
      RECT 80.645 26.095 80.815 26.265 ;
      RECT 80.645 28.815 80.815 28.985 ;
      RECT 80.645 31.535 80.815 31.705 ;
      RECT 80.645 34.255 80.815 34.425 ;
      RECT 80.645 36.975 80.815 37.145 ;
      RECT 80.645 39.695 80.815 39.865 ;
      RECT 80.645 42.415 80.815 42.585 ;
      RECT 80.645 45.135 80.815 45.305 ;
      RECT 80.645 47.855 80.815 48.025 ;
      RECT 80.645 50.575 80.815 50.745 ;
      RECT 80.645 53.295 80.815 53.465 ;
      RECT 80.645 56.015 80.815 56.185 ;
      RECT 80.645 58.735 80.815 58.905 ;
      RECT 80.47 26.945 80.64 27.115 ;
      RECT 80.185 9.775 80.355 9.945 ;
      RECT 80.185 12.495 80.355 12.665 ;
      RECT 80.185 15.215 80.355 15.385 ;
      RECT 80.185 17.935 80.355 18.105 ;
      RECT 80.185 20.655 80.355 20.825 ;
      RECT 80.185 23.375 80.355 23.545 ;
      RECT 80.185 26.095 80.355 26.265 ;
      RECT 80.185 28.815 80.355 28.985 ;
      RECT 80.185 31.535 80.355 31.705 ;
      RECT 80.185 34.255 80.355 34.425 ;
      RECT 80.185 36.975 80.355 37.145 ;
      RECT 80.185 39.695 80.355 39.865 ;
      RECT 80.185 42.415 80.355 42.585 ;
      RECT 80.185 45.135 80.355 45.305 ;
      RECT 80.185 47.855 80.355 48.025 ;
      RECT 80.185 50.575 80.355 50.745 ;
      RECT 80.185 53.295 80.355 53.465 ;
      RECT 80.185 56.015 80.355 56.185 ;
      RECT 80.185 58.735 80.355 58.905 ;
      RECT 79.955 27.285 80.125 27.455 ;
      RECT 79.725 9.775 79.895 9.945 ;
      RECT 79.725 12.495 79.895 12.665 ;
      RECT 79.725 15.215 79.895 15.385 ;
      RECT 79.725 17.935 79.895 18.105 ;
      RECT 79.725 20.655 79.895 20.825 ;
      RECT 79.725 23.375 79.895 23.545 ;
      RECT 79.725 26.095 79.895 26.265 ;
      RECT 79.725 28.815 79.895 28.985 ;
      RECT 79.725 31.535 79.895 31.705 ;
      RECT 79.725 34.255 79.895 34.425 ;
      RECT 79.725 36.975 79.895 37.145 ;
      RECT 79.725 39.695 79.895 39.865 ;
      RECT 79.725 42.415 79.895 42.585 ;
      RECT 79.725 45.135 79.895 45.305 ;
      RECT 79.725 47.855 79.895 48.025 ;
      RECT 79.725 50.575 79.895 50.745 ;
      RECT 79.725 53.295 79.895 53.465 ;
      RECT 79.725 56.015 79.895 56.185 ;
      RECT 79.725 58.735 79.895 58.905 ;
      RECT 79.715 32.725 79.885 32.895 ;
      RECT 79.28 32.385 79.45 32.555 ;
      RECT 79.265 9.775 79.435 9.945 ;
      RECT 79.265 12.495 79.435 12.665 ;
      RECT 79.265 15.215 79.435 15.385 ;
      RECT 79.265 17.935 79.435 18.105 ;
      RECT 79.265 20.655 79.435 20.825 ;
      RECT 79.265 23.375 79.435 23.545 ;
      RECT 79.265 26.095 79.435 26.265 ;
      RECT 79.265 28.815 79.435 28.985 ;
      RECT 79.265 31.535 79.435 31.705 ;
      RECT 79.265 34.255 79.435 34.425 ;
      RECT 79.265 36.975 79.435 37.145 ;
      RECT 79.265 39.695 79.435 39.865 ;
      RECT 79.265 42.415 79.435 42.585 ;
      RECT 79.265 45.135 79.435 45.305 ;
      RECT 79.265 47.855 79.435 48.025 ;
      RECT 79.265 50.575 79.435 50.745 ;
      RECT 79.265 53.295 79.435 53.465 ;
      RECT 79.265 56.015 79.435 56.185 ;
      RECT 79.265 58.735 79.435 58.905 ;
      RECT 79.19 27.625 79.36 27.795 ;
      RECT 78.805 9.775 78.975 9.945 ;
      RECT 78.805 12.495 78.975 12.665 ;
      RECT 78.805 15.215 78.975 15.385 ;
      RECT 78.805 17.935 78.975 18.105 ;
      RECT 78.805 20.655 78.975 20.825 ;
      RECT 78.805 23.375 78.975 23.545 ;
      RECT 78.805 24.565 78.975 24.735 ;
      RECT 78.805 26.095 78.975 26.265 ;
      RECT 78.805 28.815 78.975 28.985 ;
      RECT 78.805 31.535 78.975 31.705 ;
      RECT 78.805 34.255 78.975 34.425 ;
      RECT 78.805 36.975 78.975 37.145 ;
      RECT 78.805 39.695 78.975 39.865 ;
      RECT 78.805 42.415 78.975 42.585 ;
      RECT 78.805 45.135 78.975 45.305 ;
      RECT 78.805 47.855 78.975 48.025 ;
      RECT 78.805 50.575 78.975 50.745 ;
      RECT 78.805 53.295 78.975 53.465 ;
      RECT 78.805 56.015 78.975 56.185 ;
      RECT 78.805 58.735 78.975 58.905 ;
      RECT 78.795 19.465 78.965 19.635 ;
      RECT 78.765 27.285 78.935 27.455 ;
      RECT 78.37 26.945 78.54 27.115 ;
      RECT 78.36 19.805 78.53 19.975 ;
      RECT 78.345 9.775 78.515 9.945 ;
      RECT 78.345 11.305 78.515 11.475 ;
      RECT 78.345 12.495 78.515 12.665 ;
      RECT 78.345 15.215 78.515 15.385 ;
      RECT 78.345 17.935 78.515 18.105 ;
      RECT 78.345 20.655 78.515 20.825 ;
      RECT 78.345 23.375 78.515 23.545 ;
      RECT 78.345 26.095 78.515 26.265 ;
      RECT 78.345 28.815 78.515 28.985 ;
      RECT 78.345 31.535 78.515 31.705 ;
      RECT 78.345 34.255 78.515 34.425 ;
      RECT 78.345 36.975 78.515 37.145 ;
      RECT 78.345 39.695 78.515 39.865 ;
      RECT 78.345 42.415 78.515 42.585 ;
      RECT 78.345 45.135 78.515 45.305 ;
      RECT 78.345 47.855 78.515 48.025 ;
      RECT 78.345 50.575 78.515 50.745 ;
      RECT 78.345 53.295 78.515 53.465 ;
      RECT 78.345 56.015 78.515 56.185 ;
      RECT 78.345 58.735 78.515 58.905 ;
      RECT 78.115 24.565 78.285 24.735 ;
      RECT 77.885 9.775 78.055 9.945 ;
      RECT 77.885 12.495 78.055 12.665 ;
      RECT 77.885 15.215 78.055 15.385 ;
      RECT 77.885 17.935 78.055 18.105 ;
      RECT 77.885 20.655 78.055 20.825 ;
      RECT 77.885 23.375 78.055 23.545 ;
      RECT 77.885 26.095 78.055 26.265 ;
      RECT 77.885 27.285 78.055 27.455 ;
      RECT 77.885 28.815 78.055 28.985 ;
      RECT 77.885 31.535 78.055 31.705 ;
      RECT 77.885 34.255 78.055 34.425 ;
      RECT 77.885 36.975 78.055 37.145 ;
      RECT 77.885 39.695 78.055 39.865 ;
      RECT 77.885 42.415 78.055 42.585 ;
      RECT 77.885 45.135 78.055 45.305 ;
      RECT 77.885 47.855 78.055 48.025 ;
      RECT 77.885 50.575 78.055 50.745 ;
      RECT 77.885 53.295 78.055 53.465 ;
      RECT 77.885 56.015 78.055 56.185 ;
      RECT 77.885 58.735 78.055 58.905 ;
      RECT 77.71 32.385 77.88 32.555 ;
      RECT 77.425 9.775 77.595 9.945 ;
      RECT 77.425 12.495 77.595 12.665 ;
      RECT 77.425 15.215 77.595 15.385 ;
      RECT 77.425 17.935 77.595 18.105 ;
      RECT 77.425 20.655 77.595 20.825 ;
      RECT 77.425 23.375 77.595 23.545 ;
      RECT 77.425 24.225 77.595 24.395 ;
      RECT 77.425 26.095 77.595 26.265 ;
      RECT 77.425 28.815 77.595 28.985 ;
      RECT 77.425 31.535 77.595 31.705 ;
      RECT 77.425 34.255 77.595 34.425 ;
      RECT 77.425 36.975 77.595 37.145 ;
      RECT 77.425 39.695 77.595 39.865 ;
      RECT 77.425 42.415 77.595 42.585 ;
      RECT 77.425 45.135 77.595 45.305 ;
      RECT 77.425 47.855 77.595 48.025 ;
      RECT 77.425 50.575 77.595 50.745 ;
      RECT 77.425 53.295 77.595 53.465 ;
      RECT 77.425 56.015 77.595 56.185 ;
      RECT 77.425 58.735 77.595 58.905 ;
      RECT 77.195 32.725 77.365 32.895 ;
      RECT 76.965 9.775 77.135 9.945 ;
      RECT 76.965 12.495 77.135 12.665 ;
      RECT 76.965 15.215 77.135 15.385 ;
      RECT 76.965 17.935 77.135 18.105 ;
      RECT 76.965 20.655 77.135 20.825 ;
      RECT 76.965 23.375 77.135 23.545 ;
      RECT 76.965 24.565 77.135 24.735 ;
      RECT 76.965 26.095 77.135 26.265 ;
      RECT 76.965 28.815 77.135 28.985 ;
      RECT 76.965 31.535 77.135 31.705 ;
      RECT 76.965 34.255 77.135 34.425 ;
      RECT 76.965 36.975 77.135 37.145 ;
      RECT 76.965 39.695 77.135 39.865 ;
      RECT 76.965 42.415 77.135 42.585 ;
      RECT 76.965 45.135 77.135 45.305 ;
      RECT 76.965 47.855 77.135 48.025 ;
      RECT 76.965 50.575 77.135 50.745 ;
      RECT 76.965 53.295 77.135 53.465 ;
      RECT 76.965 56.015 77.135 56.185 ;
      RECT 76.965 58.735 77.135 58.905 ;
      RECT 76.79 19.805 76.96 19.975 ;
      RECT 76.505 9.775 76.675 9.945 ;
      RECT 76.505 12.495 76.675 12.665 ;
      RECT 76.505 15.215 76.675 15.385 ;
      RECT 76.505 17.935 76.675 18.105 ;
      RECT 76.505 20.655 76.675 20.825 ;
      RECT 76.505 23.375 76.675 23.545 ;
      RECT 76.505 26.095 76.675 26.265 ;
      RECT 76.505 28.815 76.675 28.985 ;
      RECT 76.505 31.535 76.675 31.705 ;
      RECT 76.505 34.255 76.675 34.425 ;
      RECT 76.505 36.975 76.675 37.145 ;
      RECT 76.505 39.695 76.675 39.865 ;
      RECT 76.505 42.415 76.675 42.585 ;
      RECT 76.505 45.135 76.675 45.305 ;
      RECT 76.505 47.855 76.675 48.025 ;
      RECT 76.505 50.575 76.675 50.745 ;
      RECT 76.505 53.295 76.675 53.465 ;
      RECT 76.505 56.015 76.675 56.185 ;
      RECT 76.505 58.735 76.675 58.905 ;
      RECT 76.43 24.565 76.6 24.735 ;
      RECT 76.43 33.405 76.6 33.575 ;
      RECT 76.275 19.465 76.445 19.635 ;
      RECT 76.045 9.775 76.215 9.945 ;
      RECT 76.045 12.495 76.215 12.665 ;
      RECT 76.045 15.215 76.215 15.385 ;
      RECT 76.045 17.935 76.215 18.105 ;
      RECT 76.045 20.655 76.215 20.825 ;
      RECT 76.045 23.375 76.215 23.545 ;
      RECT 76.045 26.095 76.215 26.265 ;
      RECT 76.045 28.815 76.215 28.985 ;
      RECT 76.045 31.535 76.215 31.705 ;
      RECT 76.045 34.255 76.215 34.425 ;
      RECT 76.045 36.975 76.215 37.145 ;
      RECT 76.045 39.695 76.215 39.865 ;
      RECT 76.045 42.415 76.215 42.585 ;
      RECT 76.045 45.135 76.215 45.305 ;
      RECT 76.045 47.855 76.215 48.025 ;
      RECT 76.045 50.575 76.215 50.745 ;
      RECT 76.045 53.295 76.215 53.465 ;
      RECT 76.045 56.015 76.215 56.185 ;
      RECT 76.045 58.735 76.215 58.905 ;
      RECT 76.005 32.725 76.175 32.895 ;
      RECT 75.61 32.385 75.78 32.555 ;
      RECT 75.585 9.775 75.755 9.945 ;
      RECT 75.585 12.495 75.755 12.665 ;
      RECT 75.585 15.215 75.755 15.385 ;
      RECT 75.585 17.935 75.755 18.105 ;
      RECT 75.585 20.655 75.755 20.825 ;
      RECT 75.585 23.375 75.755 23.545 ;
      RECT 75.585 25.585 75.755 25.755 ;
      RECT 75.585 26.095 75.755 26.265 ;
      RECT 75.585 28.815 75.755 28.985 ;
      RECT 75.585 31.535 75.755 31.705 ;
      RECT 75.585 34.255 75.755 34.425 ;
      RECT 75.585 36.975 75.755 37.145 ;
      RECT 75.585 39.695 75.755 39.865 ;
      RECT 75.585 42.415 75.755 42.585 ;
      RECT 75.585 45.135 75.755 45.305 ;
      RECT 75.585 47.855 75.755 48.025 ;
      RECT 75.585 50.575 75.755 50.745 ;
      RECT 75.585 53.295 75.755 53.465 ;
      RECT 75.585 56.015 75.755 56.185 ;
      RECT 75.585 58.735 75.755 58.905 ;
      RECT 75.54 19.135 75.71 19.305 ;
      RECT 75.125 9.775 75.295 9.945 ;
      RECT 75.125 12.495 75.295 12.665 ;
      RECT 75.125 15.215 75.295 15.385 ;
      RECT 75.125 17.935 75.295 18.105 ;
      RECT 75.125 20.655 75.295 20.825 ;
      RECT 75.125 23.375 75.295 23.545 ;
      RECT 75.125 26.095 75.295 26.265 ;
      RECT 75.125 28.815 75.295 28.985 ;
      RECT 75.125 31.535 75.295 31.705 ;
      RECT 75.125 32.725 75.295 32.895 ;
      RECT 75.125 34.255 75.295 34.425 ;
      RECT 75.125 36.975 75.295 37.145 ;
      RECT 75.125 39.695 75.295 39.865 ;
      RECT 75.125 42.415 75.295 42.585 ;
      RECT 75.125 45.135 75.295 45.305 ;
      RECT 75.125 47.855 75.295 48.025 ;
      RECT 75.125 50.575 75.295 50.745 ;
      RECT 75.125 53.295 75.295 53.465 ;
      RECT 75.125 56.015 75.295 56.185 ;
      RECT 75.125 58.735 75.295 58.905 ;
      RECT 75.085 19.465 75.255 19.635 ;
      RECT 74.69 19.805 74.86 19.975 ;
      RECT 74.665 9.775 74.835 9.945 ;
      RECT 74.665 12.495 74.835 12.665 ;
      RECT 74.665 15.215 74.835 15.385 ;
      RECT 74.665 17.935 74.835 18.105 ;
      RECT 74.665 20.655 74.835 20.825 ;
      RECT 74.665 23.375 74.835 23.545 ;
      RECT 74.665 26.095 74.835 26.265 ;
      RECT 74.665 28.815 74.835 28.985 ;
      RECT 74.665 31.535 74.835 31.705 ;
      RECT 74.665 34.255 74.835 34.425 ;
      RECT 74.665 36.975 74.835 37.145 ;
      RECT 74.665 39.695 74.835 39.865 ;
      RECT 74.665 42.415 74.835 42.585 ;
      RECT 74.665 45.135 74.835 45.305 ;
      RECT 74.665 47.855 74.835 48.025 ;
      RECT 74.665 50.575 74.835 50.745 ;
      RECT 74.665 53.295 74.835 53.465 ;
      RECT 74.665 56.015 74.835 56.185 ;
      RECT 74.665 58.735 74.835 58.905 ;
      RECT 74.205 9.775 74.375 9.945 ;
      RECT 74.205 12.495 74.375 12.665 ;
      RECT 74.205 15.215 74.375 15.385 ;
      RECT 74.205 17.935 74.375 18.105 ;
      RECT 74.205 20.655 74.375 20.825 ;
      RECT 74.205 23.375 74.375 23.545 ;
      RECT 74.205 26.095 74.375 26.265 ;
      RECT 74.205 28.815 74.375 28.985 ;
      RECT 74.205 31.535 74.375 31.705 ;
      RECT 74.205 34.255 74.375 34.425 ;
      RECT 74.205 36.975 74.375 37.145 ;
      RECT 74.205 39.695 74.375 39.865 ;
      RECT 74.205 42.415 74.375 42.585 ;
      RECT 74.205 45.135 74.375 45.305 ;
      RECT 74.205 47.855 74.375 48.025 ;
      RECT 74.205 50.575 74.375 50.745 ;
      RECT 74.205 53.295 74.375 53.465 ;
      RECT 74.205 56.015 74.375 56.185 ;
      RECT 74.205 58.735 74.375 58.905 ;
      RECT 73.745 9.775 73.915 9.945 ;
      RECT 73.745 12.495 73.915 12.665 ;
      RECT 73.745 15.215 73.915 15.385 ;
      RECT 73.745 16.745 73.915 16.915 ;
      RECT 73.745 17.935 73.915 18.105 ;
      RECT 73.745 20.655 73.915 20.825 ;
      RECT 73.745 23.375 73.915 23.545 ;
      RECT 73.745 26.095 73.915 26.265 ;
      RECT 73.745 28.815 73.915 28.985 ;
      RECT 73.745 31.535 73.915 31.705 ;
      RECT 73.745 34.255 73.915 34.425 ;
      RECT 73.745 36.975 73.915 37.145 ;
      RECT 73.745 39.695 73.915 39.865 ;
      RECT 73.745 42.415 73.915 42.585 ;
      RECT 73.745 45.135 73.915 45.305 ;
      RECT 73.745 47.855 73.915 48.025 ;
      RECT 73.745 50.575 73.915 50.745 ;
      RECT 73.745 53.295 73.915 53.465 ;
      RECT 73.745 56.015 73.915 56.185 ;
      RECT 73.745 58.735 73.915 58.905 ;
      RECT 73.285 9.775 73.455 9.945 ;
      RECT 73.285 12.495 73.455 12.665 ;
      RECT 73.285 15.215 73.455 15.385 ;
      RECT 73.285 15.725 73.455 15.895 ;
      RECT 73.285 17.935 73.455 18.105 ;
      RECT 73.285 18.785 73.455 18.955 ;
      RECT 73.285 20.655 73.455 20.825 ;
      RECT 73.285 23.375 73.455 23.545 ;
      RECT 73.285 26.095 73.455 26.265 ;
      RECT 73.285 28.815 73.455 28.985 ;
      RECT 73.285 31.535 73.455 31.705 ;
      RECT 73.285 34.255 73.455 34.425 ;
      RECT 73.285 36.975 73.455 37.145 ;
      RECT 73.285 39.695 73.455 39.865 ;
      RECT 73.285 42.415 73.455 42.585 ;
      RECT 73.285 45.135 73.455 45.305 ;
      RECT 73.285 47.855 73.455 48.025 ;
      RECT 73.285 50.575 73.455 50.745 ;
      RECT 73.285 53.295 73.455 53.465 ;
      RECT 73.285 56.015 73.455 56.185 ;
      RECT 73.285 58.735 73.455 58.905 ;
      RECT 72.825 9.775 72.995 9.945 ;
      RECT 72.825 12.495 72.995 12.665 ;
      RECT 72.825 15.215 72.995 15.385 ;
      RECT 72.825 17.935 72.995 18.105 ;
      RECT 72.825 20.655 72.995 20.825 ;
      RECT 72.825 23.375 72.995 23.545 ;
      RECT 72.825 26.095 72.995 26.265 ;
      RECT 72.825 28.815 72.995 28.985 ;
      RECT 72.825 31.535 72.995 31.705 ;
      RECT 72.825 34.255 72.995 34.425 ;
      RECT 72.825 36.975 72.995 37.145 ;
      RECT 72.825 39.695 72.995 39.865 ;
      RECT 72.825 42.415 72.995 42.585 ;
      RECT 72.825 45.135 72.995 45.305 ;
      RECT 72.825 47.855 72.995 48.025 ;
      RECT 72.825 50.575 72.995 50.745 ;
      RECT 72.825 53.295 72.995 53.465 ;
      RECT 72.825 56.015 72.995 56.185 ;
      RECT 72.825 58.735 72.995 58.905 ;
      RECT 72.365 9.775 72.535 9.945 ;
      RECT 72.365 12.495 72.535 12.665 ;
      RECT 72.365 15.215 72.535 15.385 ;
      RECT 72.365 17.935 72.535 18.105 ;
      RECT 72.365 19.125 72.535 19.295 ;
      RECT 72.365 20.655 72.535 20.825 ;
      RECT 72.365 23.375 72.535 23.545 ;
      RECT 72.365 26.095 72.535 26.265 ;
      RECT 72.365 28.815 72.535 28.985 ;
      RECT 72.365 31.535 72.535 31.705 ;
      RECT 72.365 34.255 72.535 34.425 ;
      RECT 72.365 36.975 72.535 37.145 ;
      RECT 72.365 39.695 72.535 39.865 ;
      RECT 72.365 42.415 72.535 42.585 ;
      RECT 72.365 45.135 72.535 45.305 ;
      RECT 72.365 47.855 72.535 48.025 ;
      RECT 72.365 50.575 72.535 50.745 ;
      RECT 72.365 53.295 72.535 53.465 ;
      RECT 72.365 56.015 72.535 56.185 ;
      RECT 72.365 58.735 72.535 58.905 ;
      RECT 71.905 9.775 72.075 9.945 ;
      RECT 71.905 12.495 72.075 12.665 ;
      RECT 71.905 15.215 72.075 15.385 ;
      RECT 71.905 17.935 72.075 18.105 ;
      RECT 71.905 20.655 72.075 20.825 ;
      RECT 71.905 23.375 72.075 23.545 ;
      RECT 71.905 26.095 72.075 26.265 ;
      RECT 71.905 28.815 72.075 28.985 ;
      RECT 71.905 31.535 72.075 31.705 ;
      RECT 71.905 34.255 72.075 34.425 ;
      RECT 71.905 36.975 72.075 37.145 ;
      RECT 71.905 39.695 72.075 39.865 ;
      RECT 71.905 42.415 72.075 42.585 ;
      RECT 71.905 45.135 72.075 45.305 ;
      RECT 71.905 47.855 72.075 48.025 ;
      RECT 71.905 50.575 72.075 50.745 ;
      RECT 71.905 53.295 72.075 53.465 ;
      RECT 71.905 56.015 72.075 56.185 ;
      RECT 71.905 58.735 72.075 58.905 ;
      RECT 71.445 9.775 71.615 9.945 ;
      RECT 71.445 12.495 71.615 12.665 ;
      RECT 71.445 15.215 71.615 15.385 ;
      RECT 71.445 17.935 71.615 18.105 ;
      RECT 71.445 20.655 71.615 20.825 ;
      RECT 71.445 23.375 71.615 23.545 ;
      RECT 71.445 26.095 71.615 26.265 ;
      RECT 71.445 28.815 71.615 28.985 ;
      RECT 71.445 31.535 71.615 31.705 ;
      RECT 71.445 34.255 71.615 34.425 ;
      RECT 71.445 36.975 71.615 37.145 ;
      RECT 71.445 39.695 71.615 39.865 ;
      RECT 71.445 42.415 71.615 42.585 ;
      RECT 71.445 45.135 71.615 45.305 ;
      RECT 71.445 47.855 71.615 48.025 ;
      RECT 71.445 50.575 71.615 50.745 ;
      RECT 71.445 53.295 71.615 53.465 ;
      RECT 71.445 56.015 71.615 56.185 ;
      RECT 71.445 58.735 71.615 58.905 ;
      RECT 70.985 9.775 71.155 9.945 ;
      RECT 70.985 12.495 71.155 12.665 ;
      RECT 70.985 15.215 71.155 15.385 ;
      RECT 70.985 17.935 71.155 18.105 ;
      RECT 70.985 20.655 71.155 20.825 ;
      RECT 70.985 23.375 71.155 23.545 ;
      RECT 70.985 26.095 71.155 26.265 ;
      RECT 70.985 26.605 71.155 26.775 ;
      RECT 70.985 28.815 71.155 28.985 ;
      RECT 70.985 31.535 71.155 31.705 ;
      RECT 70.985 34.255 71.155 34.425 ;
      RECT 70.985 36.975 71.155 37.145 ;
      RECT 70.985 39.695 71.155 39.865 ;
      RECT 70.985 42.415 71.155 42.585 ;
      RECT 70.985 45.135 71.155 45.305 ;
      RECT 70.985 47.855 71.155 48.025 ;
      RECT 70.985 50.575 71.155 50.745 ;
      RECT 70.985 53.295 71.155 53.465 ;
      RECT 70.985 56.015 71.155 56.185 ;
      RECT 70.985 58.735 71.155 58.905 ;
      RECT 70.975 16.405 71.145 16.575 ;
      RECT 70.54 16.065 70.71 16.235 ;
      RECT 70.525 9.775 70.695 9.945 ;
      RECT 70.525 12.495 70.695 12.665 ;
      RECT 70.525 15.215 70.695 15.385 ;
      RECT 70.525 17.935 70.695 18.105 ;
      RECT 70.525 20.655 70.695 20.825 ;
      RECT 70.525 23.375 70.695 23.545 ;
      RECT 70.525 24.565 70.695 24.735 ;
      RECT 70.525 26.095 70.695 26.265 ;
      RECT 70.525 28.815 70.695 28.985 ;
      RECT 70.525 31.535 70.695 31.705 ;
      RECT 70.525 34.255 70.695 34.425 ;
      RECT 70.525 36.975 70.695 37.145 ;
      RECT 70.525 39.695 70.695 39.865 ;
      RECT 70.525 42.415 70.695 42.585 ;
      RECT 70.525 45.135 70.695 45.305 ;
      RECT 70.525 47.855 70.695 48.025 ;
      RECT 70.525 50.575 70.695 50.745 ;
      RECT 70.525 53.295 70.695 53.465 ;
      RECT 70.525 56.015 70.695 56.185 ;
      RECT 70.525 58.735 70.695 58.905 ;
      RECT 70.065 9.775 70.235 9.945 ;
      RECT 70.065 12.495 70.235 12.665 ;
      RECT 70.065 15.215 70.235 15.385 ;
      RECT 70.065 17.935 70.235 18.105 ;
      RECT 70.065 20.655 70.235 20.825 ;
      RECT 70.065 23.375 70.235 23.545 ;
      RECT 70.065 26.095 70.235 26.265 ;
      RECT 70.065 28.815 70.235 28.985 ;
      RECT 70.065 31.535 70.235 31.705 ;
      RECT 70.065 34.255 70.235 34.425 ;
      RECT 70.065 36.975 70.235 37.145 ;
      RECT 70.065 39.695 70.235 39.865 ;
      RECT 70.065 42.415 70.235 42.585 ;
      RECT 70.065 45.135 70.235 45.305 ;
      RECT 70.065 47.855 70.235 48.025 ;
      RECT 70.065 50.575 70.235 50.745 ;
      RECT 70.065 53.295 70.235 53.465 ;
      RECT 70.065 56.015 70.235 56.185 ;
      RECT 70.065 58.735 70.235 58.905 ;
      RECT 69.92 24.565 70.09 24.735 ;
      RECT 69.605 9.775 69.775 9.945 ;
      RECT 69.605 12.495 69.775 12.665 ;
      RECT 69.605 15.215 69.775 15.385 ;
      RECT 69.605 17.935 69.775 18.105 ;
      RECT 69.605 20.655 69.775 20.825 ;
      RECT 69.605 23.375 69.775 23.545 ;
      RECT 69.605 26.095 69.775 26.265 ;
      RECT 69.605 28.815 69.775 28.985 ;
      RECT 69.605 31.535 69.775 31.705 ;
      RECT 69.605 34.255 69.775 34.425 ;
      RECT 69.605 36.975 69.775 37.145 ;
      RECT 69.605 39.695 69.775 39.865 ;
      RECT 69.605 42.415 69.775 42.585 ;
      RECT 69.605 45.135 69.775 45.305 ;
      RECT 69.605 47.855 69.775 48.025 ;
      RECT 69.605 50.575 69.775 50.745 ;
      RECT 69.605 53.295 69.775 53.465 ;
      RECT 69.605 56.015 69.775 56.185 ;
      RECT 69.605 58.735 69.775 58.905 ;
      RECT 69.145 9.775 69.315 9.945 ;
      RECT 69.145 11.305 69.315 11.475 ;
      RECT 69.145 12.495 69.315 12.665 ;
      RECT 69.145 15.215 69.315 15.385 ;
      RECT 69.145 17.935 69.315 18.105 ;
      RECT 69.145 20.655 69.315 20.825 ;
      RECT 69.145 23.375 69.315 23.545 ;
      RECT 69.145 24.565 69.315 24.735 ;
      RECT 69.145 26.095 69.315 26.265 ;
      RECT 69.145 28.815 69.315 28.985 ;
      RECT 69.145 31.535 69.315 31.705 ;
      RECT 69.145 34.255 69.315 34.425 ;
      RECT 69.145 36.975 69.315 37.145 ;
      RECT 69.145 39.695 69.315 39.865 ;
      RECT 69.145 42.415 69.315 42.585 ;
      RECT 69.145 45.135 69.315 45.305 ;
      RECT 69.145 47.855 69.315 48.025 ;
      RECT 69.145 50.575 69.315 50.745 ;
      RECT 69.145 53.295 69.315 53.465 ;
      RECT 69.145 56.015 69.315 56.185 ;
      RECT 69.145 58.735 69.315 58.905 ;
      RECT 68.97 16.065 69.14 16.235 ;
      RECT 68.685 9.775 68.855 9.945 ;
      RECT 68.685 12.495 68.855 12.665 ;
      RECT 68.685 15.215 68.855 15.385 ;
      RECT 68.685 17.935 68.855 18.105 ;
      RECT 68.685 20.655 68.855 20.825 ;
      RECT 68.685 23.375 68.855 23.545 ;
      RECT 68.685 24.225 68.855 24.395 ;
      RECT 68.685 26.095 68.855 26.265 ;
      RECT 68.685 28.815 68.855 28.985 ;
      RECT 68.685 31.535 68.855 31.705 ;
      RECT 68.685 34.255 68.855 34.425 ;
      RECT 68.685 36.975 68.855 37.145 ;
      RECT 68.685 39.695 68.855 39.865 ;
      RECT 68.685 42.415 68.855 42.585 ;
      RECT 68.685 45.135 68.855 45.305 ;
      RECT 68.685 47.855 68.855 48.025 ;
      RECT 68.685 50.575 68.855 50.745 ;
      RECT 68.685 53.295 68.855 53.465 ;
      RECT 68.685 56.015 68.855 56.185 ;
      RECT 68.685 58.735 68.855 58.905 ;
      RECT 68.675 27.285 68.845 27.455 ;
      RECT 68.455 16.405 68.625 16.575 ;
      RECT 68.24 26.945 68.41 27.115 ;
      RECT 68.225 9.775 68.395 9.945 ;
      RECT 68.225 12.495 68.395 12.665 ;
      RECT 68.225 15.215 68.395 15.385 ;
      RECT 68.225 17.935 68.395 18.105 ;
      RECT 68.225 20.655 68.395 20.825 ;
      RECT 68.225 22.865 68.395 23.035 ;
      RECT 68.225 23.375 68.395 23.545 ;
      RECT 68.225 26.095 68.395 26.265 ;
      RECT 68.225 28.815 68.395 28.985 ;
      RECT 68.225 31.535 68.395 31.705 ;
      RECT 68.225 34.255 68.395 34.425 ;
      RECT 68.225 36.975 68.395 37.145 ;
      RECT 68.225 39.695 68.395 39.865 ;
      RECT 68.225 42.415 68.395 42.585 ;
      RECT 68.225 45.135 68.395 45.305 ;
      RECT 68.225 47.855 68.395 48.025 ;
      RECT 68.225 50.575 68.395 50.745 ;
      RECT 68.225 53.295 68.395 53.465 ;
      RECT 68.225 56.015 68.395 56.185 ;
      RECT 68.225 58.735 68.395 58.905 ;
      RECT 67.995 24.565 68.165 24.735 ;
      RECT 67.765 9.775 67.935 9.945 ;
      RECT 67.765 12.495 67.935 12.665 ;
      RECT 67.765 15.215 67.935 15.385 ;
      RECT 67.765 17.935 67.935 18.105 ;
      RECT 67.765 20.145 67.935 20.315 ;
      RECT 67.765 20.655 67.935 20.825 ;
      RECT 67.765 23.375 67.935 23.545 ;
      RECT 67.765 26.095 67.935 26.265 ;
      RECT 67.765 28.815 67.935 28.985 ;
      RECT 67.765 31.535 67.935 31.705 ;
      RECT 67.765 34.255 67.935 34.425 ;
      RECT 67.765 36.975 67.935 37.145 ;
      RECT 67.765 39.695 67.935 39.865 ;
      RECT 67.765 42.415 67.935 42.585 ;
      RECT 67.765 45.135 67.935 45.305 ;
      RECT 67.765 47.855 67.935 48.025 ;
      RECT 67.765 50.575 67.935 50.745 ;
      RECT 67.765 53.295 67.935 53.465 ;
      RECT 67.765 56.015 67.935 56.185 ;
      RECT 67.765 58.735 67.935 58.905 ;
      RECT 67.69 17.085 67.86 17.255 ;
      RECT 67.535 22.185 67.705 22.355 ;
      RECT 67.305 9.775 67.475 9.945 ;
      RECT 67.305 12.495 67.475 12.665 ;
      RECT 67.305 15.215 67.475 15.385 ;
      RECT 67.305 17.935 67.475 18.105 ;
      RECT 67.305 20.655 67.475 20.825 ;
      RECT 67.305 23.375 67.475 23.545 ;
      RECT 67.305 25.585 67.475 25.755 ;
      RECT 67.305 26.095 67.475 26.265 ;
      RECT 67.305 28.815 67.475 28.985 ;
      RECT 67.305 31.535 67.475 31.705 ;
      RECT 67.305 34.255 67.475 34.425 ;
      RECT 67.305 36.975 67.475 37.145 ;
      RECT 67.305 39.695 67.475 39.865 ;
      RECT 67.305 42.415 67.475 42.585 ;
      RECT 67.305 45.135 67.475 45.305 ;
      RECT 67.305 47.855 67.475 48.025 ;
      RECT 67.305 50.575 67.475 50.745 ;
      RECT 67.305 53.295 67.475 53.465 ;
      RECT 67.305 56.015 67.475 56.185 ;
      RECT 67.305 58.735 67.475 58.905 ;
      RECT 67.265 16.405 67.435 16.575 ;
      RECT 66.87 16.065 67.04 16.235 ;
      RECT 66.87 19.125 67.04 19.295 ;
      RECT 66.845 9.775 67.015 9.945 ;
      RECT 66.845 12.495 67.015 12.665 ;
      RECT 66.845 14.705 67.015 14.875 ;
      RECT 66.845 15.215 67.015 15.385 ;
      RECT 66.845 17.935 67.015 18.105 ;
      RECT 66.845 20.655 67.015 20.825 ;
      RECT 66.845 22.525 67.015 22.695 ;
      RECT 66.845 23.375 67.015 23.545 ;
      RECT 66.845 26.095 67.015 26.265 ;
      RECT 66.845 28.815 67.015 28.985 ;
      RECT 66.845 31.535 67.015 31.705 ;
      RECT 66.845 34.255 67.015 34.425 ;
      RECT 66.845 36.975 67.015 37.145 ;
      RECT 66.845 38.505 67.015 38.675 ;
      RECT 66.845 39.695 67.015 39.865 ;
      RECT 66.845 42.415 67.015 42.585 ;
      RECT 66.845 45.135 67.015 45.305 ;
      RECT 66.845 47.855 67.015 48.025 ;
      RECT 66.845 50.575 67.015 50.745 ;
      RECT 66.845 53.295 67.015 53.465 ;
      RECT 66.845 56.015 67.015 56.185 ;
      RECT 66.845 58.735 67.015 58.905 ;
      RECT 66.67 26.945 66.84 27.115 ;
      RECT 66.385 9.775 66.555 9.945 ;
      RECT 66.385 12.495 66.555 12.665 ;
      RECT 66.385 15.215 66.555 15.385 ;
      RECT 66.385 16.745 66.555 16.915 ;
      RECT 66.385 17.935 66.555 18.105 ;
      RECT 66.385 19.125 66.555 19.295 ;
      RECT 66.385 20.655 66.555 20.825 ;
      RECT 66.385 22.525 66.555 22.695 ;
      RECT 66.385 23.375 66.555 23.545 ;
      RECT 66.385 26.095 66.555 26.265 ;
      RECT 66.385 28.815 66.555 28.985 ;
      RECT 66.385 31.535 66.555 31.705 ;
      RECT 66.385 34.255 66.555 34.425 ;
      RECT 66.385 36.975 66.555 37.145 ;
      RECT 66.385 39.695 66.555 39.865 ;
      RECT 66.385 42.415 66.555 42.585 ;
      RECT 66.385 45.135 66.555 45.305 ;
      RECT 66.385 47.855 66.555 48.025 ;
      RECT 66.385 50.575 66.555 50.745 ;
      RECT 66.385 53.295 66.555 53.465 ;
      RECT 66.385 56.015 66.555 56.185 ;
      RECT 66.385 58.735 66.555 58.905 ;
      RECT 66.155 13.685 66.325 13.855 ;
      RECT 66.155 27.285 66.325 27.455 ;
      RECT 65.925 9.775 66.095 9.945 ;
      RECT 65.925 12.495 66.095 12.665 ;
      RECT 65.925 15.215 66.095 15.385 ;
      RECT 65.925 17.935 66.095 18.105 ;
      RECT 65.925 19.125 66.095 19.295 ;
      RECT 65.925 20.655 66.095 20.825 ;
      RECT 65.925 23.375 66.095 23.545 ;
      RECT 65.925 26.095 66.095 26.265 ;
      RECT 65.925 28.815 66.095 28.985 ;
      RECT 65.925 31.535 66.095 31.705 ;
      RECT 65.925 34.255 66.095 34.425 ;
      RECT 65.925 36.975 66.095 37.145 ;
      RECT 65.925 39.695 66.095 39.865 ;
      RECT 65.925 42.415 66.095 42.585 ;
      RECT 65.925 45.135 66.095 45.305 ;
      RECT 65.925 47.855 66.095 48.025 ;
      RECT 65.925 50.575 66.095 50.745 ;
      RECT 65.925 53.295 66.095 53.465 ;
      RECT 65.925 56.015 66.095 56.185 ;
      RECT 65.925 58.735 66.095 58.905 ;
      RECT 65.695 22.185 65.865 22.355 ;
      RECT 65.465 9.775 65.635 9.945 ;
      RECT 65.465 12.495 65.635 12.665 ;
      RECT 65.465 13.685 65.635 13.855 ;
      RECT 65.465 15.215 65.635 15.385 ;
      RECT 65.465 17.935 65.635 18.105 ;
      RECT 65.465 20.655 65.635 20.825 ;
      RECT 65.465 23.375 65.635 23.545 ;
      RECT 65.465 26.095 65.635 26.265 ;
      RECT 65.465 28.815 65.635 28.985 ;
      RECT 65.465 31.535 65.635 31.705 ;
      RECT 65.465 34.255 65.635 34.425 ;
      RECT 65.465 36.975 65.635 37.145 ;
      RECT 65.465 39.695 65.635 39.865 ;
      RECT 65.465 42.415 65.635 42.585 ;
      RECT 65.465 45.135 65.635 45.305 ;
      RECT 65.465 47.855 65.635 48.025 ;
      RECT 65.465 50.575 65.635 50.745 ;
      RECT 65.465 53.295 65.635 53.465 ;
      RECT 65.465 56.015 65.635 56.185 ;
      RECT 65.465 58.735 65.635 58.905 ;
      RECT 65.39 27.965 65.56 28.135 ;
      RECT 65.01 19.135 65.18 19.305 ;
      RECT 65.005 9.775 65.175 9.945 ;
      RECT 65.005 12.495 65.175 12.665 ;
      RECT 65.005 13.345 65.175 13.515 ;
      RECT 65.005 15.215 65.175 15.385 ;
      RECT 65.005 16.745 65.175 16.915 ;
      RECT 65.005 17.935 65.175 18.105 ;
      RECT 65.005 20.655 65.175 20.825 ;
      RECT 65.005 22.185 65.175 22.355 ;
      RECT 65.005 23.375 65.175 23.545 ;
      RECT 65.005 26.095 65.175 26.265 ;
      RECT 65.005 28.815 65.175 28.985 ;
      RECT 65.005 31.535 65.175 31.705 ;
      RECT 65.005 34.255 65.175 34.425 ;
      RECT 65.005 36.975 65.175 37.145 ;
      RECT 65.005 39.695 65.175 39.865 ;
      RECT 65.005 42.415 65.175 42.585 ;
      RECT 65.005 45.135 65.175 45.305 ;
      RECT 65.005 47.855 65.175 48.025 ;
      RECT 65.005 50.575 65.175 50.745 ;
      RECT 65.005 53.295 65.175 53.465 ;
      RECT 65.005 56.015 65.175 56.185 ;
      RECT 65.005 58.735 65.175 58.905 ;
      RECT 64.965 27.285 65.135 27.455 ;
      RECT 64.57 26.945 64.74 27.115 ;
      RECT 64.545 9.775 64.715 9.945 ;
      RECT 64.545 12.495 64.715 12.665 ;
      RECT 64.545 15.215 64.715 15.385 ;
      RECT 64.545 17.935 64.715 18.105 ;
      RECT 64.545 19.125 64.715 19.295 ;
      RECT 64.545 20.655 64.715 20.825 ;
      RECT 64.545 23.375 64.715 23.545 ;
      RECT 64.545 26.095 64.715 26.265 ;
      RECT 64.545 28.815 64.715 28.985 ;
      RECT 64.545 31.535 64.715 31.705 ;
      RECT 64.545 34.255 64.715 34.425 ;
      RECT 64.545 36.975 64.715 37.145 ;
      RECT 64.545 39.695 64.715 39.865 ;
      RECT 64.545 42.415 64.715 42.585 ;
      RECT 64.545 45.135 64.715 45.305 ;
      RECT 64.545 47.855 64.715 48.025 ;
      RECT 64.545 50.575 64.715 50.745 ;
      RECT 64.545 53.295 64.715 53.465 ;
      RECT 64.545 56.015 64.715 56.185 ;
      RECT 64.545 58.735 64.715 58.905 ;
      RECT 64.315 13.685 64.485 13.855 ;
      RECT 64.085 9.775 64.255 9.945 ;
      RECT 64.085 12.495 64.255 12.665 ;
      RECT 64.085 15.215 64.255 15.385 ;
      RECT 64.085 17.935 64.255 18.105 ;
      RECT 64.085 20.655 64.255 20.825 ;
      RECT 64.085 23.375 64.255 23.545 ;
      RECT 64.085 26.095 64.255 26.265 ;
      RECT 64.085 27.625 64.255 27.795 ;
      RECT 64.085 28.815 64.255 28.985 ;
      RECT 64.085 31.535 64.255 31.705 ;
      RECT 64.085 34.255 64.255 34.425 ;
      RECT 64.085 36.975 64.255 37.145 ;
      RECT 64.085 39.695 64.255 39.865 ;
      RECT 64.085 42.415 64.255 42.585 ;
      RECT 64.085 45.135 64.255 45.305 ;
      RECT 64.085 47.855 64.255 48.025 ;
      RECT 64.085 50.575 64.255 50.745 ;
      RECT 64.085 53.295 64.255 53.465 ;
      RECT 64.085 56.015 64.255 56.185 ;
      RECT 64.085 58.735 64.255 58.905 ;
      RECT 63.625 9.775 63.795 9.945 ;
      RECT 63.625 12.495 63.795 12.665 ;
      RECT 63.625 13.685 63.795 13.855 ;
      RECT 63.625 15.215 63.795 15.385 ;
      RECT 63.625 17.935 63.795 18.105 ;
      RECT 63.625 20.655 63.795 20.825 ;
      RECT 63.625 23.375 63.795 23.545 ;
      RECT 63.625 26.095 63.795 26.265 ;
      RECT 63.625 28.815 63.795 28.985 ;
      RECT 63.625 31.535 63.795 31.705 ;
      RECT 63.625 34.255 63.795 34.425 ;
      RECT 63.625 36.975 63.795 37.145 ;
      RECT 63.625 39.695 63.795 39.865 ;
      RECT 63.625 42.415 63.795 42.585 ;
      RECT 63.625 45.135 63.795 45.305 ;
      RECT 63.625 47.855 63.795 48.025 ;
      RECT 63.625 50.575 63.795 50.745 ;
      RECT 63.625 53.295 63.795 53.465 ;
      RECT 63.625 56.015 63.795 56.185 ;
      RECT 63.625 58.735 63.795 58.905 ;
      RECT 63.165 9.775 63.335 9.945 ;
      RECT 63.165 12.495 63.335 12.665 ;
      RECT 63.165 15.215 63.335 15.385 ;
      RECT 63.165 17.935 63.335 18.105 ;
      RECT 63.165 20.655 63.335 20.825 ;
      RECT 63.165 23.375 63.335 23.545 ;
      RECT 63.165 26.095 63.335 26.265 ;
      RECT 63.165 28.815 63.335 28.985 ;
      RECT 63.165 31.535 63.335 31.705 ;
      RECT 63.165 34.255 63.335 34.425 ;
      RECT 63.165 36.975 63.335 37.145 ;
      RECT 63.165 39.695 63.335 39.865 ;
      RECT 63.165 42.415 63.335 42.585 ;
      RECT 63.165 45.135 63.335 45.305 ;
      RECT 63.165 47.855 63.335 48.025 ;
      RECT 63.165 50.575 63.335 50.745 ;
      RECT 63.165 53.295 63.335 53.465 ;
      RECT 63.165 56.015 63.335 56.185 ;
      RECT 63.165 58.735 63.335 58.905 ;
      RECT 62.705 9.775 62.875 9.945 ;
      RECT 62.705 12.495 62.875 12.665 ;
      RECT 62.705 15.215 62.875 15.385 ;
      RECT 62.705 17.935 62.875 18.105 ;
      RECT 62.705 20.655 62.875 20.825 ;
      RECT 62.705 23.375 62.875 23.545 ;
      RECT 62.705 26.095 62.875 26.265 ;
      RECT 62.705 28.815 62.875 28.985 ;
      RECT 62.705 31.535 62.875 31.705 ;
      RECT 62.705 34.255 62.875 34.425 ;
      RECT 62.705 36.975 62.875 37.145 ;
      RECT 62.705 39.695 62.875 39.865 ;
      RECT 62.705 42.415 62.875 42.585 ;
      RECT 62.705 45.135 62.875 45.305 ;
      RECT 62.705 47.855 62.875 48.025 ;
      RECT 62.705 50.575 62.875 50.745 ;
      RECT 62.705 53.295 62.875 53.465 ;
      RECT 62.705 56.015 62.875 56.185 ;
      RECT 62.705 58.735 62.875 58.905 ;
      RECT 62.245 9.775 62.415 9.945 ;
      RECT 62.245 12.495 62.415 12.665 ;
      RECT 62.245 15.215 62.415 15.385 ;
      RECT 62.245 17.935 62.415 18.105 ;
      RECT 62.245 20.655 62.415 20.825 ;
      RECT 62.245 23.375 62.415 23.545 ;
      RECT 62.245 26.095 62.415 26.265 ;
      RECT 62.245 28.815 62.415 28.985 ;
      RECT 62.245 31.535 62.415 31.705 ;
      RECT 62.245 34.255 62.415 34.425 ;
      RECT 62.245 36.975 62.415 37.145 ;
      RECT 62.245 39.695 62.415 39.865 ;
      RECT 62.245 42.415 62.415 42.585 ;
      RECT 62.245 45.135 62.415 45.305 ;
      RECT 62.245 47.855 62.415 48.025 ;
      RECT 62.245 50.575 62.415 50.745 ;
      RECT 62.245 53.295 62.415 53.465 ;
      RECT 62.245 56.015 62.415 56.185 ;
      RECT 62.245 58.735 62.415 58.905 ;
      RECT 61.785 9.775 61.955 9.945 ;
      RECT 61.785 12.495 61.955 12.665 ;
      RECT 61.785 15.215 61.955 15.385 ;
      RECT 61.785 17.935 61.955 18.105 ;
      RECT 61.785 20.655 61.955 20.825 ;
      RECT 61.785 23.375 61.955 23.545 ;
      RECT 61.785 26.095 61.955 26.265 ;
      RECT 61.785 28.815 61.955 28.985 ;
      RECT 61.785 31.535 61.955 31.705 ;
      RECT 61.785 34.255 61.955 34.425 ;
      RECT 61.785 36.975 61.955 37.145 ;
      RECT 61.785 39.695 61.955 39.865 ;
      RECT 61.785 42.415 61.955 42.585 ;
      RECT 61.785 45.135 61.955 45.305 ;
      RECT 61.785 47.855 61.955 48.025 ;
      RECT 61.785 50.575 61.955 50.745 ;
      RECT 61.785 53.295 61.955 53.465 ;
      RECT 61.785 56.015 61.955 56.185 ;
      RECT 61.785 58.735 61.955 58.905 ;
      RECT 61.325 9.775 61.495 9.945 ;
      RECT 61.325 12.495 61.495 12.665 ;
      RECT 61.325 15.215 61.495 15.385 ;
      RECT 61.325 17.935 61.495 18.105 ;
      RECT 61.325 19.125 61.495 19.295 ;
      RECT 61.325 20.655 61.495 20.825 ;
      RECT 61.325 23.375 61.495 23.545 ;
      RECT 61.325 26.095 61.495 26.265 ;
      RECT 61.325 28.815 61.495 28.985 ;
      RECT 61.325 31.535 61.495 31.705 ;
      RECT 61.325 34.255 61.495 34.425 ;
      RECT 61.325 36.975 61.495 37.145 ;
      RECT 61.325 39.695 61.495 39.865 ;
      RECT 61.325 42.415 61.495 42.585 ;
      RECT 61.325 45.135 61.495 45.305 ;
      RECT 61.325 47.855 61.495 48.025 ;
      RECT 61.325 50.575 61.495 50.745 ;
      RECT 61.325 53.295 61.495 53.465 ;
      RECT 61.325 56.015 61.495 56.185 ;
      RECT 61.325 58.735 61.495 58.905 ;
      RECT 60.865 9.775 61.035 9.945 ;
      RECT 60.865 12.495 61.035 12.665 ;
      RECT 60.865 15.215 61.035 15.385 ;
      RECT 60.865 17.935 61.035 18.105 ;
      RECT 60.865 20.655 61.035 20.825 ;
      RECT 60.865 23.375 61.035 23.545 ;
      RECT 60.865 26.095 61.035 26.265 ;
      RECT 60.865 28.815 61.035 28.985 ;
      RECT 60.865 31.535 61.035 31.705 ;
      RECT 60.865 34.255 61.035 34.425 ;
      RECT 60.865 36.975 61.035 37.145 ;
      RECT 60.865 39.695 61.035 39.865 ;
      RECT 60.865 42.415 61.035 42.585 ;
      RECT 60.865 45.135 61.035 45.305 ;
      RECT 60.865 47.855 61.035 48.025 ;
      RECT 60.865 50.575 61.035 50.745 ;
      RECT 60.865 53.295 61.035 53.465 ;
      RECT 60.865 56.015 61.035 56.185 ;
      RECT 60.865 58.735 61.035 58.905 ;
      RECT 60.405 9.775 60.575 9.945 ;
      RECT 60.405 12.495 60.575 12.665 ;
      RECT 60.405 15.215 60.575 15.385 ;
      RECT 60.405 17.935 60.575 18.105 ;
      RECT 60.405 20.655 60.575 20.825 ;
      RECT 60.405 23.375 60.575 23.545 ;
      RECT 60.405 26.095 60.575 26.265 ;
      RECT 60.405 28.815 60.575 28.985 ;
      RECT 60.405 31.535 60.575 31.705 ;
      RECT 60.405 34.255 60.575 34.425 ;
      RECT 60.405 36.975 60.575 37.145 ;
      RECT 60.405 39.695 60.575 39.865 ;
      RECT 60.405 42.415 60.575 42.585 ;
      RECT 60.405 45.135 60.575 45.305 ;
      RECT 60.405 47.855 60.575 48.025 ;
      RECT 60.405 50.575 60.575 50.745 ;
      RECT 60.405 53.295 60.575 53.465 ;
      RECT 60.405 56.015 60.575 56.185 ;
      RECT 60.405 58.735 60.575 58.905 ;
      RECT 59.945 9.775 60.115 9.945 ;
      RECT 59.945 11.985 60.115 12.155 ;
      RECT 59.945 12.495 60.115 12.665 ;
      RECT 59.945 15.215 60.115 15.385 ;
      RECT 59.945 17.935 60.115 18.105 ;
      RECT 59.945 20.655 60.115 20.825 ;
      RECT 59.945 23.375 60.115 23.545 ;
      RECT 59.945 26.095 60.115 26.265 ;
      RECT 59.945 28.815 60.115 28.985 ;
      RECT 59.945 31.535 60.115 31.705 ;
      RECT 59.945 34.255 60.115 34.425 ;
      RECT 59.945 36.975 60.115 37.145 ;
      RECT 59.945 39.695 60.115 39.865 ;
      RECT 59.945 42.415 60.115 42.585 ;
      RECT 59.945 45.135 60.115 45.305 ;
      RECT 59.945 47.855 60.115 48.025 ;
      RECT 59.945 50.575 60.115 50.745 ;
      RECT 59.945 53.295 60.115 53.465 ;
      RECT 59.945 56.015 60.115 56.185 ;
      RECT 59.945 58.735 60.115 58.905 ;
      RECT 59.485 9.775 59.655 9.945 ;
      RECT 59.485 12.495 59.655 12.665 ;
      RECT 59.485 15.215 59.655 15.385 ;
      RECT 59.485 17.935 59.655 18.105 ;
      RECT 59.485 19.125 59.655 19.295 ;
      RECT 59.485 20.655 59.655 20.825 ;
      RECT 59.485 23.375 59.655 23.545 ;
      RECT 59.485 26.095 59.655 26.265 ;
      RECT 59.485 28.815 59.655 28.985 ;
      RECT 59.485 31.535 59.655 31.705 ;
      RECT 59.485 34.255 59.655 34.425 ;
      RECT 59.485 36.975 59.655 37.145 ;
      RECT 59.485 39.695 59.655 39.865 ;
      RECT 59.485 42.415 59.655 42.585 ;
      RECT 59.485 45.135 59.655 45.305 ;
      RECT 59.485 47.855 59.655 48.025 ;
      RECT 59.485 50.575 59.655 50.745 ;
      RECT 59.485 53.295 59.655 53.465 ;
      RECT 59.485 56.015 59.655 56.185 ;
      RECT 59.485 58.735 59.655 58.905 ;
      RECT 59.025 9.775 59.195 9.945 ;
      RECT 59.025 12.495 59.195 12.665 ;
      RECT 59.025 15.215 59.195 15.385 ;
      RECT 59.025 17.935 59.195 18.105 ;
      RECT 59.025 20.655 59.195 20.825 ;
      RECT 59.025 23.375 59.195 23.545 ;
      RECT 59.025 26.095 59.195 26.265 ;
      RECT 59.025 28.815 59.195 28.985 ;
      RECT 59.025 31.535 59.195 31.705 ;
      RECT 59.025 34.255 59.195 34.425 ;
      RECT 59.025 36.975 59.195 37.145 ;
      RECT 59.025 39.695 59.195 39.865 ;
      RECT 59.025 42.415 59.195 42.585 ;
      RECT 59.025 45.135 59.195 45.305 ;
      RECT 59.025 47.855 59.195 48.025 ;
      RECT 59.025 50.575 59.195 50.745 ;
      RECT 59.025 53.295 59.195 53.465 ;
      RECT 59.025 56.015 59.195 56.185 ;
      RECT 59.025 58.735 59.195 58.905 ;
      RECT 58.565 9.775 58.735 9.945 ;
      RECT 58.565 12.495 58.735 12.665 ;
      RECT 58.565 15.215 58.735 15.385 ;
      RECT 58.565 15.725 58.735 15.895 ;
      RECT 58.565 17.425 58.735 17.595 ;
      RECT 58.565 17.935 58.735 18.105 ;
      RECT 58.565 20.655 58.735 20.825 ;
      RECT 58.565 23.375 58.735 23.545 ;
      RECT 58.565 26.095 58.735 26.265 ;
      RECT 58.565 26.605 58.735 26.775 ;
      RECT 58.565 28.815 58.735 28.985 ;
      RECT 58.565 31.535 58.735 31.705 ;
      RECT 58.565 34.255 58.735 34.425 ;
      RECT 58.565 36.975 58.735 37.145 ;
      RECT 58.565 39.695 58.735 39.865 ;
      RECT 58.565 42.415 58.735 42.585 ;
      RECT 58.565 45.135 58.735 45.305 ;
      RECT 58.565 47.855 58.735 48.025 ;
      RECT 58.565 50.575 58.735 50.745 ;
      RECT 58.565 53.295 58.735 53.465 ;
      RECT 58.565 56.015 58.735 56.185 ;
      RECT 58.565 58.735 58.735 58.905 ;
      RECT 58.105 9.775 58.275 9.945 ;
      RECT 58.105 12.495 58.275 12.665 ;
      RECT 58.105 15.215 58.275 15.385 ;
      RECT 58.105 17.935 58.275 18.105 ;
      RECT 58.105 20.655 58.275 20.825 ;
      RECT 58.105 23.375 58.275 23.545 ;
      RECT 58.105 26.095 58.275 26.265 ;
      RECT 58.105 28.815 58.275 28.985 ;
      RECT 58.105 31.535 58.275 31.705 ;
      RECT 58.105 34.255 58.275 34.425 ;
      RECT 58.105 36.975 58.275 37.145 ;
      RECT 58.105 39.695 58.275 39.865 ;
      RECT 58.105 42.415 58.275 42.585 ;
      RECT 58.105 45.135 58.275 45.305 ;
      RECT 58.105 47.855 58.275 48.025 ;
      RECT 58.105 50.575 58.275 50.745 ;
      RECT 58.105 53.295 58.275 53.465 ;
      RECT 58.105 56.015 58.275 56.185 ;
      RECT 58.105 58.735 58.275 58.905 ;
      RECT 57.645 9.775 57.815 9.945 ;
      RECT 57.645 12.495 57.815 12.665 ;
      RECT 57.645 15.215 57.815 15.385 ;
      RECT 57.645 17.935 57.815 18.105 ;
      RECT 57.645 20.655 57.815 20.825 ;
      RECT 57.645 23.375 57.815 23.545 ;
      RECT 57.645 26.095 57.815 26.265 ;
      RECT 57.645 28.815 57.815 28.985 ;
      RECT 57.645 31.535 57.815 31.705 ;
      RECT 57.645 34.255 57.815 34.425 ;
      RECT 57.645 36.975 57.815 37.145 ;
      RECT 57.645 39.695 57.815 39.865 ;
      RECT 57.645 42.415 57.815 42.585 ;
      RECT 57.645 45.135 57.815 45.305 ;
      RECT 57.645 47.855 57.815 48.025 ;
      RECT 57.645 50.575 57.815 50.745 ;
      RECT 57.645 53.295 57.815 53.465 ;
      RECT 57.645 56.015 57.815 56.185 ;
      RECT 57.645 58.735 57.815 58.905 ;
      RECT 57.185 9.775 57.355 9.945 ;
      RECT 57.185 12.495 57.355 12.665 ;
      RECT 57.185 15.215 57.355 15.385 ;
      RECT 57.185 17.935 57.355 18.105 ;
      RECT 57.185 20.655 57.355 20.825 ;
      RECT 57.185 23.375 57.355 23.545 ;
      RECT 57.185 26.095 57.355 26.265 ;
      RECT 57.185 28.815 57.355 28.985 ;
      RECT 57.185 31.535 57.355 31.705 ;
      RECT 57.185 34.255 57.355 34.425 ;
      RECT 57.185 36.975 57.355 37.145 ;
      RECT 57.185 39.695 57.355 39.865 ;
      RECT 57.185 42.415 57.355 42.585 ;
      RECT 57.185 45.135 57.355 45.305 ;
      RECT 57.185 47.855 57.355 48.025 ;
      RECT 57.185 50.575 57.355 50.745 ;
      RECT 57.185 53.295 57.355 53.465 ;
      RECT 57.185 56.015 57.355 56.185 ;
      RECT 57.185 58.735 57.355 58.905 ;
      RECT 56.725 9.775 56.895 9.945 ;
      RECT 56.725 12.495 56.895 12.665 ;
      RECT 56.725 15.215 56.895 15.385 ;
      RECT 56.725 17.935 56.895 18.105 ;
      RECT 56.725 20.655 56.895 20.825 ;
      RECT 56.725 23.375 56.895 23.545 ;
      RECT 56.725 26.095 56.895 26.265 ;
      RECT 56.725 28.815 56.895 28.985 ;
      RECT 56.725 31.535 56.895 31.705 ;
      RECT 56.725 34.255 56.895 34.425 ;
      RECT 56.725 36.975 56.895 37.145 ;
      RECT 56.725 39.695 56.895 39.865 ;
      RECT 56.725 42.415 56.895 42.585 ;
      RECT 56.725 45.135 56.895 45.305 ;
      RECT 56.725 47.855 56.895 48.025 ;
      RECT 56.725 50.575 56.895 50.745 ;
      RECT 56.725 53.295 56.895 53.465 ;
      RECT 56.725 56.015 56.895 56.185 ;
      RECT 56.725 58.735 56.895 58.905 ;
      RECT 56.265 9.775 56.435 9.945 ;
      RECT 56.265 12.495 56.435 12.665 ;
      RECT 56.265 15.215 56.435 15.385 ;
      RECT 56.265 17.935 56.435 18.105 ;
      RECT 56.265 20.655 56.435 20.825 ;
      RECT 56.265 23.375 56.435 23.545 ;
      RECT 56.265 26.095 56.435 26.265 ;
      RECT 56.265 28.815 56.435 28.985 ;
      RECT 56.265 31.535 56.435 31.705 ;
      RECT 56.265 34.255 56.435 34.425 ;
      RECT 56.265 36.975 56.435 37.145 ;
      RECT 56.265 39.695 56.435 39.865 ;
      RECT 56.265 42.415 56.435 42.585 ;
      RECT 56.265 45.135 56.435 45.305 ;
      RECT 56.265 47.855 56.435 48.025 ;
      RECT 56.265 50.575 56.435 50.745 ;
      RECT 56.265 53.295 56.435 53.465 ;
      RECT 56.265 56.015 56.435 56.185 ;
      RECT 56.265 58.735 56.435 58.905 ;
      RECT 56.255 16.405 56.425 16.575 ;
      RECT 56.255 27.285 56.425 27.455 ;
      RECT 55.82 16.065 55.99 16.235 ;
      RECT 55.82 26.945 55.99 27.115 ;
      RECT 55.805 9.775 55.975 9.945 ;
      RECT 55.805 12.495 55.975 12.665 ;
      RECT 55.805 13.685 55.975 13.855 ;
      RECT 55.805 15.215 55.975 15.385 ;
      RECT 55.805 17.935 55.975 18.105 ;
      RECT 55.805 20.655 55.975 20.825 ;
      RECT 55.805 23.375 55.975 23.545 ;
      RECT 55.805 26.095 55.975 26.265 ;
      RECT 55.805 28.815 55.975 28.985 ;
      RECT 55.805 31.535 55.975 31.705 ;
      RECT 55.805 34.255 55.975 34.425 ;
      RECT 55.805 36.975 55.975 37.145 ;
      RECT 55.805 39.695 55.975 39.865 ;
      RECT 55.805 42.415 55.975 42.585 ;
      RECT 55.805 45.135 55.975 45.305 ;
      RECT 55.805 47.855 55.975 48.025 ;
      RECT 55.805 50.575 55.975 50.745 ;
      RECT 55.805 53.295 55.975 53.465 ;
      RECT 55.805 56.015 55.975 56.185 ;
      RECT 55.805 58.735 55.975 58.905 ;
      RECT 55.345 9.775 55.515 9.945 ;
      RECT 55.345 12.495 55.515 12.665 ;
      RECT 55.345 15.215 55.515 15.385 ;
      RECT 55.345 17.935 55.515 18.105 ;
      RECT 55.345 20.655 55.515 20.825 ;
      RECT 55.345 23.375 55.515 23.545 ;
      RECT 55.345 26.095 55.515 26.265 ;
      RECT 55.345 28.815 55.515 28.985 ;
      RECT 55.345 31.535 55.515 31.705 ;
      RECT 55.345 34.255 55.515 34.425 ;
      RECT 55.345 36.975 55.515 37.145 ;
      RECT 55.345 39.695 55.515 39.865 ;
      RECT 55.345 42.415 55.515 42.585 ;
      RECT 55.345 45.135 55.515 45.305 ;
      RECT 55.345 47.855 55.515 48.025 ;
      RECT 55.345 50.575 55.515 50.745 ;
      RECT 55.345 53.295 55.515 53.465 ;
      RECT 55.345 56.015 55.515 56.185 ;
      RECT 55.345 58.735 55.515 58.905 ;
      RECT 55.115 13.685 55.285 13.855 ;
      RECT 54.885 9.775 55.055 9.945 ;
      RECT 54.885 12.495 55.055 12.665 ;
      RECT 54.885 15.215 55.055 15.385 ;
      RECT 54.885 17.935 55.055 18.105 ;
      RECT 54.885 20.655 55.055 20.825 ;
      RECT 54.885 23.375 55.055 23.545 ;
      RECT 54.885 26.095 55.055 26.265 ;
      RECT 54.885 28.815 55.055 28.985 ;
      RECT 54.885 31.535 55.055 31.705 ;
      RECT 54.885 34.255 55.055 34.425 ;
      RECT 54.885 36.975 55.055 37.145 ;
      RECT 54.885 39.695 55.055 39.865 ;
      RECT 54.885 42.415 55.055 42.585 ;
      RECT 54.885 45.135 55.055 45.305 ;
      RECT 54.885 47.855 55.055 48.025 ;
      RECT 54.885 50.575 55.055 50.745 ;
      RECT 54.885 53.295 55.055 53.465 ;
      RECT 54.885 56.015 55.055 56.185 ;
      RECT 54.885 58.735 55.055 58.905 ;
      RECT 54.425 9.775 54.595 9.945 ;
      RECT 54.425 12.495 54.595 12.665 ;
      RECT 54.425 13.685 54.595 13.855 ;
      RECT 54.425 15.215 54.595 15.385 ;
      RECT 54.425 17.935 54.595 18.105 ;
      RECT 54.425 20.655 54.595 20.825 ;
      RECT 54.425 23.375 54.595 23.545 ;
      RECT 54.425 26.095 54.595 26.265 ;
      RECT 54.425 28.815 54.595 28.985 ;
      RECT 54.425 31.535 54.595 31.705 ;
      RECT 54.425 34.255 54.595 34.425 ;
      RECT 54.425 36.975 54.595 37.145 ;
      RECT 54.425 39.695 54.595 39.865 ;
      RECT 54.425 42.415 54.595 42.585 ;
      RECT 54.425 45.135 54.595 45.305 ;
      RECT 54.425 47.855 54.595 48.025 ;
      RECT 54.425 50.575 54.595 50.745 ;
      RECT 54.425 53.295 54.595 53.465 ;
      RECT 54.425 56.015 54.595 56.185 ;
      RECT 54.425 58.735 54.595 58.905 ;
      RECT 54.25 16.065 54.42 16.235 ;
      RECT 54.25 26.945 54.42 27.115 ;
      RECT 53.965 9.775 54.135 9.945 ;
      RECT 53.965 12.495 54.135 12.665 ;
      RECT 53.965 13.345 54.135 13.515 ;
      RECT 53.965 15.215 54.135 15.385 ;
      RECT 53.965 17.935 54.135 18.105 ;
      RECT 53.965 18.445 54.135 18.615 ;
      RECT 53.965 20.655 54.135 20.825 ;
      RECT 53.965 23.375 54.135 23.545 ;
      RECT 53.965 26.095 54.135 26.265 ;
      RECT 53.965 28.815 54.135 28.985 ;
      RECT 53.965 31.535 54.135 31.705 ;
      RECT 53.965 34.255 54.135 34.425 ;
      RECT 53.965 36.975 54.135 37.145 ;
      RECT 53.965 39.695 54.135 39.865 ;
      RECT 53.965 42.415 54.135 42.585 ;
      RECT 53.965 45.135 54.135 45.305 ;
      RECT 53.965 47.855 54.135 48.025 ;
      RECT 53.965 50.575 54.135 50.745 ;
      RECT 53.965 53.295 54.135 53.465 ;
      RECT 53.965 56.015 54.135 56.185 ;
      RECT 53.965 58.735 54.135 58.905 ;
      RECT 53.735 16.405 53.905 16.575 ;
      RECT 53.735 27.285 53.905 27.455 ;
      RECT 53.505 9.775 53.675 9.945 ;
      RECT 53.505 12.495 53.675 12.665 ;
      RECT 53.505 15.215 53.675 15.385 ;
      RECT 53.505 17.935 53.675 18.105 ;
      RECT 53.505 20.655 53.675 20.825 ;
      RECT 53.505 23.375 53.675 23.545 ;
      RECT 53.505 26.095 53.675 26.265 ;
      RECT 53.505 28.815 53.675 28.985 ;
      RECT 53.505 31.535 53.675 31.705 ;
      RECT 53.505 34.255 53.675 34.425 ;
      RECT 53.505 36.975 53.675 37.145 ;
      RECT 53.505 39.695 53.675 39.865 ;
      RECT 53.505 42.415 53.675 42.585 ;
      RECT 53.505 45.135 53.675 45.305 ;
      RECT 53.505 47.855 53.675 48.025 ;
      RECT 53.505 50.575 53.675 50.745 ;
      RECT 53.505 53.295 53.675 53.465 ;
      RECT 53.505 56.015 53.675 56.185 ;
      RECT 53.505 58.735 53.675 58.905 ;
      RECT 53.275 13.685 53.445 13.855 ;
      RECT 53.045 9.775 53.215 9.945 ;
      RECT 53.045 12.495 53.215 12.665 ;
      RECT 53.045 15.215 53.215 15.385 ;
      RECT 53.045 17.935 53.215 18.105 ;
      RECT 53.045 20.655 53.215 20.825 ;
      RECT 53.045 23.375 53.215 23.545 ;
      RECT 53.045 26.095 53.215 26.265 ;
      RECT 53.045 28.815 53.215 28.985 ;
      RECT 53.045 31.535 53.215 31.705 ;
      RECT 53.045 34.255 53.215 34.425 ;
      RECT 53.045 36.975 53.215 37.145 ;
      RECT 53.045 39.695 53.215 39.865 ;
      RECT 53.045 42.415 53.215 42.585 ;
      RECT 53.045 45.135 53.215 45.305 ;
      RECT 53.045 47.855 53.215 48.025 ;
      RECT 53.045 50.575 53.215 50.745 ;
      RECT 53.045 53.295 53.215 53.465 ;
      RECT 53.045 56.015 53.215 56.185 ;
      RECT 53.045 58.735 53.215 58.905 ;
      RECT 52.97 27.965 53.14 28.135 ;
      RECT 52.89 17.085 53.06 17.255 ;
      RECT 52.585 9.775 52.755 9.945 ;
      RECT 52.585 12.495 52.755 12.665 ;
      RECT 52.585 14.705 52.755 14.875 ;
      RECT 52.585 15.215 52.755 15.385 ;
      RECT 52.585 17.935 52.755 18.105 ;
      RECT 52.585 20.655 52.755 20.825 ;
      RECT 52.585 23.375 52.755 23.545 ;
      RECT 52.585 26.095 52.755 26.265 ;
      RECT 52.585 28.815 52.755 28.985 ;
      RECT 52.585 31.535 52.755 31.705 ;
      RECT 52.585 34.255 52.755 34.425 ;
      RECT 52.585 36.975 52.755 37.145 ;
      RECT 52.585 39.695 52.755 39.865 ;
      RECT 52.585 42.415 52.755 42.585 ;
      RECT 52.585 45.135 52.755 45.305 ;
      RECT 52.585 47.855 52.755 48.025 ;
      RECT 52.585 50.575 52.755 50.745 ;
      RECT 52.585 53.295 52.755 53.465 ;
      RECT 52.585 56.015 52.755 56.185 ;
      RECT 52.585 58.735 52.755 58.905 ;
      RECT 52.545 16.405 52.715 16.575 ;
      RECT 52.545 27.285 52.715 27.455 ;
      RECT 52.15 16.065 52.32 16.235 ;
      RECT 52.15 26.945 52.32 27.115 ;
      RECT 52.125 9.775 52.295 9.945 ;
      RECT 52.125 12.495 52.295 12.665 ;
      RECT 52.125 15.215 52.295 15.385 ;
      RECT 52.125 17.935 52.295 18.105 ;
      RECT 52.125 20.655 52.295 20.825 ;
      RECT 52.125 23.375 52.295 23.545 ;
      RECT 52.125 26.095 52.295 26.265 ;
      RECT 52.125 28.815 52.295 28.985 ;
      RECT 52.125 31.535 52.295 31.705 ;
      RECT 52.125 34.255 52.295 34.425 ;
      RECT 52.125 36.975 52.295 37.145 ;
      RECT 52.125 39.695 52.295 39.865 ;
      RECT 52.125 42.415 52.295 42.585 ;
      RECT 52.125 45.135 52.295 45.305 ;
      RECT 52.125 47.855 52.295 48.025 ;
      RECT 52.125 50.575 52.295 50.745 ;
      RECT 52.125 53.295 52.295 53.465 ;
      RECT 52.125 56.015 52.295 56.185 ;
      RECT 52.125 58.735 52.295 58.905 ;
      RECT 51.665 9.775 51.835 9.945 ;
      RECT 51.665 12.495 51.835 12.665 ;
      RECT 51.665 15.215 51.835 15.385 ;
      RECT 51.665 16.745 51.835 16.915 ;
      RECT 51.665 17.935 51.835 18.105 ;
      RECT 51.665 20.655 51.835 20.825 ;
      RECT 51.665 23.375 51.835 23.545 ;
      RECT 51.665 26.095 51.835 26.265 ;
      RECT 51.665 27.625 51.835 27.795 ;
      RECT 51.665 28.815 51.835 28.985 ;
      RECT 51.665 31.535 51.835 31.705 ;
      RECT 51.665 34.255 51.835 34.425 ;
      RECT 51.665 36.975 51.835 37.145 ;
      RECT 51.665 39.695 51.835 39.865 ;
      RECT 51.665 42.415 51.835 42.585 ;
      RECT 51.665 45.135 51.835 45.305 ;
      RECT 51.665 47.855 51.835 48.025 ;
      RECT 51.665 50.575 51.835 50.745 ;
      RECT 51.665 53.295 51.835 53.465 ;
      RECT 51.665 56.015 51.835 56.185 ;
      RECT 51.665 58.735 51.835 58.905 ;
      RECT 51.655 19.465 51.825 19.635 ;
      RECT 51.22 19.805 51.39 19.975 ;
      RECT 51.205 9.775 51.375 9.945 ;
      RECT 51.205 12.495 51.375 12.665 ;
      RECT 51.205 15.215 51.375 15.385 ;
      RECT 51.205 17.935 51.375 18.105 ;
      RECT 51.205 20.655 51.375 20.825 ;
      RECT 51.205 23.375 51.375 23.545 ;
      RECT 51.205 26.095 51.375 26.265 ;
      RECT 51.205 28.815 51.375 28.985 ;
      RECT 51.205 31.535 51.375 31.705 ;
      RECT 51.205 34.255 51.375 34.425 ;
      RECT 51.205 36.975 51.375 37.145 ;
      RECT 51.205 39.695 51.375 39.865 ;
      RECT 51.205 42.415 51.375 42.585 ;
      RECT 51.205 45.135 51.375 45.305 ;
      RECT 51.205 47.855 51.375 48.025 ;
      RECT 51.205 50.575 51.375 50.745 ;
      RECT 51.205 53.295 51.375 53.465 ;
      RECT 51.205 56.015 51.375 56.185 ;
      RECT 51.205 58.735 51.375 58.905 ;
      RECT 50.745 9.775 50.915 9.945 ;
      RECT 50.745 12.495 50.915 12.665 ;
      RECT 50.745 15.215 50.915 15.385 ;
      RECT 50.745 17.935 50.915 18.105 ;
      RECT 50.745 20.655 50.915 20.825 ;
      RECT 50.745 23.375 50.915 23.545 ;
      RECT 50.745 26.095 50.915 26.265 ;
      RECT 50.745 28.815 50.915 28.985 ;
      RECT 50.745 31.535 50.915 31.705 ;
      RECT 50.745 34.255 50.915 34.425 ;
      RECT 50.745 36.975 50.915 37.145 ;
      RECT 50.745 39.695 50.915 39.865 ;
      RECT 50.745 42.415 50.915 42.585 ;
      RECT 50.745 45.135 50.915 45.305 ;
      RECT 50.745 47.855 50.915 48.025 ;
      RECT 50.745 50.575 50.915 50.745 ;
      RECT 50.745 53.295 50.915 53.465 ;
      RECT 50.745 56.015 50.915 56.185 ;
      RECT 50.745 58.735 50.915 58.905 ;
      RECT 50.285 9.775 50.455 9.945 ;
      RECT 50.285 12.495 50.455 12.665 ;
      RECT 50.285 15.215 50.455 15.385 ;
      RECT 50.285 17.935 50.455 18.105 ;
      RECT 50.285 20.655 50.455 20.825 ;
      RECT 50.285 23.375 50.455 23.545 ;
      RECT 50.285 26.095 50.455 26.265 ;
      RECT 50.285 28.815 50.455 28.985 ;
      RECT 50.285 31.535 50.455 31.705 ;
      RECT 50.285 34.255 50.455 34.425 ;
      RECT 50.285 36.975 50.455 37.145 ;
      RECT 50.285 39.695 50.455 39.865 ;
      RECT 50.285 42.415 50.455 42.585 ;
      RECT 50.285 45.135 50.455 45.305 ;
      RECT 50.285 47.855 50.455 48.025 ;
      RECT 50.285 50.575 50.455 50.745 ;
      RECT 50.285 53.295 50.455 53.465 ;
      RECT 50.285 56.015 50.455 56.185 ;
      RECT 50.285 58.735 50.455 58.905 ;
      RECT 49.825 9.775 49.995 9.945 ;
      RECT 49.825 12.495 49.995 12.665 ;
      RECT 49.825 15.215 49.995 15.385 ;
      RECT 49.825 17.935 49.995 18.105 ;
      RECT 49.825 20.655 49.995 20.825 ;
      RECT 49.825 23.375 49.995 23.545 ;
      RECT 49.825 26.095 49.995 26.265 ;
      RECT 49.825 28.815 49.995 28.985 ;
      RECT 49.825 31.535 49.995 31.705 ;
      RECT 49.825 34.255 49.995 34.425 ;
      RECT 49.825 36.975 49.995 37.145 ;
      RECT 49.825 39.695 49.995 39.865 ;
      RECT 49.825 42.415 49.995 42.585 ;
      RECT 49.825 45.135 49.995 45.305 ;
      RECT 49.825 47.855 49.995 48.025 ;
      RECT 49.825 50.575 49.995 50.745 ;
      RECT 49.825 53.295 49.995 53.465 ;
      RECT 49.825 56.015 49.995 56.185 ;
      RECT 49.825 58.735 49.995 58.905 ;
      RECT 49.65 19.805 49.82 19.975 ;
      RECT 49.365 9.775 49.535 9.945 ;
      RECT 49.365 12.495 49.535 12.665 ;
      RECT 49.365 14.705 49.535 14.875 ;
      RECT 49.365 15.215 49.535 15.385 ;
      RECT 49.365 17.935 49.535 18.105 ;
      RECT 49.365 20.655 49.535 20.825 ;
      RECT 49.365 23.375 49.535 23.545 ;
      RECT 49.365 24.565 49.535 24.735 ;
      RECT 49.365 26.095 49.535 26.265 ;
      RECT 49.365 28.815 49.535 28.985 ;
      RECT 49.365 31.535 49.535 31.705 ;
      RECT 49.365 34.255 49.535 34.425 ;
      RECT 49.365 36.975 49.535 37.145 ;
      RECT 49.365 39.695 49.535 39.865 ;
      RECT 49.365 42.415 49.535 42.585 ;
      RECT 49.365 45.135 49.535 45.305 ;
      RECT 49.365 47.855 49.535 48.025 ;
      RECT 49.365 50.575 49.535 50.745 ;
      RECT 49.365 53.295 49.535 53.465 ;
      RECT 49.365 56.015 49.535 56.185 ;
      RECT 49.365 58.735 49.535 58.905 ;
      RECT 49.135 19.465 49.305 19.635 ;
      RECT 48.905 9.775 49.075 9.945 ;
      RECT 48.905 12.495 49.075 12.665 ;
      RECT 48.905 15.215 49.075 15.385 ;
      RECT 48.905 17.935 49.075 18.105 ;
      RECT 48.905 20.655 49.075 20.825 ;
      RECT 48.905 23.375 49.075 23.545 ;
      RECT 48.905 26.095 49.075 26.265 ;
      RECT 48.905 28.815 49.075 28.985 ;
      RECT 48.905 31.535 49.075 31.705 ;
      RECT 48.905 34.255 49.075 34.425 ;
      RECT 48.905 36.975 49.075 37.145 ;
      RECT 48.905 39.695 49.075 39.865 ;
      RECT 48.905 42.415 49.075 42.585 ;
      RECT 48.905 45.135 49.075 45.305 ;
      RECT 48.905 47.855 49.075 48.025 ;
      RECT 48.905 50.575 49.075 50.745 ;
      RECT 48.905 53.295 49.075 53.465 ;
      RECT 48.905 56.015 49.075 56.185 ;
      RECT 48.905 58.735 49.075 58.905 ;
      RECT 48.675 13.685 48.845 13.855 ;
      RECT 48.445 9.775 48.615 9.945 ;
      RECT 48.445 12.495 48.615 12.665 ;
      RECT 48.445 15.215 48.615 15.385 ;
      RECT 48.445 17.935 48.615 18.105 ;
      RECT 48.445 20.655 48.615 20.825 ;
      RECT 48.445 23.375 48.615 23.545 ;
      RECT 48.445 26.095 48.615 26.265 ;
      RECT 48.445 28.815 48.615 28.985 ;
      RECT 48.445 31.535 48.615 31.705 ;
      RECT 48.445 34.255 48.615 34.425 ;
      RECT 48.445 36.975 48.615 37.145 ;
      RECT 48.445 39.695 48.615 39.865 ;
      RECT 48.445 42.415 48.615 42.585 ;
      RECT 48.445 45.135 48.615 45.305 ;
      RECT 48.445 47.855 48.615 48.025 ;
      RECT 48.445 50.575 48.615 50.745 ;
      RECT 48.445 53.295 48.615 53.465 ;
      RECT 48.445 56.015 48.615 56.185 ;
      RECT 48.445 58.735 48.615 58.905 ;
      RECT 48.37 18.785 48.54 18.955 ;
      RECT 47.985 9.775 48.155 9.945 ;
      RECT 47.985 12.495 48.155 12.665 ;
      RECT 47.985 13.345 48.155 13.515 ;
      RECT 47.985 15.215 48.155 15.385 ;
      RECT 47.985 17.935 48.155 18.105 ;
      RECT 47.985 20.655 48.155 20.825 ;
      RECT 47.985 23.375 48.155 23.545 ;
      RECT 47.985 26.095 48.155 26.265 ;
      RECT 47.985 28.815 48.155 28.985 ;
      RECT 47.985 31.535 48.155 31.705 ;
      RECT 47.985 34.255 48.155 34.425 ;
      RECT 47.985 36.975 48.155 37.145 ;
      RECT 47.985 39.695 48.155 39.865 ;
      RECT 47.985 42.415 48.155 42.585 ;
      RECT 47.985 45.135 48.155 45.305 ;
      RECT 47.985 47.855 48.155 48.025 ;
      RECT 47.985 50.575 48.155 50.745 ;
      RECT 47.985 53.295 48.155 53.465 ;
      RECT 47.985 56.015 48.155 56.185 ;
      RECT 47.985 58.735 48.155 58.905 ;
      RECT 47.945 19.465 48.115 19.635 ;
      RECT 47.55 19.805 47.72 19.975 ;
      RECT 47.525 9.775 47.695 9.945 ;
      RECT 47.525 11.305 47.695 11.475 ;
      RECT 47.525 12.495 47.695 12.665 ;
      RECT 47.525 13.685 47.695 13.855 ;
      RECT 47.525 15.215 47.695 15.385 ;
      RECT 47.525 17.935 47.695 18.105 ;
      RECT 47.525 20.655 47.695 20.825 ;
      RECT 47.525 23.375 47.695 23.545 ;
      RECT 47.525 26.095 47.695 26.265 ;
      RECT 47.525 28.815 47.695 28.985 ;
      RECT 47.525 31.535 47.695 31.705 ;
      RECT 47.525 34.255 47.695 34.425 ;
      RECT 47.525 36.975 47.695 37.145 ;
      RECT 47.525 39.695 47.695 39.865 ;
      RECT 47.525 42.415 47.695 42.585 ;
      RECT 47.525 45.135 47.695 45.305 ;
      RECT 47.525 47.855 47.695 48.025 ;
      RECT 47.525 50.575 47.695 50.745 ;
      RECT 47.525 53.295 47.695 53.465 ;
      RECT 47.525 56.015 47.695 56.185 ;
      RECT 47.525 58.735 47.695 58.905 ;
      RECT 47.065 9.775 47.235 9.945 ;
      RECT 47.065 12.495 47.235 12.665 ;
      RECT 47.065 15.215 47.235 15.385 ;
      RECT 47.065 17.935 47.235 18.105 ;
      RECT 47.065 19.125 47.235 19.295 ;
      RECT 47.065 20.655 47.235 20.825 ;
      RECT 47.065 23.375 47.235 23.545 ;
      RECT 47.065 26.095 47.235 26.265 ;
      RECT 47.065 28.815 47.235 28.985 ;
      RECT 47.065 31.535 47.235 31.705 ;
      RECT 47.065 34.255 47.235 34.425 ;
      RECT 47.065 36.975 47.235 37.145 ;
      RECT 47.065 39.695 47.235 39.865 ;
      RECT 47.065 42.415 47.235 42.585 ;
      RECT 47.065 45.135 47.235 45.305 ;
      RECT 47.065 47.855 47.235 48.025 ;
      RECT 47.065 50.575 47.235 50.745 ;
      RECT 47.065 53.295 47.235 53.465 ;
      RECT 47.065 56.015 47.235 56.185 ;
      RECT 47.065 58.735 47.235 58.905 ;
      RECT 46.745 13.685 46.915 13.855 ;
      RECT 46.605 9.775 46.775 9.945 ;
      RECT 46.605 12.495 46.775 12.665 ;
      RECT 46.605 15.215 46.775 15.385 ;
      RECT 46.605 17.935 46.775 18.105 ;
      RECT 46.605 20.655 46.775 20.825 ;
      RECT 46.605 23.375 46.775 23.545 ;
      RECT 46.605 26.095 46.775 26.265 ;
      RECT 46.605 28.815 46.775 28.985 ;
      RECT 46.605 31.535 46.775 31.705 ;
      RECT 46.605 34.255 46.775 34.425 ;
      RECT 46.605 36.975 46.775 37.145 ;
      RECT 46.605 39.695 46.775 39.865 ;
      RECT 46.605 42.415 46.775 42.585 ;
      RECT 46.605 45.135 46.775 45.305 ;
      RECT 46.605 47.855 46.775 48.025 ;
      RECT 46.605 50.575 46.775 50.745 ;
      RECT 46.605 53.295 46.775 53.465 ;
      RECT 46.605 56.015 46.775 56.185 ;
      RECT 46.605 58.735 46.775 58.905 ;
      RECT 46.145 9.775 46.315 9.945 ;
      RECT 46.145 12.495 46.315 12.665 ;
      RECT 46.145 13.685 46.315 13.855 ;
      RECT 46.145 15.215 46.315 15.385 ;
      RECT 46.145 17.935 46.315 18.105 ;
      RECT 46.145 20.655 46.315 20.825 ;
      RECT 46.145 23.375 46.315 23.545 ;
      RECT 46.145 26.095 46.315 26.265 ;
      RECT 46.145 28.815 46.315 28.985 ;
      RECT 46.145 31.535 46.315 31.705 ;
      RECT 46.145 34.255 46.315 34.425 ;
      RECT 46.145 36.975 46.315 37.145 ;
      RECT 46.145 39.695 46.315 39.865 ;
      RECT 46.145 42.415 46.315 42.585 ;
      RECT 46.145 45.135 46.315 45.305 ;
      RECT 46.145 47.855 46.315 48.025 ;
      RECT 46.145 50.575 46.315 50.745 ;
      RECT 46.145 53.295 46.315 53.465 ;
      RECT 46.145 56.015 46.315 56.185 ;
      RECT 46.145 58.735 46.315 58.905 ;
      RECT 45.685 9.775 45.855 9.945 ;
      RECT 45.685 12.495 45.855 12.665 ;
      RECT 45.685 15.215 45.855 15.385 ;
      RECT 45.685 17.935 45.855 18.105 ;
      RECT 45.685 20.655 45.855 20.825 ;
      RECT 45.685 23.375 45.855 23.545 ;
      RECT 45.685 26.095 45.855 26.265 ;
      RECT 45.685 28.815 45.855 28.985 ;
      RECT 45.685 31.535 45.855 31.705 ;
      RECT 45.685 34.255 45.855 34.425 ;
      RECT 45.685 36.975 45.855 37.145 ;
      RECT 45.685 39.695 45.855 39.865 ;
      RECT 45.685 42.415 45.855 42.585 ;
      RECT 45.685 45.135 45.855 45.305 ;
      RECT 45.685 47.855 45.855 48.025 ;
      RECT 45.685 50.575 45.855 50.745 ;
      RECT 45.685 53.295 45.855 53.465 ;
      RECT 45.685 56.015 45.855 56.185 ;
      RECT 45.685 58.735 45.855 58.905 ;
      RECT 45.225 9.775 45.395 9.945 ;
      RECT 45.225 12.495 45.395 12.665 ;
      RECT 45.225 15.215 45.395 15.385 ;
      RECT 45.225 17.935 45.395 18.105 ;
      RECT 45.225 20.655 45.395 20.825 ;
      RECT 45.225 23.375 45.395 23.545 ;
      RECT 45.225 26.095 45.395 26.265 ;
      RECT 45.225 28.815 45.395 28.985 ;
      RECT 45.225 31.535 45.395 31.705 ;
      RECT 45.225 34.255 45.395 34.425 ;
      RECT 45.225 36.975 45.395 37.145 ;
      RECT 45.225 39.695 45.395 39.865 ;
      RECT 45.225 42.415 45.395 42.585 ;
      RECT 45.225 45.135 45.395 45.305 ;
      RECT 45.225 47.855 45.395 48.025 ;
      RECT 45.225 50.575 45.395 50.745 ;
      RECT 45.225 53.295 45.395 53.465 ;
      RECT 45.225 56.015 45.395 56.185 ;
      RECT 45.225 58.735 45.395 58.905 ;
      RECT 44.765 9.775 44.935 9.945 ;
      RECT 44.765 12.495 44.935 12.665 ;
      RECT 44.765 15.215 44.935 15.385 ;
      RECT 44.765 17.935 44.935 18.105 ;
      RECT 44.765 20.655 44.935 20.825 ;
      RECT 44.765 23.375 44.935 23.545 ;
      RECT 44.765 26.095 44.935 26.265 ;
      RECT 44.765 28.815 44.935 28.985 ;
      RECT 44.765 31.535 44.935 31.705 ;
      RECT 44.765 34.255 44.935 34.425 ;
      RECT 44.765 36.975 44.935 37.145 ;
      RECT 44.765 39.695 44.935 39.865 ;
      RECT 44.765 42.415 44.935 42.585 ;
      RECT 44.765 45.135 44.935 45.305 ;
      RECT 44.765 47.855 44.935 48.025 ;
      RECT 44.765 50.575 44.935 50.745 ;
      RECT 44.765 53.295 44.935 53.465 ;
      RECT 44.765 56.015 44.935 56.185 ;
      RECT 44.765 58.735 44.935 58.905 ;
      RECT 44.305 9.775 44.475 9.945 ;
      RECT 44.305 12.495 44.475 12.665 ;
      RECT 44.305 15.215 44.475 15.385 ;
      RECT 44.305 17.935 44.475 18.105 ;
      RECT 44.305 20.655 44.475 20.825 ;
      RECT 44.305 23.375 44.475 23.545 ;
      RECT 44.305 26.095 44.475 26.265 ;
      RECT 44.305 28.815 44.475 28.985 ;
      RECT 44.305 31.535 44.475 31.705 ;
      RECT 44.305 34.255 44.475 34.425 ;
      RECT 44.305 36.975 44.475 37.145 ;
      RECT 44.305 39.695 44.475 39.865 ;
      RECT 44.305 42.415 44.475 42.585 ;
      RECT 44.305 45.135 44.475 45.305 ;
      RECT 44.305 47.855 44.475 48.025 ;
      RECT 44.305 50.575 44.475 50.745 ;
      RECT 44.305 53.295 44.475 53.465 ;
      RECT 44.305 56.015 44.475 56.185 ;
      RECT 44.305 58.735 44.475 58.905 ;
      RECT 43.845 9.775 44.015 9.945 ;
      RECT 43.845 12.495 44.015 12.665 ;
      RECT 43.845 15.215 44.015 15.385 ;
      RECT 43.845 17.935 44.015 18.105 ;
      RECT 43.845 20.655 44.015 20.825 ;
      RECT 43.845 22.865 44.015 23.035 ;
      RECT 43.845 23.375 44.015 23.545 ;
      RECT 43.845 26.095 44.015 26.265 ;
      RECT 43.845 26.945 44.015 27.115 ;
      RECT 43.845 28.815 44.015 28.985 ;
      RECT 43.845 31.535 44.015 31.705 ;
      RECT 43.845 34.255 44.015 34.425 ;
      RECT 43.845 36.975 44.015 37.145 ;
      RECT 43.845 39.695 44.015 39.865 ;
      RECT 43.845 42.415 44.015 42.585 ;
      RECT 43.845 45.135 44.015 45.305 ;
      RECT 43.845 47.855 44.015 48.025 ;
      RECT 43.845 50.575 44.015 50.745 ;
      RECT 43.845 53.295 44.015 53.465 ;
      RECT 43.845 56.015 44.015 56.185 ;
      RECT 43.845 58.735 44.015 58.905 ;
      RECT 43.385 9.775 43.555 9.945 ;
      RECT 43.385 12.495 43.555 12.665 ;
      RECT 43.385 15.215 43.555 15.385 ;
      RECT 43.385 17.935 43.555 18.105 ;
      RECT 43.385 20.655 43.555 20.825 ;
      RECT 43.385 23.375 43.555 23.545 ;
      RECT 43.385 26.095 43.555 26.265 ;
      RECT 43.385 28.815 43.555 28.985 ;
      RECT 43.385 31.535 43.555 31.705 ;
      RECT 43.385 34.255 43.555 34.425 ;
      RECT 43.385 36.975 43.555 37.145 ;
      RECT 43.385 39.695 43.555 39.865 ;
      RECT 43.385 42.415 43.555 42.585 ;
      RECT 43.385 45.135 43.555 45.305 ;
      RECT 43.385 47.855 43.555 48.025 ;
      RECT 43.385 50.575 43.555 50.745 ;
      RECT 43.385 53.295 43.555 53.465 ;
      RECT 43.385 56.015 43.555 56.185 ;
      RECT 43.385 58.735 43.555 58.905 ;
      RECT 42.925 9.775 43.095 9.945 ;
      RECT 42.925 12.495 43.095 12.665 ;
      RECT 42.925 15.215 43.095 15.385 ;
      RECT 42.925 17.935 43.095 18.105 ;
      RECT 42.925 20.655 43.095 20.825 ;
      RECT 42.925 23.375 43.095 23.545 ;
      RECT 42.925 26.095 43.095 26.265 ;
      RECT 42.925 28.815 43.095 28.985 ;
      RECT 42.925 31.535 43.095 31.705 ;
      RECT 42.925 34.255 43.095 34.425 ;
      RECT 42.925 36.975 43.095 37.145 ;
      RECT 42.925 39.695 43.095 39.865 ;
      RECT 42.925 42.415 43.095 42.585 ;
      RECT 42.925 45.135 43.095 45.305 ;
      RECT 42.925 47.855 43.095 48.025 ;
      RECT 42.925 50.575 43.095 50.745 ;
      RECT 42.925 53.295 43.095 53.465 ;
      RECT 42.925 56.015 43.095 56.185 ;
      RECT 42.925 58.735 43.095 58.905 ;
      RECT 42.465 9.775 42.635 9.945 ;
      RECT 42.465 12.495 42.635 12.665 ;
      RECT 42.465 15.215 42.635 15.385 ;
      RECT 42.465 17.935 42.635 18.105 ;
      RECT 42.465 20.655 42.635 20.825 ;
      RECT 42.465 23.375 42.635 23.545 ;
      RECT 42.465 26.095 42.635 26.265 ;
      RECT 42.465 28.815 42.635 28.985 ;
      RECT 42.465 31.535 42.635 31.705 ;
      RECT 42.465 34.255 42.635 34.425 ;
      RECT 42.465 36.975 42.635 37.145 ;
      RECT 42.465 39.695 42.635 39.865 ;
      RECT 42.465 42.415 42.635 42.585 ;
      RECT 42.465 45.135 42.635 45.305 ;
      RECT 42.465 47.855 42.635 48.025 ;
      RECT 42.465 50.575 42.635 50.745 ;
      RECT 42.465 53.295 42.635 53.465 ;
      RECT 42.465 56.015 42.635 56.185 ;
      RECT 42.465 58.735 42.635 58.905 ;
      RECT 42.005 9.775 42.175 9.945 ;
      RECT 42.005 12.495 42.175 12.665 ;
      RECT 42.005 15.215 42.175 15.385 ;
      RECT 42.005 17.935 42.175 18.105 ;
      RECT 42.005 20.655 42.175 20.825 ;
      RECT 42.005 23.375 42.175 23.545 ;
      RECT 42.005 26.095 42.175 26.265 ;
      RECT 42.005 28.815 42.175 28.985 ;
      RECT 42.005 31.535 42.175 31.705 ;
      RECT 42.005 34.255 42.175 34.425 ;
      RECT 42.005 36.975 42.175 37.145 ;
      RECT 42.005 39.695 42.175 39.865 ;
      RECT 42.005 42.415 42.175 42.585 ;
      RECT 42.005 45.135 42.175 45.305 ;
      RECT 42.005 47.855 42.175 48.025 ;
      RECT 42.005 50.575 42.175 50.745 ;
      RECT 42.005 53.295 42.175 53.465 ;
      RECT 42.005 56.015 42.175 56.185 ;
      RECT 42.005 58.735 42.175 58.905 ;
      RECT 41.545 9.775 41.715 9.945 ;
      RECT 41.545 12.495 41.715 12.665 ;
      RECT 41.545 15.215 41.715 15.385 ;
      RECT 41.545 17.935 41.715 18.105 ;
      RECT 41.545 20.655 41.715 20.825 ;
      RECT 41.545 23.375 41.715 23.545 ;
      RECT 41.545 26.095 41.715 26.265 ;
      RECT 41.545 28.815 41.715 28.985 ;
      RECT 41.545 31.535 41.715 31.705 ;
      RECT 41.545 34.255 41.715 34.425 ;
      RECT 41.545 36.975 41.715 37.145 ;
      RECT 41.545 39.695 41.715 39.865 ;
      RECT 41.545 42.415 41.715 42.585 ;
      RECT 41.545 45.135 41.715 45.305 ;
      RECT 41.545 47.855 41.715 48.025 ;
      RECT 41.545 50.575 41.715 50.745 ;
      RECT 41.545 53.295 41.715 53.465 ;
      RECT 41.545 56.015 41.715 56.185 ;
      RECT 41.545 58.735 41.715 58.905 ;
      RECT 41.535 27.285 41.705 27.455 ;
      RECT 41.1 26.945 41.27 27.115 ;
      RECT 41.085 9.775 41.255 9.945 ;
      RECT 41.085 12.495 41.255 12.665 ;
      RECT 41.085 15.215 41.255 15.385 ;
      RECT 41.085 17.935 41.255 18.105 ;
      RECT 41.085 20.655 41.255 20.825 ;
      RECT 41.085 23.375 41.255 23.545 ;
      RECT 41.085 26.095 41.255 26.265 ;
      RECT 41.085 28.815 41.255 28.985 ;
      RECT 41.085 31.535 41.255 31.705 ;
      RECT 41.085 34.255 41.255 34.425 ;
      RECT 41.085 36.975 41.255 37.145 ;
      RECT 41.085 39.695 41.255 39.865 ;
      RECT 41.085 42.415 41.255 42.585 ;
      RECT 41.085 45.135 41.255 45.305 ;
      RECT 41.085 47.855 41.255 48.025 ;
      RECT 41.085 50.575 41.255 50.745 ;
      RECT 41.085 53.295 41.255 53.465 ;
      RECT 41.085 56.015 41.255 56.185 ;
      RECT 41.085 58.735 41.255 58.905 ;
      RECT 40.625 9.775 40.795 9.945 ;
      RECT 40.625 12.495 40.795 12.665 ;
      RECT 40.625 15.215 40.795 15.385 ;
      RECT 40.625 17.935 40.795 18.105 ;
      RECT 40.625 18.445 40.795 18.615 ;
      RECT 40.625 20.655 40.795 20.825 ;
      RECT 40.625 23.375 40.795 23.545 ;
      RECT 40.625 26.095 40.795 26.265 ;
      RECT 40.625 28.815 40.795 28.985 ;
      RECT 40.625 31.535 40.795 31.705 ;
      RECT 40.625 34.255 40.795 34.425 ;
      RECT 40.625 36.975 40.795 37.145 ;
      RECT 40.625 39.695 40.795 39.865 ;
      RECT 40.625 42.415 40.795 42.585 ;
      RECT 40.625 45.135 40.795 45.305 ;
      RECT 40.625 47.855 40.795 48.025 ;
      RECT 40.625 50.575 40.795 50.745 ;
      RECT 40.625 53.295 40.795 53.465 ;
      RECT 40.625 56.015 40.795 56.185 ;
      RECT 40.625 58.735 40.795 58.905 ;
      RECT 40.165 9.775 40.335 9.945 ;
      RECT 40.165 12.495 40.335 12.665 ;
      RECT 40.165 15.215 40.335 15.385 ;
      RECT 40.165 15.725 40.335 15.895 ;
      RECT 40.165 17.935 40.335 18.105 ;
      RECT 40.165 20.655 40.335 20.825 ;
      RECT 40.165 23.375 40.335 23.545 ;
      RECT 40.165 26.095 40.335 26.265 ;
      RECT 40.165 28.815 40.335 28.985 ;
      RECT 40.165 31.535 40.335 31.705 ;
      RECT 40.165 34.255 40.335 34.425 ;
      RECT 40.165 34.765 40.335 34.935 ;
      RECT 40.165 36.975 40.335 37.145 ;
      RECT 40.165 39.695 40.335 39.865 ;
      RECT 40.165 42.415 40.335 42.585 ;
      RECT 40.165 45.135 40.335 45.305 ;
      RECT 40.165 47.855 40.335 48.025 ;
      RECT 40.165 50.575 40.335 50.745 ;
      RECT 40.165 53.295 40.335 53.465 ;
      RECT 40.165 56.015 40.335 56.185 ;
      RECT 40.165 58.735 40.335 58.905 ;
      RECT 39.705 9.775 39.875 9.945 ;
      RECT 39.705 12.495 39.875 12.665 ;
      RECT 39.705 15.215 39.875 15.385 ;
      RECT 39.705 17.935 39.875 18.105 ;
      RECT 39.705 20.655 39.875 20.825 ;
      RECT 39.705 23.375 39.875 23.545 ;
      RECT 39.705 26.095 39.875 26.265 ;
      RECT 39.705 28.815 39.875 28.985 ;
      RECT 39.705 31.535 39.875 31.705 ;
      RECT 39.705 34.255 39.875 34.425 ;
      RECT 39.705 36.975 39.875 37.145 ;
      RECT 39.705 39.695 39.875 39.865 ;
      RECT 39.705 42.415 39.875 42.585 ;
      RECT 39.705 45.135 39.875 45.305 ;
      RECT 39.705 47.855 39.875 48.025 ;
      RECT 39.705 50.575 39.875 50.745 ;
      RECT 39.705 53.295 39.875 53.465 ;
      RECT 39.705 56.015 39.875 56.185 ;
      RECT 39.705 58.735 39.875 58.905 ;
      RECT 39.53 26.945 39.7 27.115 ;
      RECT 39.245 9.775 39.415 9.945 ;
      RECT 39.245 12.495 39.415 12.665 ;
      RECT 39.245 15.215 39.415 15.385 ;
      RECT 39.245 17.935 39.415 18.105 ;
      RECT 39.245 20.655 39.415 20.825 ;
      RECT 39.245 23.375 39.415 23.545 ;
      RECT 39.245 26.095 39.415 26.265 ;
      RECT 39.245 28.815 39.415 28.985 ;
      RECT 39.245 31.535 39.415 31.705 ;
      RECT 39.245 34.255 39.415 34.425 ;
      RECT 39.245 36.975 39.415 37.145 ;
      RECT 39.245 39.695 39.415 39.865 ;
      RECT 39.245 42.415 39.415 42.585 ;
      RECT 39.245 45.135 39.415 45.305 ;
      RECT 39.245 47.855 39.415 48.025 ;
      RECT 39.245 50.575 39.415 50.745 ;
      RECT 39.245 53.295 39.415 53.465 ;
      RECT 39.245 56.015 39.415 56.185 ;
      RECT 39.245 58.735 39.415 58.905 ;
      RECT 39.015 27.285 39.185 27.455 ;
      RECT 38.785 9.775 38.955 9.945 ;
      RECT 38.785 12.495 38.955 12.665 ;
      RECT 38.785 15.215 38.955 15.385 ;
      RECT 38.785 17.935 38.955 18.105 ;
      RECT 38.785 20.655 38.955 20.825 ;
      RECT 38.785 23.375 38.955 23.545 ;
      RECT 38.785 26.095 38.955 26.265 ;
      RECT 38.785 28.815 38.955 28.985 ;
      RECT 38.785 31.535 38.955 31.705 ;
      RECT 38.785 34.255 38.955 34.425 ;
      RECT 38.785 36.975 38.955 37.145 ;
      RECT 38.785 39.695 38.955 39.865 ;
      RECT 38.785 42.415 38.955 42.585 ;
      RECT 38.785 45.135 38.955 45.305 ;
      RECT 38.785 47.855 38.955 48.025 ;
      RECT 38.785 50.575 38.955 50.745 ;
      RECT 38.785 53.295 38.955 53.465 ;
      RECT 38.785 56.015 38.955 56.185 ;
      RECT 38.785 58.735 38.955 58.905 ;
      RECT 38.325 9.775 38.495 9.945 ;
      RECT 38.325 12.495 38.495 12.665 ;
      RECT 38.325 14.705 38.495 14.875 ;
      RECT 38.325 15.215 38.495 15.385 ;
      RECT 38.325 17.935 38.495 18.105 ;
      RECT 38.325 20.655 38.495 20.825 ;
      RECT 38.325 23.375 38.495 23.545 ;
      RECT 38.325 25.585 38.495 25.755 ;
      RECT 38.325 26.095 38.495 26.265 ;
      RECT 38.325 28.815 38.495 28.985 ;
      RECT 38.325 29.325 38.495 29.495 ;
      RECT 38.325 31.535 38.495 31.705 ;
      RECT 38.325 33.745 38.495 33.915 ;
      RECT 38.325 34.255 38.495 34.425 ;
      RECT 38.325 36.975 38.495 37.145 ;
      RECT 38.325 39.695 38.495 39.865 ;
      RECT 38.325 42.415 38.495 42.585 ;
      RECT 38.325 45.135 38.495 45.305 ;
      RECT 38.325 47.855 38.495 48.025 ;
      RECT 38.325 50.575 38.495 50.745 ;
      RECT 38.325 53.295 38.495 53.465 ;
      RECT 38.325 56.015 38.495 56.185 ;
      RECT 38.325 58.735 38.495 58.905 ;
      RECT 38.315 19.465 38.485 19.635 ;
      RECT 38.25 27.965 38.42 28.135 ;
      RECT 37.88 19.805 38.05 19.975 ;
      RECT 37.865 9.775 38.035 9.945 ;
      RECT 37.865 12.495 38.035 12.665 ;
      RECT 37.865 15.215 38.035 15.385 ;
      RECT 37.865 17.935 38.035 18.105 ;
      RECT 37.865 20.655 38.035 20.825 ;
      RECT 37.865 23.375 38.035 23.545 ;
      RECT 37.865 26.095 38.035 26.265 ;
      RECT 37.865 28.815 38.035 28.985 ;
      RECT 37.865 31.535 38.035 31.705 ;
      RECT 37.865 34.255 38.035 34.425 ;
      RECT 37.865 36.975 38.035 37.145 ;
      RECT 37.865 39.695 38.035 39.865 ;
      RECT 37.865 42.415 38.035 42.585 ;
      RECT 37.865 45.135 38.035 45.305 ;
      RECT 37.865 47.855 38.035 48.025 ;
      RECT 37.865 50.575 38.035 50.745 ;
      RECT 37.865 53.295 38.035 53.465 ;
      RECT 37.865 56.015 38.035 56.185 ;
      RECT 37.865 58.735 38.035 58.905 ;
      RECT 37.855 16.405 38.025 16.575 ;
      RECT 37.855 35.785 38.025 35.955 ;
      RECT 37.825 27.285 37.995 27.455 ;
      RECT 37.635 13.685 37.805 13.855 ;
      RECT 37.635 24.565 37.805 24.735 ;
      RECT 37.635 30.005 37.805 30.175 ;
      RECT 37.635 33.065 37.805 33.235 ;
      RECT 37.43 26.945 37.6 27.115 ;
      RECT 37.42 16.065 37.59 16.235 ;
      RECT 37.42 36.125 37.59 36.295 ;
      RECT 37.405 9.775 37.575 9.945 ;
      RECT 37.405 12.495 37.575 12.665 ;
      RECT 37.405 15.215 37.575 15.385 ;
      RECT 37.405 17.935 37.575 18.105 ;
      RECT 37.405 20.655 37.575 20.825 ;
      RECT 37.405 23.375 37.575 23.545 ;
      RECT 37.405 26.095 37.575 26.265 ;
      RECT 37.405 28.815 37.575 28.985 ;
      RECT 37.405 31.535 37.575 31.705 ;
      RECT 37.405 34.255 37.575 34.425 ;
      RECT 37.405 36.975 37.575 37.145 ;
      RECT 37.405 39.695 37.575 39.865 ;
      RECT 37.405 42.415 37.575 42.585 ;
      RECT 37.405 45.135 37.575 45.305 ;
      RECT 37.405 47.855 37.575 48.025 ;
      RECT 37.405 50.575 37.575 50.745 ;
      RECT 37.405 53.295 37.575 53.465 ;
      RECT 37.405 56.015 37.575 56.185 ;
      RECT 37.405 58.735 37.575 58.905 ;
      RECT 36.945 9.775 37.115 9.945 ;
      RECT 36.945 12.495 37.115 12.665 ;
      RECT 36.945 13.685 37.115 13.855 ;
      RECT 36.945 15.215 37.115 15.385 ;
      RECT 36.945 17.935 37.115 18.105 ;
      RECT 36.945 20.655 37.115 20.825 ;
      RECT 36.945 23.375 37.115 23.545 ;
      RECT 36.945 24.225 37.115 24.395 ;
      RECT 36.945 26.095 37.115 26.265 ;
      RECT 36.945 27.625 37.115 27.795 ;
      RECT 36.945 28.815 37.115 28.985 ;
      RECT 36.945 29.665 37.115 29.835 ;
      RECT 36.945 31.535 37.115 31.705 ;
      RECT 36.945 33.065 37.115 33.235 ;
      RECT 36.945 34.255 37.115 34.425 ;
      RECT 36.945 36.975 37.115 37.145 ;
      RECT 36.945 39.695 37.115 39.865 ;
      RECT 36.945 42.415 37.115 42.585 ;
      RECT 36.945 45.135 37.115 45.305 ;
      RECT 36.945 47.855 37.115 48.025 ;
      RECT 36.945 50.575 37.115 50.745 ;
      RECT 36.945 53.295 37.115 53.465 ;
      RECT 36.945 56.015 37.115 56.185 ;
      RECT 36.945 58.735 37.115 58.905 ;
      RECT 36.485 9.775 36.655 9.945 ;
      RECT 36.485 10.965 36.655 11.135 ;
      RECT 36.485 12.495 36.655 12.665 ;
      RECT 36.485 13.345 36.655 13.515 ;
      RECT 36.485 15.215 36.655 15.385 ;
      RECT 36.485 17.935 36.655 18.105 ;
      RECT 36.485 20.655 36.655 20.825 ;
      RECT 36.485 23.375 36.655 23.545 ;
      RECT 36.485 24.225 36.655 24.395 ;
      RECT 36.485 26.095 36.655 26.265 ;
      RECT 36.485 28.815 36.655 28.985 ;
      RECT 36.485 29.665 36.655 29.835 ;
      RECT 36.485 31.535 36.655 31.705 ;
      RECT 36.485 33.065 36.655 33.235 ;
      RECT 36.485 34.255 36.655 34.425 ;
      RECT 36.485 36.975 36.655 37.145 ;
      RECT 36.485 39.695 36.655 39.865 ;
      RECT 36.485 42.415 36.655 42.585 ;
      RECT 36.485 45.135 36.655 45.305 ;
      RECT 36.485 47.855 36.655 48.025 ;
      RECT 36.485 50.575 36.655 50.745 ;
      RECT 36.485 53.295 36.655 53.465 ;
      RECT 36.485 56.015 36.655 56.185 ;
      RECT 36.485 58.735 36.655 58.905 ;
      RECT 36.31 19.805 36.48 19.975 ;
      RECT 36.025 9.775 36.195 9.945 ;
      RECT 36.025 11.645 36.195 11.815 ;
      RECT 36.025 12.495 36.195 12.665 ;
      RECT 36.025 15.215 36.195 15.385 ;
      RECT 36.025 17.935 36.195 18.105 ;
      RECT 36.025 20.655 36.195 20.825 ;
      RECT 36.025 23.375 36.195 23.545 ;
      RECT 36.025 26.095 36.195 26.265 ;
      RECT 36.025 28.815 36.195 28.985 ;
      RECT 36.025 31.535 36.195 31.705 ;
      RECT 36.025 34.255 36.195 34.425 ;
      RECT 36.025 36.975 36.195 37.145 ;
      RECT 36.025 39.695 36.195 39.865 ;
      RECT 36.025 42.415 36.195 42.585 ;
      RECT 36.025 45.135 36.195 45.305 ;
      RECT 36.025 47.855 36.195 48.025 ;
      RECT 36.025 50.575 36.195 50.745 ;
      RECT 36.025 53.295 36.195 53.465 ;
      RECT 36.025 56.015 36.195 56.185 ;
      RECT 36.025 58.735 36.195 58.905 ;
      RECT 35.85 16.065 36.02 16.235 ;
      RECT 35.85 36.125 36.02 36.295 ;
      RECT 35.795 13.685 35.965 13.855 ;
      RECT 35.795 19.465 35.965 19.635 ;
      RECT 35.795 24.565 35.965 24.735 ;
      RECT 35.795 30.005 35.965 30.175 ;
      RECT 35.795 33.065 35.965 33.235 ;
      RECT 35.565 9.775 35.735 9.945 ;
      RECT 35.565 11.305 35.735 11.475 ;
      RECT 35.565 12.495 35.735 12.665 ;
      RECT 35.565 15.215 35.735 15.385 ;
      RECT 35.565 17.935 35.735 18.105 ;
      RECT 35.565 20.655 35.735 20.825 ;
      RECT 35.565 23.375 35.735 23.545 ;
      RECT 35.565 26.095 35.735 26.265 ;
      RECT 35.565 28.815 35.735 28.985 ;
      RECT 35.565 31.535 35.735 31.705 ;
      RECT 35.565 34.255 35.735 34.425 ;
      RECT 35.565 36.975 35.735 37.145 ;
      RECT 35.565 39.695 35.735 39.865 ;
      RECT 35.565 42.415 35.735 42.585 ;
      RECT 35.565 45.135 35.735 45.305 ;
      RECT 35.565 47.855 35.735 48.025 ;
      RECT 35.565 50.575 35.735 50.745 ;
      RECT 35.565 53.295 35.735 53.465 ;
      RECT 35.565 56.015 35.735 56.185 ;
      RECT 35.565 58.735 35.735 58.905 ;
      RECT 35.335 16.405 35.505 16.575 ;
      RECT 35.335 35.785 35.505 35.955 ;
      RECT 35.105 9.775 35.275 9.945 ;
      RECT 35.105 10.965 35.275 11.135 ;
      RECT 35.105 12.495 35.275 12.665 ;
      RECT 35.105 13.685 35.275 13.855 ;
      RECT 35.105 15.215 35.275 15.385 ;
      RECT 35.105 17.935 35.275 18.105 ;
      RECT 35.105 20.655 35.275 20.825 ;
      RECT 35.105 22.185 35.275 22.355 ;
      RECT 35.105 23.375 35.275 23.545 ;
      RECT 35.105 24.565 35.275 24.735 ;
      RECT 35.105 26.095 35.275 26.265 ;
      RECT 35.105 28.815 35.275 28.985 ;
      RECT 35.105 30.005 35.275 30.175 ;
      RECT 35.105 31.535 35.275 31.705 ;
      RECT 35.105 33.065 35.275 33.235 ;
      RECT 35.105 34.255 35.275 34.425 ;
      RECT 35.105 36.975 35.275 37.145 ;
      RECT 35.105 39.695 35.275 39.865 ;
      RECT 35.105 42.415 35.275 42.585 ;
      RECT 35.105 45.135 35.275 45.305 ;
      RECT 35.105 47.855 35.275 48.025 ;
      RECT 35.105 50.575 35.275 50.745 ;
      RECT 35.105 53.295 35.275 53.465 ;
      RECT 35.105 56.015 35.275 56.185 ;
      RECT 35.105 58.735 35.275 58.905 ;
      RECT 35.03 18.785 35.2 18.955 ;
      RECT 34.645 9.775 34.815 9.945 ;
      RECT 34.645 10.285 34.815 10.455 ;
      RECT 34.645 12.495 34.815 12.665 ;
      RECT 34.645 15.215 34.815 15.385 ;
      RECT 34.645 17.935 34.815 18.105 ;
      RECT 34.645 20.655 34.815 20.825 ;
      RECT 34.645 23.375 34.815 23.545 ;
      RECT 34.645 26.095 34.815 26.265 ;
      RECT 34.645 28.815 34.815 28.985 ;
      RECT 34.645 31.535 34.815 31.705 ;
      RECT 34.645 34.255 34.815 34.425 ;
      RECT 34.645 36.975 34.815 37.145 ;
      RECT 34.645 39.695 34.815 39.865 ;
      RECT 34.645 42.415 34.815 42.585 ;
      RECT 34.645 45.135 34.815 45.305 ;
      RECT 34.645 47.855 34.815 48.025 ;
      RECT 34.645 50.575 34.815 50.745 ;
      RECT 34.645 53.295 34.815 53.465 ;
      RECT 34.645 56.015 34.815 56.185 ;
      RECT 34.645 58.735 34.815 58.905 ;
      RECT 34.605 19.465 34.775 19.635 ;
      RECT 34.57 16.745 34.74 16.915 ;
      RECT 34.57 35.105 34.74 35.275 ;
      RECT 34.21 19.805 34.38 19.975 ;
      RECT 34.185 9.775 34.355 9.945 ;
      RECT 34.185 12.495 34.355 12.665 ;
      RECT 34.185 15.215 34.355 15.385 ;
      RECT 34.185 17.935 34.355 18.105 ;
      RECT 34.185 20.655 34.355 20.825 ;
      RECT 34.185 23.375 34.355 23.545 ;
      RECT 34.185 26.095 34.355 26.265 ;
      RECT 34.185 28.815 34.355 28.985 ;
      RECT 34.185 31.535 34.355 31.705 ;
      RECT 34.185 34.255 34.355 34.425 ;
      RECT 34.185 36.975 34.355 37.145 ;
      RECT 34.185 39.695 34.355 39.865 ;
      RECT 34.185 42.415 34.355 42.585 ;
      RECT 34.185 45.135 34.355 45.305 ;
      RECT 34.185 47.855 34.355 48.025 ;
      RECT 34.185 50.575 34.355 50.745 ;
      RECT 34.185 53.295 34.355 53.465 ;
      RECT 34.185 56.015 34.355 56.185 ;
      RECT 34.185 58.735 34.355 58.905 ;
      RECT 34.145 16.405 34.315 16.575 ;
      RECT 34.145 35.785 34.315 35.955 ;
      RECT 33.75 16.065 33.92 16.235 ;
      RECT 33.75 36.125 33.92 36.295 ;
      RECT 33.725 9.775 33.895 9.945 ;
      RECT 33.725 11.985 33.895 12.155 ;
      RECT 33.725 12.495 33.895 12.665 ;
      RECT 33.725 15.215 33.895 15.385 ;
      RECT 33.725 17.935 33.895 18.105 ;
      RECT 33.725 19.125 33.895 19.295 ;
      RECT 33.725 20.655 33.895 20.825 ;
      RECT 33.725 23.375 33.895 23.545 ;
      RECT 33.725 26.095 33.895 26.265 ;
      RECT 33.725 28.815 33.895 28.985 ;
      RECT 33.725 31.535 33.895 31.705 ;
      RECT 33.725 34.255 33.895 34.425 ;
      RECT 33.725 36.975 33.895 37.145 ;
      RECT 33.725 39.695 33.895 39.865 ;
      RECT 33.725 42.415 33.895 42.585 ;
      RECT 33.725 45.135 33.895 45.305 ;
      RECT 33.725 47.855 33.895 48.025 ;
      RECT 33.725 50.575 33.895 50.745 ;
      RECT 33.725 53.295 33.895 53.465 ;
      RECT 33.725 56.015 33.895 56.185 ;
      RECT 33.725 58.735 33.895 58.905 ;
      RECT 33.265 9.775 33.435 9.945 ;
      RECT 33.265 12.495 33.435 12.665 ;
      RECT 33.265 15.215 33.435 15.385 ;
      RECT 33.265 16.745 33.435 16.915 ;
      RECT 33.265 17.935 33.435 18.105 ;
      RECT 33.265 20.655 33.435 20.825 ;
      RECT 33.265 23.375 33.435 23.545 ;
      RECT 33.265 26.095 33.435 26.265 ;
      RECT 33.265 28.815 33.435 28.985 ;
      RECT 33.265 31.535 33.435 31.705 ;
      RECT 33.265 34.255 33.435 34.425 ;
      RECT 33.265 35.445 33.435 35.615 ;
      RECT 33.265 36.975 33.435 37.145 ;
      RECT 33.265 39.695 33.435 39.865 ;
      RECT 33.265 42.415 33.435 42.585 ;
      RECT 33.265 45.135 33.435 45.305 ;
      RECT 33.265 47.855 33.435 48.025 ;
      RECT 33.265 50.575 33.435 50.745 ;
      RECT 33.265 53.295 33.435 53.465 ;
      RECT 33.265 56.015 33.435 56.185 ;
      RECT 33.265 58.735 33.435 58.905 ;
      RECT 32.805 9.775 32.975 9.945 ;
      RECT 32.805 12.495 32.975 12.665 ;
      RECT 32.805 15.215 32.975 15.385 ;
      RECT 32.805 17.935 32.975 18.105 ;
      RECT 32.805 20.655 32.975 20.825 ;
      RECT 32.805 23.375 32.975 23.545 ;
      RECT 32.805 26.095 32.975 26.265 ;
      RECT 32.805 28.815 32.975 28.985 ;
      RECT 32.805 31.535 32.975 31.705 ;
      RECT 32.805 34.255 32.975 34.425 ;
      RECT 32.805 36.975 32.975 37.145 ;
      RECT 32.805 39.695 32.975 39.865 ;
      RECT 32.805 42.415 32.975 42.585 ;
      RECT 32.805 45.135 32.975 45.305 ;
      RECT 32.805 47.855 32.975 48.025 ;
      RECT 32.805 50.575 32.975 50.745 ;
      RECT 32.805 53.295 32.975 53.465 ;
      RECT 32.805 56.015 32.975 56.185 ;
      RECT 32.805 58.735 32.975 58.905 ;
      RECT 32.345 9.775 32.515 9.945 ;
      RECT 32.345 12.495 32.515 12.665 ;
      RECT 32.345 15.215 32.515 15.385 ;
      RECT 32.345 17.935 32.515 18.105 ;
      RECT 32.345 20.655 32.515 20.825 ;
      RECT 32.345 23.375 32.515 23.545 ;
      RECT 32.345 26.095 32.515 26.265 ;
      RECT 32.345 28.815 32.515 28.985 ;
      RECT 32.345 31.535 32.515 31.705 ;
      RECT 32.345 34.255 32.515 34.425 ;
      RECT 32.345 36.975 32.515 37.145 ;
      RECT 32.345 39.695 32.515 39.865 ;
      RECT 32.345 42.415 32.515 42.585 ;
      RECT 32.345 45.135 32.515 45.305 ;
      RECT 32.345 47.855 32.515 48.025 ;
      RECT 32.345 50.575 32.515 50.745 ;
      RECT 32.345 53.295 32.515 53.465 ;
      RECT 32.345 56.015 32.515 56.185 ;
      RECT 32.345 58.735 32.515 58.905 ;
      RECT 31.885 9.775 32.055 9.945 ;
      RECT 31.885 12.495 32.055 12.665 ;
      RECT 31.885 15.215 32.055 15.385 ;
      RECT 31.885 17.935 32.055 18.105 ;
      RECT 31.885 20.655 32.055 20.825 ;
      RECT 31.885 23.375 32.055 23.545 ;
      RECT 31.885 26.095 32.055 26.265 ;
      RECT 31.885 28.815 32.055 28.985 ;
      RECT 31.885 31.535 32.055 31.705 ;
      RECT 31.885 34.255 32.055 34.425 ;
      RECT 31.885 36.975 32.055 37.145 ;
      RECT 31.885 39.695 32.055 39.865 ;
      RECT 31.885 42.415 32.055 42.585 ;
      RECT 31.885 45.135 32.055 45.305 ;
      RECT 31.885 47.855 32.055 48.025 ;
      RECT 31.885 50.575 32.055 50.745 ;
      RECT 31.885 53.295 32.055 53.465 ;
      RECT 31.885 56.015 32.055 56.185 ;
      RECT 31.885 58.735 32.055 58.905 ;
      RECT 31.425 9.775 31.595 9.945 ;
      RECT 31.425 12.495 31.595 12.665 ;
      RECT 31.425 15.215 31.595 15.385 ;
      RECT 31.425 17.935 31.595 18.105 ;
      RECT 31.425 20.655 31.595 20.825 ;
      RECT 31.425 23.375 31.595 23.545 ;
      RECT 31.425 26.095 31.595 26.265 ;
      RECT 31.425 28.815 31.595 28.985 ;
      RECT 31.425 31.535 31.595 31.705 ;
      RECT 31.425 34.255 31.595 34.425 ;
      RECT 31.425 36.975 31.595 37.145 ;
      RECT 31.425 39.695 31.595 39.865 ;
      RECT 31.425 42.415 31.595 42.585 ;
      RECT 31.425 45.135 31.595 45.305 ;
      RECT 31.425 47.855 31.595 48.025 ;
      RECT 31.425 50.575 31.595 50.745 ;
      RECT 31.425 53.295 31.595 53.465 ;
      RECT 31.425 56.015 31.595 56.185 ;
      RECT 31.425 58.735 31.595 58.905 ;
      RECT 30.965 9.775 31.135 9.945 ;
      RECT 30.965 12.495 31.135 12.665 ;
      RECT 30.965 15.215 31.135 15.385 ;
      RECT 30.965 17.935 31.135 18.105 ;
      RECT 30.965 20.655 31.135 20.825 ;
      RECT 30.965 23.375 31.135 23.545 ;
      RECT 30.965 26.095 31.135 26.265 ;
      RECT 30.965 28.815 31.135 28.985 ;
      RECT 30.965 31.535 31.135 31.705 ;
      RECT 30.965 34.255 31.135 34.425 ;
      RECT 30.965 36.975 31.135 37.145 ;
      RECT 30.965 39.695 31.135 39.865 ;
      RECT 30.965 42.415 31.135 42.585 ;
      RECT 30.965 45.135 31.135 45.305 ;
      RECT 30.965 47.855 31.135 48.025 ;
      RECT 30.965 50.575 31.135 50.745 ;
      RECT 30.965 53.295 31.135 53.465 ;
      RECT 30.965 56.015 31.135 56.185 ;
      RECT 30.965 58.735 31.135 58.905 ;
      RECT 30.505 9.775 30.675 9.945 ;
      RECT 30.505 12.495 30.675 12.665 ;
      RECT 30.505 15.215 30.675 15.385 ;
      RECT 30.505 17.935 30.675 18.105 ;
      RECT 30.505 20.655 30.675 20.825 ;
      RECT 30.505 23.375 30.675 23.545 ;
      RECT 30.505 26.095 30.675 26.265 ;
      RECT 30.505 28.815 30.675 28.985 ;
      RECT 30.505 31.535 30.675 31.705 ;
      RECT 30.505 34.255 30.675 34.425 ;
      RECT 30.505 36.975 30.675 37.145 ;
      RECT 30.505 39.695 30.675 39.865 ;
      RECT 30.505 42.415 30.675 42.585 ;
      RECT 30.505 45.135 30.675 45.305 ;
      RECT 30.505 47.855 30.675 48.025 ;
      RECT 30.505 50.575 30.675 50.745 ;
      RECT 30.505 53.295 30.675 53.465 ;
      RECT 30.505 56.015 30.675 56.185 ;
      RECT 30.505 58.735 30.675 58.905 ;
      RECT 30.045 9.775 30.215 9.945 ;
      RECT 30.045 12.495 30.215 12.665 ;
      RECT 30.045 15.215 30.215 15.385 ;
      RECT 30.045 17.935 30.215 18.105 ;
      RECT 30.045 20.655 30.215 20.825 ;
      RECT 30.045 23.375 30.215 23.545 ;
      RECT 30.045 26.095 30.215 26.265 ;
      RECT 30.045 28.815 30.215 28.985 ;
      RECT 30.045 31.535 30.215 31.705 ;
      RECT 30.045 34.255 30.215 34.425 ;
      RECT 30.045 36.975 30.215 37.145 ;
      RECT 30.045 39.695 30.215 39.865 ;
      RECT 30.045 42.415 30.215 42.585 ;
      RECT 30.045 45.135 30.215 45.305 ;
      RECT 30.045 47.855 30.215 48.025 ;
      RECT 30.045 50.575 30.215 50.745 ;
      RECT 30.045 53.295 30.215 53.465 ;
      RECT 30.045 56.015 30.215 56.185 ;
      RECT 30.045 58.735 30.215 58.905 ;
      RECT 29.585 9.775 29.755 9.945 ;
      RECT 29.585 12.495 29.755 12.665 ;
      RECT 29.585 15.215 29.755 15.385 ;
      RECT 29.585 17.935 29.755 18.105 ;
      RECT 29.585 20.655 29.755 20.825 ;
      RECT 29.585 23.375 29.755 23.545 ;
      RECT 29.585 26.095 29.755 26.265 ;
      RECT 29.585 28.815 29.755 28.985 ;
      RECT 29.585 31.535 29.755 31.705 ;
      RECT 29.585 34.255 29.755 34.425 ;
      RECT 29.585 36.975 29.755 37.145 ;
      RECT 29.585 39.695 29.755 39.865 ;
      RECT 29.585 42.415 29.755 42.585 ;
      RECT 29.585 45.135 29.755 45.305 ;
      RECT 29.585 47.855 29.755 48.025 ;
      RECT 29.585 50.575 29.755 50.745 ;
      RECT 29.585 53.295 29.755 53.465 ;
      RECT 29.585 56.015 29.755 56.185 ;
      RECT 29.585 58.735 29.755 58.905 ;
      RECT 29.125 9.775 29.295 9.945 ;
      RECT 29.125 12.495 29.295 12.665 ;
      RECT 29.125 15.215 29.295 15.385 ;
      RECT 29.125 17.935 29.295 18.105 ;
      RECT 29.125 20.655 29.295 20.825 ;
      RECT 29.125 23.375 29.295 23.545 ;
      RECT 29.125 26.095 29.295 26.265 ;
      RECT 29.125 26.605 29.295 26.775 ;
      RECT 29.125 28.815 29.295 28.985 ;
      RECT 29.125 31.535 29.295 31.705 ;
      RECT 29.125 34.255 29.295 34.425 ;
      RECT 29.125 36.975 29.295 37.145 ;
      RECT 29.125 39.695 29.295 39.865 ;
      RECT 29.125 42.415 29.295 42.585 ;
      RECT 29.125 45.135 29.295 45.305 ;
      RECT 29.125 47.855 29.295 48.025 ;
      RECT 29.125 50.575 29.295 50.745 ;
      RECT 29.125 53.295 29.295 53.465 ;
      RECT 29.125 56.015 29.295 56.185 ;
      RECT 29.125 58.735 29.295 58.905 ;
      RECT 28.665 9.775 28.835 9.945 ;
      RECT 28.665 12.495 28.835 12.665 ;
      RECT 28.665 15.215 28.835 15.385 ;
      RECT 28.665 17.935 28.835 18.105 ;
      RECT 28.665 20.655 28.835 20.825 ;
      RECT 28.665 23.375 28.835 23.545 ;
      RECT 28.665 26.095 28.835 26.265 ;
      RECT 28.665 28.815 28.835 28.985 ;
      RECT 28.665 31.535 28.835 31.705 ;
      RECT 28.665 34.255 28.835 34.425 ;
      RECT 28.665 36.975 28.835 37.145 ;
      RECT 28.665 39.695 28.835 39.865 ;
      RECT 28.665 42.415 28.835 42.585 ;
      RECT 28.665 45.135 28.835 45.305 ;
      RECT 28.665 47.855 28.835 48.025 ;
      RECT 28.665 50.575 28.835 50.745 ;
      RECT 28.665 53.295 28.835 53.465 ;
      RECT 28.665 56.015 28.835 56.185 ;
      RECT 28.665 58.735 28.835 58.905 ;
      RECT 28.205 9.775 28.375 9.945 ;
      RECT 28.205 12.495 28.375 12.665 ;
      RECT 28.205 15.215 28.375 15.385 ;
      RECT 28.205 17.935 28.375 18.105 ;
      RECT 28.205 20.655 28.375 20.825 ;
      RECT 28.205 23.375 28.375 23.545 ;
      RECT 28.205 26.095 28.375 26.265 ;
      RECT 28.205 28.815 28.375 28.985 ;
      RECT 28.205 31.535 28.375 31.705 ;
      RECT 28.205 34.255 28.375 34.425 ;
      RECT 28.205 36.975 28.375 37.145 ;
      RECT 28.205 39.695 28.375 39.865 ;
      RECT 28.205 42.415 28.375 42.585 ;
      RECT 28.205 45.135 28.375 45.305 ;
      RECT 28.205 47.855 28.375 48.025 ;
      RECT 28.205 50.575 28.375 50.745 ;
      RECT 28.205 53.295 28.375 53.465 ;
      RECT 28.205 56.015 28.375 56.185 ;
      RECT 28.205 58.735 28.375 58.905 ;
      RECT 27.745 9.775 27.915 9.945 ;
      RECT 27.745 12.495 27.915 12.665 ;
      RECT 27.745 15.215 27.915 15.385 ;
      RECT 27.745 17.935 27.915 18.105 ;
      RECT 27.745 20.655 27.915 20.825 ;
      RECT 27.745 23.375 27.915 23.545 ;
      RECT 27.745 26.095 27.915 26.265 ;
      RECT 27.745 28.815 27.915 28.985 ;
      RECT 27.745 31.535 27.915 31.705 ;
      RECT 27.745 34.255 27.915 34.425 ;
      RECT 27.745 36.975 27.915 37.145 ;
      RECT 27.745 39.695 27.915 39.865 ;
      RECT 27.745 42.415 27.915 42.585 ;
      RECT 27.745 45.135 27.915 45.305 ;
      RECT 27.745 47.855 27.915 48.025 ;
      RECT 27.745 50.575 27.915 50.745 ;
      RECT 27.745 53.295 27.915 53.465 ;
      RECT 27.745 56.015 27.915 56.185 ;
      RECT 27.745 58.735 27.915 58.905 ;
      RECT 27.285 9.775 27.455 9.945 ;
      RECT 27.285 12.495 27.455 12.665 ;
      RECT 27.285 15.215 27.455 15.385 ;
      RECT 27.285 17.935 27.455 18.105 ;
      RECT 27.285 20.655 27.455 20.825 ;
      RECT 27.285 23.375 27.455 23.545 ;
      RECT 27.285 26.095 27.455 26.265 ;
      RECT 27.285 28.815 27.455 28.985 ;
      RECT 27.285 31.535 27.455 31.705 ;
      RECT 27.285 34.255 27.455 34.425 ;
      RECT 27.285 36.975 27.455 37.145 ;
      RECT 27.285 39.695 27.455 39.865 ;
      RECT 27.285 42.415 27.455 42.585 ;
      RECT 27.285 45.135 27.455 45.305 ;
      RECT 27.285 47.855 27.455 48.025 ;
      RECT 27.285 50.575 27.455 50.745 ;
      RECT 27.285 53.295 27.455 53.465 ;
      RECT 27.285 56.015 27.455 56.185 ;
      RECT 27.285 58.735 27.455 58.905 ;
      RECT 26.825 9.775 26.995 9.945 ;
      RECT 26.825 12.495 26.995 12.665 ;
      RECT 26.825 15.215 26.995 15.385 ;
      RECT 26.825 17.935 26.995 18.105 ;
      RECT 26.825 20.655 26.995 20.825 ;
      RECT 26.825 23.375 26.995 23.545 ;
      RECT 26.825 26.095 26.995 26.265 ;
      RECT 26.825 28.815 26.995 28.985 ;
      RECT 26.825 31.535 26.995 31.705 ;
      RECT 26.825 34.255 26.995 34.425 ;
      RECT 26.825 36.975 26.995 37.145 ;
      RECT 26.825 39.695 26.995 39.865 ;
      RECT 26.825 42.415 26.995 42.585 ;
      RECT 26.825 45.135 26.995 45.305 ;
      RECT 26.825 47.855 26.995 48.025 ;
      RECT 26.825 50.575 26.995 50.745 ;
      RECT 26.825 53.295 26.995 53.465 ;
      RECT 26.825 56.015 26.995 56.185 ;
      RECT 26.825 58.735 26.995 58.905 ;
      RECT 26.815 27.285 26.985 27.455 ;
      RECT 26.38 26.945 26.55 27.115 ;
      RECT 26.365 9.775 26.535 9.945 ;
      RECT 26.365 12.495 26.535 12.665 ;
      RECT 26.365 15.215 26.535 15.385 ;
      RECT 26.365 17.935 26.535 18.105 ;
      RECT 26.365 20.655 26.535 20.825 ;
      RECT 26.365 23.375 26.535 23.545 ;
      RECT 26.365 26.095 26.535 26.265 ;
      RECT 26.365 28.815 26.535 28.985 ;
      RECT 26.365 31.535 26.535 31.705 ;
      RECT 26.365 34.255 26.535 34.425 ;
      RECT 26.365 36.975 26.535 37.145 ;
      RECT 26.365 39.695 26.535 39.865 ;
      RECT 26.365 42.415 26.535 42.585 ;
      RECT 26.365 45.135 26.535 45.305 ;
      RECT 26.365 47.855 26.535 48.025 ;
      RECT 26.365 50.575 26.535 50.745 ;
      RECT 26.365 53.295 26.535 53.465 ;
      RECT 26.365 56.015 26.535 56.185 ;
      RECT 26.365 58.735 26.535 58.905 ;
      RECT 25.905 9.775 26.075 9.945 ;
      RECT 25.905 12.495 26.075 12.665 ;
      RECT 25.905 15.215 26.075 15.385 ;
      RECT 25.905 17.935 26.075 18.105 ;
      RECT 25.905 20.655 26.075 20.825 ;
      RECT 25.905 23.375 26.075 23.545 ;
      RECT 25.905 26.095 26.075 26.265 ;
      RECT 25.905 28.815 26.075 28.985 ;
      RECT 25.905 31.535 26.075 31.705 ;
      RECT 25.905 34.255 26.075 34.425 ;
      RECT 25.905 36.975 26.075 37.145 ;
      RECT 25.905 39.695 26.075 39.865 ;
      RECT 25.905 42.415 26.075 42.585 ;
      RECT 25.905 45.135 26.075 45.305 ;
      RECT 25.905 47.855 26.075 48.025 ;
      RECT 25.905 50.575 26.075 50.745 ;
      RECT 25.905 53.295 26.075 53.465 ;
      RECT 25.905 56.015 26.075 56.185 ;
      RECT 25.905 58.735 26.075 58.905 ;
      RECT 25.445 9.775 25.615 9.945 ;
      RECT 25.445 12.495 25.615 12.665 ;
      RECT 25.445 15.215 25.615 15.385 ;
      RECT 25.445 17.935 25.615 18.105 ;
      RECT 25.445 20.655 25.615 20.825 ;
      RECT 25.445 23.375 25.615 23.545 ;
      RECT 25.445 26.095 25.615 26.265 ;
      RECT 25.445 28.815 25.615 28.985 ;
      RECT 25.445 31.535 25.615 31.705 ;
      RECT 25.445 34.255 25.615 34.425 ;
      RECT 25.445 36.975 25.615 37.145 ;
      RECT 25.445 39.695 25.615 39.865 ;
      RECT 25.445 42.415 25.615 42.585 ;
      RECT 25.445 45.135 25.615 45.305 ;
      RECT 25.445 47.855 25.615 48.025 ;
      RECT 25.445 50.575 25.615 50.745 ;
      RECT 25.445 53.295 25.615 53.465 ;
      RECT 25.445 56.015 25.615 56.185 ;
      RECT 25.445 58.735 25.615 58.905 ;
      RECT 24.985 9.775 25.155 9.945 ;
      RECT 24.985 11.305 25.155 11.475 ;
      RECT 24.985 12.495 25.155 12.665 ;
      RECT 24.985 15.215 25.155 15.385 ;
      RECT 24.985 17.935 25.155 18.105 ;
      RECT 24.985 20.655 25.155 20.825 ;
      RECT 24.985 23.375 25.155 23.545 ;
      RECT 24.985 26.095 25.155 26.265 ;
      RECT 24.985 28.815 25.155 28.985 ;
      RECT 24.985 31.535 25.155 31.705 ;
      RECT 24.985 34.255 25.155 34.425 ;
      RECT 24.985 36.975 25.155 37.145 ;
      RECT 24.985 39.695 25.155 39.865 ;
      RECT 24.985 42.415 25.155 42.585 ;
      RECT 24.985 45.135 25.155 45.305 ;
      RECT 24.985 47.855 25.155 48.025 ;
      RECT 24.985 50.575 25.155 50.745 ;
      RECT 24.985 53.295 25.155 53.465 ;
      RECT 24.985 56.015 25.155 56.185 ;
      RECT 24.985 58.735 25.155 58.905 ;
      RECT 24.81 26.945 24.98 27.115 ;
      RECT 24.525 9.775 24.695 9.945 ;
      RECT 24.525 12.495 24.695 12.665 ;
      RECT 24.525 15.215 24.695 15.385 ;
      RECT 24.525 17.935 24.695 18.105 ;
      RECT 24.525 20.655 24.695 20.825 ;
      RECT 24.525 23.375 24.695 23.545 ;
      RECT 24.525 26.095 24.695 26.265 ;
      RECT 24.525 28.815 24.695 28.985 ;
      RECT 24.525 31.535 24.695 31.705 ;
      RECT 24.525 34.255 24.695 34.425 ;
      RECT 24.525 36.975 24.695 37.145 ;
      RECT 24.525 39.695 24.695 39.865 ;
      RECT 24.525 42.415 24.695 42.585 ;
      RECT 24.525 45.135 24.695 45.305 ;
      RECT 24.525 47.855 24.695 48.025 ;
      RECT 24.525 50.575 24.695 50.745 ;
      RECT 24.525 53.295 24.695 53.465 ;
      RECT 24.525 56.015 24.695 56.185 ;
      RECT 24.525 58.735 24.695 58.905 ;
      RECT 24.295 27.285 24.465 27.455 ;
      RECT 24.065 9.775 24.235 9.945 ;
      RECT 24.065 12.495 24.235 12.665 ;
      RECT 24.065 15.215 24.235 15.385 ;
      RECT 24.065 17.935 24.235 18.105 ;
      RECT 24.065 20.655 24.235 20.825 ;
      RECT 24.065 23.375 24.235 23.545 ;
      RECT 24.065 26.095 24.235 26.265 ;
      RECT 24.065 28.815 24.235 28.985 ;
      RECT 24.065 31.535 24.235 31.705 ;
      RECT 24.065 34.255 24.235 34.425 ;
      RECT 24.065 36.975 24.235 37.145 ;
      RECT 24.065 39.695 24.235 39.865 ;
      RECT 24.065 42.415 24.235 42.585 ;
      RECT 24.065 45.135 24.235 45.305 ;
      RECT 24.065 47.855 24.235 48.025 ;
      RECT 24.065 50.575 24.235 50.745 ;
      RECT 24.065 53.295 24.235 53.465 ;
      RECT 24.065 56.015 24.235 56.185 ;
      RECT 24.065 58.735 24.235 58.905 ;
      RECT 23.605 9.775 23.775 9.945 ;
      RECT 23.605 12.495 23.775 12.665 ;
      RECT 23.605 15.215 23.775 15.385 ;
      RECT 23.605 17.935 23.775 18.105 ;
      RECT 23.605 20.655 23.775 20.825 ;
      RECT 23.605 23.375 23.775 23.545 ;
      RECT 23.605 26.095 23.775 26.265 ;
      RECT 23.605 28.815 23.775 28.985 ;
      RECT 23.605 31.535 23.775 31.705 ;
      RECT 23.605 34.255 23.775 34.425 ;
      RECT 23.605 36.975 23.775 37.145 ;
      RECT 23.605 39.695 23.775 39.865 ;
      RECT 23.605 42.415 23.775 42.585 ;
      RECT 23.605 45.135 23.775 45.305 ;
      RECT 23.605 47.855 23.775 48.025 ;
      RECT 23.605 50.575 23.775 50.745 ;
      RECT 23.605 53.295 23.775 53.465 ;
      RECT 23.605 56.015 23.775 56.185 ;
      RECT 23.605 58.735 23.775 58.905 ;
      RECT 23.53 27.965 23.7 28.135 ;
      RECT 23.145 9.775 23.315 9.945 ;
      RECT 23.145 12.495 23.315 12.665 ;
      RECT 23.145 15.215 23.315 15.385 ;
      RECT 23.145 17.935 23.315 18.105 ;
      RECT 23.145 20.655 23.315 20.825 ;
      RECT 23.145 23.375 23.315 23.545 ;
      RECT 23.145 26.095 23.315 26.265 ;
      RECT 23.145 28.815 23.315 28.985 ;
      RECT 23.145 31.535 23.315 31.705 ;
      RECT 23.145 34.255 23.315 34.425 ;
      RECT 23.145 36.975 23.315 37.145 ;
      RECT 23.145 39.695 23.315 39.865 ;
      RECT 23.145 42.415 23.315 42.585 ;
      RECT 23.145 45.135 23.315 45.305 ;
      RECT 23.145 47.855 23.315 48.025 ;
      RECT 23.145 50.575 23.315 50.745 ;
      RECT 23.145 53.295 23.315 53.465 ;
      RECT 23.145 56.015 23.315 56.185 ;
      RECT 23.145 58.735 23.315 58.905 ;
      RECT 23.105 27.285 23.275 27.455 ;
      RECT 22.71 26.945 22.88 27.115 ;
      RECT 22.685 9.775 22.855 9.945 ;
      RECT 22.685 12.495 22.855 12.665 ;
      RECT 22.685 15.215 22.855 15.385 ;
      RECT 22.685 17.935 22.855 18.105 ;
      RECT 22.685 20.655 22.855 20.825 ;
      RECT 22.685 23.375 22.855 23.545 ;
      RECT 22.685 26.095 22.855 26.265 ;
      RECT 22.685 28.815 22.855 28.985 ;
      RECT 22.685 31.535 22.855 31.705 ;
      RECT 22.685 34.255 22.855 34.425 ;
      RECT 22.685 36.975 22.855 37.145 ;
      RECT 22.685 39.695 22.855 39.865 ;
      RECT 22.685 42.415 22.855 42.585 ;
      RECT 22.685 45.135 22.855 45.305 ;
      RECT 22.685 47.855 22.855 48.025 ;
      RECT 22.685 50.575 22.855 50.745 ;
      RECT 22.685 53.295 22.855 53.465 ;
      RECT 22.685 56.015 22.855 56.185 ;
      RECT 22.685 58.735 22.855 58.905 ;
      RECT 22.225 9.775 22.395 9.945 ;
      RECT 22.225 12.495 22.395 12.665 ;
      RECT 22.225 15.215 22.395 15.385 ;
      RECT 22.225 17.935 22.395 18.105 ;
      RECT 22.225 20.655 22.395 20.825 ;
      RECT 22.225 23.375 22.395 23.545 ;
      RECT 22.225 26.095 22.395 26.265 ;
      RECT 22.225 27.625 22.395 27.795 ;
      RECT 22.225 28.815 22.395 28.985 ;
      RECT 22.225 31.535 22.395 31.705 ;
      RECT 22.225 34.255 22.395 34.425 ;
      RECT 22.225 36.975 22.395 37.145 ;
      RECT 22.225 39.695 22.395 39.865 ;
      RECT 22.225 42.415 22.395 42.585 ;
      RECT 22.225 45.135 22.395 45.305 ;
      RECT 22.225 47.855 22.395 48.025 ;
      RECT 22.225 50.575 22.395 50.745 ;
      RECT 22.225 53.295 22.395 53.465 ;
      RECT 22.225 56.015 22.395 56.185 ;
      RECT 22.225 58.735 22.395 58.905 ;
      RECT 21.765 9.775 21.935 9.945 ;
      RECT 21.765 12.495 21.935 12.665 ;
      RECT 21.765 15.215 21.935 15.385 ;
      RECT 21.765 17.935 21.935 18.105 ;
      RECT 21.765 20.655 21.935 20.825 ;
      RECT 21.765 23.375 21.935 23.545 ;
      RECT 21.765 26.095 21.935 26.265 ;
      RECT 21.765 28.815 21.935 28.985 ;
      RECT 21.765 31.535 21.935 31.705 ;
      RECT 21.765 34.255 21.935 34.425 ;
      RECT 21.765 36.975 21.935 37.145 ;
      RECT 21.765 39.695 21.935 39.865 ;
      RECT 21.765 42.415 21.935 42.585 ;
      RECT 21.765 45.135 21.935 45.305 ;
      RECT 21.765 47.855 21.935 48.025 ;
      RECT 21.765 50.575 21.935 50.745 ;
      RECT 21.765 53.295 21.935 53.465 ;
      RECT 21.765 56.015 21.935 56.185 ;
      RECT 21.765 58.735 21.935 58.905 ;
      RECT 21.305 9.775 21.475 9.945 ;
      RECT 21.305 12.495 21.475 12.665 ;
      RECT 21.305 15.215 21.475 15.385 ;
      RECT 21.305 17.935 21.475 18.105 ;
      RECT 21.305 19.125 21.475 19.295 ;
      RECT 21.305 20.655 21.475 20.825 ;
      RECT 21.305 23.375 21.475 23.545 ;
      RECT 21.305 26.095 21.475 26.265 ;
      RECT 21.305 28.815 21.475 28.985 ;
      RECT 21.305 31.535 21.475 31.705 ;
      RECT 21.305 34.255 21.475 34.425 ;
      RECT 21.305 36.975 21.475 37.145 ;
      RECT 21.305 39.695 21.475 39.865 ;
      RECT 21.305 42.415 21.475 42.585 ;
      RECT 21.305 45.135 21.475 45.305 ;
      RECT 21.305 47.855 21.475 48.025 ;
      RECT 21.305 50.575 21.475 50.745 ;
      RECT 21.305 53.295 21.475 53.465 ;
      RECT 21.305 56.015 21.475 56.185 ;
      RECT 21.305 58.735 21.475 58.905 ;
      RECT 20.845 9.775 21.015 9.945 ;
      RECT 20.845 12.495 21.015 12.665 ;
      RECT 20.845 15.215 21.015 15.385 ;
      RECT 20.845 17.935 21.015 18.105 ;
      RECT 20.845 20.655 21.015 20.825 ;
      RECT 20.845 23.375 21.015 23.545 ;
      RECT 20.845 26.095 21.015 26.265 ;
      RECT 20.845 28.815 21.015 28.985 ;
      RECT 20.845 31.535 21.015 31.705 ;
      RECT 20.845 34.255 21.015 34.425 ;
      RECT 20.845 36.975 21.015 37.145 ;
      RECT 20.845 39.695 21.015 39.865 ;
      RECT 20.845 42.415 21.015 42.585 ;
      RECT 20.845 45.135 21.015 45.305 ;
      RECT 20.845 47.855 21.015 48.025 ;
      RECT 20.845 50.575 21.015 50.745 ;
      RECT 20.845 53.295 21.015 53.465 ;
      RECT 20.845 56.015 21.015 56.185 ;
      RECT 20.845 58.735 21.015 58.905 ;
      RECT 20.385 9.775 20.555 9.945 ;
      RECT 20.385 12.495 20.555 12.665 ;
      RECT 20.385 15.215 20.555 15.385 ;
      RECT 20.385 17.935 20.555 18.105 ;
      RECT 20.385 20.655 20.555 20.825 ;
      RECT 20.385 23.375 20.555 23.545 ;
      RECT 20.385 26.095 20.555 26.265 ;
      RECT 20.385 28.815 20.555 28.985 ;
      RECT 20.385 31.535 20.555 31.705 ;
      RECT 20.385 34.255 20.555 34.425 ;
      RECT 20.385 36.975 20.555 37.145 ;
      RECT 20.385 39.695 20.555 39.865 ;
      RECT 20.385 42.415 20.555 42.585 ;
      RECT 20.385 45.135 20.555 45.305 ;
      RECT 20.385 47.855 20.555 48.025 ;
      RECT 20.385 50.575 20.555 50.745 ;
      RECT 20.385 53.295 20.555 53.465 ;
      RECT 20.385 56.015 20.555 56.185 ;
      RECT 20.385 58.735 20.555 58.905 ;
      RECT 19.925 9.775 20.095 9.945 ;
      RECT 19.925 12.495 20.095 12.665 ;
      RECT 19.925 15.215 20.095 15.385 ;
      RECT 19.925 17.935 20.095 18.105 ;
      RECT 19.925 20.655 20.095 20.825 ;
      RECT 19.925 23.375 20.095 23.545 ;
      RECT 19.925 26.095 20.095 26.265 ;
      RECT 19.925 28.815 20.095 28.985 ;
      RECT 19.925 31.535 20.095 31.705 ;
      RECT 19.925 34.255 20.095 34.425 ;
      RECT 19.925 36.975 20.095 37.145 ;
      RECT 19.925 39.695 20.095 39.865 ;
      RECT 19.925 42.415 20.095 42.585 ;
      RECT 19.925 45.135 20.095 45.305 ;
      RECT 19.925 47.855 20.095 48.025 ;
      RECT 19.925 50.575 20.095 50.745 ;
      RECT 19.925 53.295 20.095 53.465 ;
      RECT 19.925 56.015 20.095 56.185 ;
      RECT 19.925 58.735 20.095 58.905 ;
      RECT 19.465 9.775 19.635 9.945 ;
      RECT 19.465 12.495 19.635 12.665 ;
      RECT 19.465 15.215 19.635 15.385 ;
      RECT 19.465 17.935 19.635 18.105 ;
      RECT 19.465 20.655 19.635 20.825 ;
      RECT 19.465 23.375 19.635 23.545 ;
      RECT 19.465 26.095 19.635 26.265 ;
      RECT 19.465 28.815 19.635 28.985 ;
      RECT 19.465 31.535 19.635 31.705 ;
      RECT 19.465 34.255 19.635 34.425 ;
      RECT 19.465 36.975 19.635 37.145 ;
      RECT 19.465 39.695 19.635 39.865 ;
      RECT 19.465 42.415 19.635 42.585 ;
      RECT 19.465 45.135 19.635 45.305 ;
      RECT 19.465 47.855 19.635 48.025 ;
      RECT 19.465 50.575 19.635 50.745 ;
      RECT 19.465 53.295 19.635 53.465 ;
      RECT 19.465 56.015 19.635 56.185 ;
      RECT 19.465 58.735 19.635 58.905 ;
      RECT 19.005 9.775 19.175 9.945 ;
      RECT 19.005 12.495 19.175 12.665 ;
      RECT 19.005 15.215 19.175 15.385 ;
      RECT 19.005 17.935 19.175 18.105 ;
      RECT 19.005 20.655 19.175 20.825 ;
      RECT 19.005 23.375 19.175 23.545 ;
      RECT 19.005 26.095 19.175 26.265 ;
      RECT 19.005 28.815 19.175 28.985 ;
      RECT 19.005 31.535 19.175 31.705 ;
      RECT 19.005 34.255 19.175 34.425 ;
      RECT 19.005 36.975 19.175 37.145 ;
      RECT 19.005 39.695 19.175 39.865 ;
      RECT 19.005 42.415 19.175 42.585 ;
      RECT 19.005 45.135 19.175 45.305 ;
      RECT 19.005 47.855 19.175 48.025 ;
      RECT 19.005 50.575 19.175 50.745 ;
      RECT 19.005 53.295 19.175 53.465 ;
      RECT 19.005 56.015 19.175 56.185 ;
      RECT 19.005 58.735 19.175 58.905 ;
      RECT 18.545 9.775 18.715 9.945 ;
      RECT 18.545 12.495 18.715 12.665 ;
      RECT 18.545 15.215 18.715 15.385 ;
      RECT 18.545 17.935 18.715 18.105 ;
      RECT 18.545 20.655 18.715 20.825 ;
      RECT 18.545 22.185 18.715 22.355 ;
      RECT 18.545 23.375 18.715 23.545 ;
      RECT 18.545 26.095 18.715 26.265 ;
      RECT 18.545 28.815 18.715 28.985 ;
      RECT 18.545 31.535 18.715 31.705 ;
      RECT 18.545 34.255 18.715 34.425 ;
      RECT 18.545 36.975 18.715 37.145 ;
      RECT 18.545 39.695 18.715 39.865 ;
      RECT 18.545 42.415 18.715 42.585 ;
      RECT 18.545 45.135 18.715 45.305 ;
      RECT 18.545 47.855 18.715 48.025 ;
      RECT 18.545 50.575 18.715 50.745 ;
      RECT 18.545 53.295 18.715 53.465 ;
      RECT 18.545 56.015 18.715 56.185 ;
      RECT 18.545 58.735 18.715 58.905 ;
      RECT 18.085 9.775 18.255 9.945 ;
      RECT 18.085 12.495 18.255 12.665 ;
      RECT 18.085 15.215 18.255 15.385 ;
      RECT 18.085 17.935 18.255 18.105 ;
      RECT 18.085 20.655 18.255 20.825 ;
      RECT 18.085 23.375 18.255 23.545 ;
      RECT 18.085 26.095 18.255 26.265 ;
      RECT 18.085 28.815 18.255 28.985 ;
      RECT 18.085 31.535 18.255 31.705 ;
      RECT 18.085 34.255 18.255 34.425 ;
      RECT 18.085 36.975 18.255 37.145 ;
      RECT 18.085 39.695 18.255 39.865 ;
      RECT 18.085 42.415 18.255 42.585 ;
      RECT 18.085 45.135 18.255 45.305 ;
      RECT 18.085 47.855 18.255 48.025 ;
      RECT 18.085 50.575 18.255 50.745 ;
      RECT 18.085 53.295 18.255 53.465 ;
      RECT 18.085 56.015 18.255 56.185 ;
      RECT 18.085 58.735 18.255 58.905 ;
      RECT 17.625 9.775 17.795 9.945 ;
      RECT 17.625 12.495 17.795 12.665 ;
      RECT 17.625 15.215 17.795 15.385 ;
      RECT 17.625 17.935 17.795 18.105 ;
      RECT 17.625 20.655 17.795 20.825 ;
      RECT 17.625 23.375 17.795 23.545 ;
      RECT 17.625 26.095 17.795 26.265 ;
      RECT 17.625 28.815 17.795 28.985 ;
      RECT 17.625 31.535 17.795 31.705 ;
      RECT 17.625 34.255 17.795 34.425 ;
      RECT 17.625 36.975 17.795 37.145 ;
      RECT 17.625 39.695 17.795 39.865 ;
      RECT 17.625 42.415 17.795 42.585 ;
      RECT 17.625 45.135 17.795 45.305 ;
      RECT 17.625 47.855 17.795 48.025 ;
      RECT 17.625 50.575 17.795 50.745 ;
      RECT 17.625 53.295 17.795 53.465 ;
      RECT 17.625 56.015 17.795 56.185 ;
      RECT 17.625 58.735 17.795 58.905 ;
      RECT 17.165 9.775 17.335 9.945 ;
      RECT 17.165 12.495 17.335 12.665 ;
      RECT 17.165 15.215 17.335 15.385 ;
      RECT 17.165 17.935 17.335 18.105 ;
      RECT 17.165 20.655 17.335 20.825 ;
      RECT 17.165 23.375 17.335 23.545 ;
      RECT 17.165 26.095 17.335 26.265 ;
      RECT 17.165 28.815 17.335 28.985 ;
      RECT 17.165 31.535 17.335 31.705 ;
      RECT 17.165 34.255 17.335 34.425 ;
      RECT 17.165 36.975 17.335 37.145 ;
      RECT 17.165 39.695 17.335 39.865 ;
      RECT 17.165 42.415 17.335 42.585 ;
      RECT 17.165 45.135 17.335 45.305 ;
      RECT 17.165 47.855 17.335 48.025 ;
      RECT 17.165 50.575 17.335 50.745 ;
      RECT 17.165 53.295 17.335 53.465 ;
      RECT 17.165 56.015 17.335 56.185 ;
      RECT 17.165 58.735 17.335 58.905 ;
      RECT 16.705 9.775 16.875 9.945 ;
      RECT 16.705 11.305 16.875 11.475 ;
      RECT 16.705 12.495 16.875 12.665 ;
      RECT 16.705 15.215 16.875 15.385 ;
      RECT 16.705 17.935 16.875 18.105 ;
      RECT 16.705 20.655 16.875 20.825 ;
      RECT 16.705 23.375 16.875 23.545 ;
      RECT 16.705 26.095 16.875 26.265 ;
      RECT 16.705 28.815 16.875 28.985 ;
      RECT 16.705 31.535 16.875 31.705 ;
      RECT 16.705 34.255 16.875 34.425 ;
      RECT 16.705 36.975 16.875 37.145 ;
      RECT 16.705 39.695 16.875 39.865 ;
      RECT 16.705 42.415 16.875 42.585 ;
      RECT 16.705 45.135 16.875 45.305 ;
      RECT 16.705 47.855 16.875 48.025 ;
      RECT 16.705 50.575 16.875 50.745 ;
      RECT 16.705 53.295 16.875 53.465 ;
      RECT 16.705 56.015 16.875 56.185 ;
      RECT 16.705 58.735 16.875 58.905 ;
      RECT 16.245 9.775 16.415 9.945 ;
      RECT 16.245 12.495 16.415 12.665 ;
      RECT 16.245 15.215 16.415 15.385 ;
      RECT 16.245 17.935 16.415 18.105 ;
      RECT 16.245 20.655 16.415 20.825 ;
      RECT 16.245 23.375 16.415 23.545 ;
      RECT 16.245 26.095 16.415 26.265 ;
      RECT 16.245 28.815 16.415 28.985 ;
      RECT 16.245 31.535 16.415 31.705 ;
      RECT 16.245 34.255 16.415 34.425 ;
      RECT 16.245 36.975 16.415 37.145 ;
      RECT 16.245 39.695 16.415 39.865 ;
      RECT 16.245 42.415 16.415 42.585 ;
      RECT 16.245 45.135 16.415 45.305 ;
      RECT 16.245 47.855 16.415 48.025 ;
      RECT 16.245 50.575 16.415 50.745 ;
      RECT 16.245 53.295 16.415 53.465 ;
      RECT 16.245 56.015 16.415 56.185 ;
      RECT 16.245 58.735 16.415 58.905 ;
      RECT 15.785 9.775 15.955 9.945 ;
      RECT 15.785 12.495 15.955 12.665 ;
      RECT 15.785 15.215 15.955 15.385 ;
      RECT 15.785 17.935 15.955 18.105 ;
      RECT 15.785 20.655 15.955 20.825 ;
      RECT 15.785 23.375 15.955 23.545 ;
      RECT 15.785 26.095 15.955 26.265 ;
      RECT 15.785 28.815 15.955 28.985 ;
      RECT 15.785 31.535 15.955 31.705 ;
      RECT 15.785 34.255 15.955 34.425 ;
      RECT 15.785 36.975 15.955 37.145 ;
      RECT 15.785 39.695 15.955 39.865 ;
      RECT 15.785 42.415 15.955 42.585 ;
      RECT 15.785 45.135 15.955 45.305 ;
      RECT 15.785 47.855 15.955 48.025 ;
      RECT 15.785 50.575 15.955 50.745 ;
      RECT 15.785 53.295 15.955 53.465 ;
      RECT 15.785 56.015 15.955 56.185 ;
      RECT 15.785 58.735 15.955 58.905 ;
      RECT 15.325 9.775 15.495 9.945 ;
      RECT 15.325 12.495 15.495 12.665 ;
      RECT 15.325 15.215 15.495 15.385 ;
      RECT 15.325 17.935 15.495 18.105 ;
      RECT 15.325 20.655 15.495 20.825 ;
      RECT 15.325 23.375 15.495 23.545 ;
      RECT 15.325 26.095 15.495 26.265 ;
      RECT 15.325 28.815 15.495 28.985 ;
      RECT 15.325 31.535 15.495 31.705 ;
      RECT 15.325 34.255 15.495 34.425 ;
      RECT 15.325 36.975 15.495 37.145 ;
      RECT 15.325 39.695 15.495 39.865 ;
      RECT 15.325 42.415 15.495 42.585 ;
      RECT 15.325 45.135 15.495 45.305 ;
      RECT 15.325 47.855 15.495 48.025 ;
      RECT 15.325 50.575 15.495 50.745 ;
      RECT 15.325 53.295 15.495 53.465 ;
      RECT 15.325 56.015 15.495 56.185 ;
      RECT 15.325 58.735 15.495 58.905 ;
      RECT 14.865 9.775 15.035 9.945 ;
      RECT 14.865 12.495 15.035 12.665 ;
      RECT 14.865 15.215 15.035 15.385 ;
      RECT 14.865 17.935 15.035 18.105 ;
      RECT 14.865 20.655 15.035 20.825 ;
      RECT 14.865 23.375 15.035 23.545 ;
      RECT 14.865 26.095 15.035 26.265 ;
      RECT 14.865 28.815 15.035 28.985 ;
      RECT 14.865 31.535 15.035 31.705 ;
      RECT 14.865 34.255 15.035 34.425 ;
      RECT 14.865 36.975 15.035 37.145 ;
      RECT 14.865 39.695 15.035 39.865 ;
      RECT 14.865 42.415 15.035 42.585 ;
      RECT 14.865 45.135 15.035 45.305 ;
      RECT 14.865 47.855 15.035 48.025 ;
      RECT 14.865 50.575 15.035 50.745 ;
      RECT 14.865 53.295 15.035 53.465 ;
      RECT 14.865 56.015 15.035 56.185 ;
      RECT 14.865 58.735 15.035 58.905 ;
      RECT 14.405 9.775 14.575 9.945 ;
      RECT 14.405 12.495 14.575 12.665 ;
      RECT 14.405 15.215 14.575 15.385 ;
      RECT 14.405 17.935 14.575 18.105 ;
      RECT 14.405 20.655 14.575 20.825 ;
      RECT 14.405 23.375 14.575 23.545 ;
      RECT 14.405 26.095 14.575 26.265 ;
      RECT 14.405 28.815 14.575 28.985 ;
      RECT 14.405 31.535 14.575 31.705 ;
      RECT 14.405 34.255 14.575 34.425 ;
      RECT 14.405 36.975 14.575 37.145 ;
      RECT 14.405 39.695 14.575 39.865 ;
      RECT 14.405 42.415 14.575 42.585 ;
      RECT 14.405 45.135 14.575 45.305 ;
      RECT 14.405 47.855 14.575 48.025 ;
      RECT 14.405 50.575 14.575 50.745 ;
      RECT 14.405 53.295 14.575 53.465 ;
      RECT 14.405 56.015 14.575 56.185 ;
      RECT 14.405 58.735 14.575 58.905 ;
      RECT 13.945 9.775 14.115 9.945 ;
      RECT 13.945 12.495 14.115 12.665 ;
      RECT 13.945 15.215 14.115 15.385 ;
      RECT 13.945 17.935 14.115 18.105 ;
      RECT 13.945 20.655 14.115 20.825 ;
      RECT 13.945 23.375 14.115 23.545 ;
      RECT 13.945 26.095 14.115 26.265 ;
      RECT 13.945 28.815 14.115 28.985 ;
      RECT 13.945 31.535 14.115 31.705 ;
      RECT 13.945 34.255 14.115 34.425 ;
      RECT 13.945 36.975 14.115 37.145 ;
      RECT 13.945 39.695 14.115 39.865 ;
      RECT 13.945 42.415 14.115 42.585 ;
      RECT 13.945 45.135 14.115 45.305 ;
      RECT 13.945 47.855 14.115 48.025 ;
      RECT 13.945 50.575 14.115 50.745 ;
      RECT 13.945 53.295 14.115 53.465 ;
      RECT 13.945 56.015 14.115 56.185 ;
      RECT 13.945 58.735 14.115 58.905 ;
      RECT 13.485 9.775 13.655 9.945 ;
      RECT 13.485 12.495 13.655 12.665 ;
      RECT 13.485 15.215 13.655 15.385 ;
      RECT 13.485 17.935 13.655 18.105 ;
      RECT 13.485 20.655 13.655 20.825 ;
      RECT 13.485 23.375 13.655 23.545 ;
      RECT 13.485 26.095 13.655 26.265 ;
      RECT 13.485 28.815 13.655 28.985 ;
      RECT 13.485 31.535 13.655 31.705 ;
      RECT 13.485 34.255 13.655 34.425 ;
      RECT 13.485 36.975 13.655 37.145 ;
      RECT 13.485 39.695 13.655 39.865 ;
      RECT 13.485 42.415 13.655 42.585 ;
      RECT 13.485 45.135 13.655 45.305 ;
      RECT 13.485 47.855 13.655 48.025 ;
      RECT 13.485 50.575 13.655 50.745 ;
      RECT 13.485 53.295 13.655 53.465 ;
      RECT 13.485 56.015 13.655 56.185 ;
      RECT 13.485 58.735 13.655 58.905 ;
      RECT 13.025 9.775 13.195 9.945 ;
      RECT 13.025 12.495 13.195 12.665 ;
      RECT 13.025 15.215 13.195 15.385 ;
      RECT 13.025 17.935 13.195 18.105 ;
      RECT 13.025 20.655 13.195 20.825 ;
      RECT 13.025 23.375 13.195 23.545 ;
      RECT 13.025 26.095 13.195 26.265 ;
      RECT 13.025 28.815 13.195 28.985 ;
      RECT 13.025 31.535 13.195 31.705 ;
      RECT 13.025 34.255 13.195 34.425 ;
      RECT 13.025 36.975 13.195 37.145 ;
      RECT 13.025 39.695 13.195 39.865 ;
      RECT 13.025 42.415 13.195 42.585 ;
      RECT 13.025 45.135 13.195 45.305 ;
      RECT 13.025 47.855 13.195 48.025 ;
      RECT 13.025 50.575 13.195 50.745 ;
      RECT 13.025 53.295 13.195 53.465 ;
      RECT 13.025 56.015 13.195 56.185 ;
      RECT 13.025 58.735 13.195 58.905 ;
      RECT 12.565 9.775 12.735 9.945 ;
      RECT 12.565 12.495 12.735 12.665 ;
      RECT 12.565 15.215 12.735 15.385 ;
      RECT 12.565 17.935 12.735 18.105 ;
      RECT 12.565 20.655 12.735 20.825 ;
      RECT 12.565 23.375 12.735 23.545 ;
      RECT 12.565 26.095 12.735 26.265 ;
      RECT 12.565 28.815 12.735 28.985 ;
      RECT 12.565 31.535 12.735 31.705 ;
      RECT 12.565 34.255 12.735 34.425 ;
      RECT 12.565 36.975 12.735 37.145 ;
      RECT 12.565 39.695 12.735 39.865 ;
      RECT 12.565 42.415 12.735 42.585 ;
      RECT 12.565 45.135 12.735 45.305 ;
      RECT 12.565 47.855 12.735 48.025 ;
      RECT 12.565 50.575 12.735 50.745 ;
      RECT 12.565 53.295 12.735 53.465 ;
      RECT 12.565 56.015 12.735 56.185 ;
      RECT 12.565 58.735 12.735 58.905 ;
      RECT 12.105 9.775 12.275 9.945 ;
      RECT 12.105 12.495 12.275 12.665 ;
      RECT 12.105 15.215 12.275 15.385 ;
      RECT 12.105 17.935 12.275 18.105 ;
      RECT 12.105 20.655 12.275 20.825 ;
      RECT 12.105 23.375 12.275 23.545 ;
      RECT 12.105 26.095 12.275 26.265 ;
      RECT 12.105 28.815 12.275 28.985 ;
      RECT 12.105 31.535 12.275 31.705 ;
      RECT 12.105 34.255 12.275 34.425 ;
      RECT 12.105 36.975 12.275 37.145 ;
      RECT 12.105 39.695 12.275 39.865 ;
      RECT 12.105 42.415 12.275 42.585 ;
      RECT 12.105 45.135 12.275 45.305 ;
      RECT 12.105 47.855 12.275 48.025 ;
      RECT 12.105 50.575 12.275 50.745 ;
      RECT 12.105 53.295 12.275 53.465 ;
      RECT 12.105 56.015 12.275 56.185 ;
      RECT 12.105 58.735 12.275 58.905 ;
      RECT 11.645 9.775 11.815 9.945 ;
      RECT 11.645 12.495 11.815 12.665 ;
      RECT 11.645 15.215 11.815 15.385 ;
      RECT 11.645 17.935 11.815 18.105 ;
      RECT 11.645 20.655 11.815 20.825 ;
      RECT 11.645 23.375 11.815 23.545 ;
      RECT 11.645 26.095 11.815 26.265 ;
      RECT 11.645 28.815 11.815 28.985 ;
      RECT 11.645 31.535 11.815 31.705 ;
      RECT 11.645 34.255 11.815 34.425 ;
      RECT 11.645 36.975 11.815 37.145 ;
      RECT 11.645 39.695 11.815 39.865 ;
      RECT 11.645 42.415 11.815 42.585 ;
      RECT 11.645 45.135 11.815 45.305 ;
      RECT 11.645 47.855 11.815 48.025 ;
      RECT 11.645 50.575 11.815 50.745 ;
      RECT 11.645 53.295 11.815 53.465 ;
      RECT 11.645 56.015 11.815 56.185 ;
      RECT 11.645 58.735 11.815 58.905 ;
      RECT 11.185 9.775 11.355 9.945 ;
      RECT 11.185 12.495 11.355 12.665 ;
      RECT 11.185 15.215 11.355 15.385 ;
      RECT 11.185 17.935 11.355 18.105 ;
      RECT 11.185 20.655 11.355 20.825 ;
      RECT 11.185 23.375 11.355 23.545 ;
      RECT 11.185 26.095 11.355 26.265 ;
      RECT 11.185 28.815 11.355 28.985 ;
      RECT 11.185 31.535 11.355 31.705 ;
      RECT 11.185 34.255 11.355 34.425 ;
      RECT 11.185 36.975 11.355 37.145 ;
      RECT 11.185 39.695 11.355 39.865 ;
      RECT 11.185 42.415 11.355 42.585 ;
      RECT 11.185 45.135 11.355 45.305 ;
      RECT 11.185 47.855 11.355 48.025 ;
      RECT 11.185 50.575 11.355 50.745 ;
      RECT 11.185 53.295 11.355 53.465 ;
      RECT 11.185 56.015 11.355 56.185 ;
      RECT 11.185 58.735 11.355 58.905 ;
      RECT 10.725 9.775 10.895 9.945 ;
      RECT 10.725 12.495 10.895 12.665 ;
      RECT 10.725 15.215 10.895 15.385 ;
      RECT 10.725 17.935 10.895 18.105 ;
      RECT 10.725 20.655 10.895 20.825 ;
      RECT 10.725 23.375 10.895 23.545 ;
      RECT 10.725 26.095 10.895 26.265 ;
      RECT 10.725 28.815 10.895 28.985 ;
      RECT 10.725 31.535 10.895 31.705 ;
      RECT 10.725 34.255 10.895 34.425 ;
      RECT 10.725 36.975 10.895 37.145 ;
      RECT 10.725 39.695 10.895 39.865 ;
      RECT 10.725 42.415 10.895 42.585 ;
      RECT 10.725 45.135 10.895 45.305 ;
      RECT 10.725 47.855 10.895 48.025 ;
      RECT 10.725 50.575 10.895 50.745 ;
      RECT 10.725 53.295 10.895 53.465 ;
      RECT 10.725 56.015 10.895 56.185 ;
      RECT 10.725 58.735 10.895 58.905 ;
      RECT 10.265 9.775 10.435 9.945 ;
      RECT 10.265 12.495 10.435 12.665 ;
      RECT 10.265 15.215 10.435 15.385 ;
      RECT 10.265 17.935 10.435 18.105 ;
      RECT 10.265 20.655 10.435 20.825 ;
      RECT 10.265 23.375 10.435 23.545 ;
      RECT 10.265 26.095 10.435 26.265 ;
      RECT 10.265 28.815 10.435 28.985 ;
      RECT 10.265 31.535 10.435 31.705 ;
      RECT 10.265 34.255 10.435 34.425 ;
      RECT 10.265 36.975 10.435 37.145 ;
      RECT 10.265 39.695 10.435 39.865 ;
      RECT 10.265 42.415 10.435 42.585 ;
      RECT 10.265 45.135 10.435 45.305 ;
      RECT 10.265 47.855 10.435 48.025 ;
      RECT 10.265 50.575 10.435 50.745 ;
      RECT 10.265 53.295 10.435 53.465 ;
      RECT 10.265 56.015 10.435 56.185 ;
      RECT 10.265 58.735 10.435 58.905 ;
    LAYER met1 ;
      RECT 177.17 15.68 177.49 15.94 ;
      RECT 184.085 15.695 184.375 15.925 ;
      RECT 177.17 15.74 184.375 15.88 ;
      RECT 179.93 11.94 180.25 12.2 ;
      RECT 183.625 11.955 183.915 12.185 ;
      RECT 179.93 12 183.915 12.14 ;
      RECT 181.775 16.375 182.065 16.605 ;
      RECT 179.255 16.375 179.545 16.605 ;
      RECT 178.065 16.375 178.355 16.605 ;
      RECT 178.065 16.42 182.065 16.56 ;
      RECT 181.34 16.035 181.63 16.265 ;
      RECT 179.77 16.035 180.06 16.265 ;
      RECT 177.67 16.035 177.96 16.265 ;
      RECT 177.67 16.08 181.63 16.22 ;
      RECT 179.93 16.7 180.25 16.96 ;
      RECT 177.72 16.76 180.25 16.9 ;
      RECT 177.72 16.42 177.86 16.9 ;
      RECT 170.285 16.375 170.575 16.605 ;
      RECT 177.26 16.42 177.86 16.56 ;
      RECT 177.26 16.08 177.4 16.56 ;
      RECT 170.36 16.08 170.5 16.605 ;
      RECT 167.14 16.08 177.4 16.22 ;
      RECT 167.14 15.74 167.28 16.22 ;
      RECT 163.37 15.68 163.69 15.94 ;
      RECT 163.37 15.74 167.28 15.88 ;
      RECT 177.17 17.38 177.49 17.64 ;
      RECT 177.26 17.1 177.4 17.64 ;
      RECT 178.49 17.055 178.78 17.285 ;
      RECT 177.26 17.1 178.78 17.24 ;
      RECT 177.17 19.42 177.49 19.68 ;
      RECT 171.205 19.435 171.495 19.665 ;
      RECT 174.96 19.48 177.49 19.62 ;
      RECT 171.205 19.48 172.8 19.62 ;
      RECT 172.66 19.14 172.8 19.62 ;
      RECT 174.96 19.14 175.1 19.62 ;
      RECT 172.66 19.14 175.1 19.28 ;
      RECT 160.61 16.7 160.93 16.96 ;
      RECT 177.185 16.715 177.475 16.945 ;
      RECT 162.465 16.715 162.755 16.945 ;
      RECT 147.745 16.715 148.035 16.945 ;
      RECT 147.745 16.76 177.475 16.9 ;
      RECT 174.425 19.775 174.715 20.005 ;
      RECT 169.9 19.82 174.715 19.96 ;
      RECT 169.9 19.14 170.04 19.96 ;
      RECT 168.905 19.095 169.195 19.325 ;
      RECT 168.905 19.14 170.04 19.28 ;
      RECT 171.65 17.38 171.97 17.64 ;
      RECT 173.045 17.395 173.335 17.625 ;
      RECT 171.65 17.44 173.335 17.58 ;
      RECT 170.285 19.095 170.575 19.325 ;
      RECT 170.285 19.14 171.42 19.28 ;
      RECT 171.28 18.8 171.42 19.28 ;
      RECT 171.28 18.8 171.88 18.94 ;
      RECT 171.74 18.4 171.88 18.94 ;
      RECT 171.65 18.4 171.97 18.66 ;
      RECT 171.65 20.1 171.97 20.36 ;
      RECT 168.06 20.16 171.97 20.3 ;
      RECT 159.78 20.16 161.76 20.3 ;
      RECT 161.62 19.48 161.76 20.3 ;
      RECT 149.2 20.16 151.18 20.3 ;
      RECT 151.04 19.82 151.18 20.3 ;
      RECT 168.06 19.48 168.2 20.3 ;
      RECT 159.78 19.99 159.92 20.3 ;
      RECT 149.2 19.14 149.34 20.3 ;
      RECT 157.02 19.99 159.92 20.13 ;
      RECT 152.33 19.76 152.65 20.02 ;
      RECT 157.02 19.82 157.16 20.13 ;
      RECT 151.04 19.82 157.16 19.96 ;
      RECT 153.48 19.095 153.62 19.96 ;
      RECT 161.62 19.48 168.2 19.62 ;
      RECT 153.405 19.095 153.695 19.325 ;
      RECT 148.435 19.095 148.725 19.325 ;
      RECT 148.435 19.14 149.34 19.28 ;
      RECT 168.89 22.14 169.21 22.4 ;
      RECT 171.205 22.155 171.495 22.385 ;
      RECT 168.89 22.2 171.495 22.34 ;
      RECT 160.61 29.96 160.93 30.22 ;
      RECT 171.205 29.975 171.495 30.205 ;
      RECT 160.61 30.02 171.495 30.16 ;
      RECT 168.89 15.68 169.21 15.94 ;
      RECT 169.365 15.695 169.655 15.925 ;
      RECT 168.89 15.74 169.655 15.88 ;
      RECT 168.89 18.4 169.21 18.66 ;
      RECT 169.365 18.415 169.655 18.645 ;
      RECT 168.89 18.46 169.655 18.6 ;
      RECT 154.645 27.595 154.935 27.825 ;
      RECT 154.72 27.3 154.86 27.825 ;
      RECT 157.85 27.24 158.17 27.5 ;
      RECT 154.72 27.3 169.12 27.44 ;
      RECT 168.98 26.9 169.12 27.44 ;
      RECT 168.89 26.9 169.21 27.16 ;
      RECT 167.055 16.375 167.345 16.605 ;
      RECT 164.535 16.375 164.825 16.605 ;
      RECT 163.345 16.375 163.635 16.605 ;
      RECT 163.345 16.42 167.345 16.56 ;
      RECT 166.62 16.035 166.91 16.265 ;
      RECT 165.05 16.035 165.34 16.265 ;
      RECT 162.95 16.035 163.24 16.265 ;
      RECT 162.95 16.08 166.91 16.22 ;
      RECT 157.85 17.38 158.17 17.64 ;
      RECT 157.85 17.44 163.985 17.58 ;
      RECT 163.845 17.055 163.985 17.58 ;
      RECT 163.77 17.055 164.06 17.285 ;
      RECT 163.37 14.32 163.69 14.58 ;
      RECT 146.81 14.32 147.13 14.58 ;
      RECT 162.54 14.38 163.69 14.52 ;
      RECT 146.81 14.38 152.56 14.52 ;
      RECT 152.42 14.04 152.56 14.52 ;
      RECT 162.54 14.04 162.68 14.52 ;
      RECT 152.42 14.04 162.68 14.18 ;
      RECT 158.86 24.58 162.68 24.72 ;
      RECT 162.54 23.9 162.68 24.72 ;
      RECT 158.86 24.24 159 24.72 ;
      RECT 156.1 24.24 159 24.38 ;
      RECT 156.1 24.07 156.24 24.38 ;
      RECT 153.34 24.07 156.24 24.21 ;
      RECT 163.37 23.84 163.69 24.1 ;
      RECT 152.33 23.84 152.65 24.1 ;
      RECT 153.34 23.9 153.48 24.21 ;
      RECT 162.54 23.9 163.69 24.04 ;
      RECT 152.33 23.9 153.48 24.04 ;
      RECT 155.09 11.26 155.41 11.52 ;
      RECT 162.005 11.275 162.295 11.505 ;
      RECT 159.78 11.32 162.295 11.46 ;
      RECT 155.09 11.32 156.7 11.46 ;
      RECT 156.56 10.98 156.7 11.46 ;
      RECT 159.78 10.98 159.92 11.46 ;
      RECT 156.56 10.98 159.92 11.12 ;
      RECT 160.61 19.42 160.93 19.68 ;
      RECT 157.48 19.48 160.93 19.62 ;
      RECT 157.48 19.14 157.62 19.62 ;
      RECT 155.335 19.095 155.625 19.325 ;
      RECT 155.335 19.14 157.62 19.28 ;
      RECT 160.61 33.36 160.93 33.62 ;
      RECT 130.25 33.36 130.57 33.62 ;
      RECT 154.645 33.375 154.935 33.605 ;
      RECT 96.225 33.375 96.515 33.605 ;
      RECT 151.5 33.42 160.93 33.56 ;
      RECT 129.42 33.42 131.4 33.56 ;
      RECT 131.26 33.08 131.4 33.56 ;
      RECT 96.225 33.42 101.04 33.56 ;
      RECT 100.9 33.08 101.04 33.56 ;
      RECT 151.5 33.08 151.64 33.56 ;
      RECT 129.42 33.08 129.56 33.56 ;
      RECT 131.26 33.08 151.64 33.22 ;
      RECT 100.9 33.08 129.56 33.22 ;
      RECT 157.85 34.72 158.17 34.98 ;
      RECT 135.77 34.72 136.09 34.98 ;
      RECT 158.325 34.735 158.615 34.965 ;
      RECT 135.77 34.78 158.615 34.92 ;
      RECT 157.85 18.4 158.17 18.66 ;
      RECT 156.025 18.415 156.315 18.645 ;
      RECT 156.025 18.46 158.17 18.6 ;
      RECT 157.85 19.08 158.17 19.34 ;
      RECT 157.94 18.8 158.08 19.34 ;
      RECT 154.645 18.755 154.935 18.985 ;
      RECT 154.645 18.8 158.08 18.94 ;
      RECT 157.85 25.2 158.17 25.46 ;
      RECT 149.57 25.2 149.89 25.46 ;
      RECT 149.57 25.26 158.17 25.4 ;
      RECT 157.85 27.92 158.17 28.18 ;
      RECT 157.94 27.64 158.08 28.18 ;
      RECT 155.335 27.595 155.625 27.825 ;
      RECT 155.335 27.64 158.08 27.78 ;
      RECT 155.335 33.035 155.625 33.265 ;
      RECT 155.41 32.74 155.55 33.265 ;
      RECT 157.85 32.68 158.17 32.94 ;
      RECT 155.41 32.74 158.17 32.88 ;
      RECT 155.09 29.28 155.41 29.54 ;
      RECT 157.865 29.295 158.155 29.525 ;
      RECT 155.09 29.34 158.155 29.48 ;
      RECT 152.33 28.26 152.65 28.52 ;
      RECT 156.025 28.275 156.315 28.505 ;
      RECT 152.33 28.32 156.315 28.46 ;
      RECT 155.09 33.7 155.41 33.96 ;
      RECT 156.025 33.715 156.315 33.945 ;
      RECT 155.09 33.76 156.315 33.9 ;
      RECT 156.015 35.755 156.305 35.985 ;
      RECT 153.495 35.755 153.785 35.985 ;
      RECT 152.305 35.755 152.595 35.985 ;
      RECT 152.305 35.8 156.305 35.94 ;
      RECT 155.58 36.095 155.87 36.325 ;
      RECT 154.01 36.095 154.3 36.325 ;
      RECT 151.91 36.095 152.2 36.325 ;
      RECT 151.91 36.14 155.87 36.28 ;
      RECT 155.555 30.315 155.845 30.545 ;
      RECT 153.035 30.315 153.325 30.545 ;
      RECT 151.845 30.315 152.135 30.545 ;
      RECT 151.845 30.36 155.845 30.5 ;
      RECT 155.09 24.52 155.41 24.78 ;
      RECT 145.98 24.58 155.41 24.72 ;
      RECT 145.98 24.24 146.12 24.72 ;
      RECT 142.225 24.195 142.515 24.425 ;
      RECT 142.225 24.24 146.12 24.38 ;
      RECT 155.12 30.655 155.41 30.885 ;
      RECT 153.55 30.655 153.84 30.885 ;
      RECT 151.45 30.655 151.74 30.885 ;
      RECT 151.45 30.7 155.41 30.84 ;
      RECT 154.185 33.035 154.475 33.265 ;
      RECT 154.26 32.4 154.4 33.265 ;
      RECT 155.09 32.34 155.41 32.6 ;
      RECT 154.26 32.4 155.41 32.54 ;
      RECT 152.73 35.415 153.02 35.645 ;
      RECT 152.73 35.46 155.32 35.6 ;
      RECT 155.18 35.06 155.32 35.6 ;
      RECT 155.09 35.06 155.41 35.32 ;
      RECT 152.33 15.68 152.65 15.94 ;
      RECT 154.645 15.695 154.935 15.925 ;
      RECT 152.33 15.74 154.935 15.88 ;
      RECT 154.185 18.755 154.475 18.985 ;
      RECT 152.42 18.8 154.475 18.94 ;
      RECT 152.42 18.4 152.56 18.94 ;
      RECT 152.33 18.4 152.65 18.66 ;
      RECT 154.185 22.155 154.475 22.385 ;
      RECT 136.245 22.155 136.535 22.385 ;
      RECT 154.26 21.52 154.4 22.385 ;
      RECT 136.32 21.18 136.46 22.385 ;
      RECT 151.96 21.52 154.4 21.66 ;
      RECT 151.96 21.18 152.1 21.66 ;
      RECT 137.24 21.35 142.44 21.49 ;
      RECT 142.3 21.18 142.44 21.49 ;
      RECT 146.81 21.12 147.13 21.38 ;
      RECT 137.24 21.18 137.38 21.49 ;
      RECT 142.3 21.18 152.1 21.32 ;
      RECT 136.32 21.18 137.38 21.32 ;
      RECT 145.445 28.275 145.735 28.505 ;
      RECT 145.445 28.32 146.58 28.46 ;
      RECT 146.44 27.64 146.58 28.46 ;
      RECT 154.185 27.935 154.475 28.165 ;
      RECT 151.5 27.98 154.475 28.12 ;
      RECT 151.5 27.64 151.64 28.12 ;
      RECT 146.44 27.64 151.64 27.78 ;
      RECT 153.495 27.595 153.785 27.825 ;
      RECT 153.57 26.62 153.71 27.825 ;
      RECT 152.33 26.56 152.65 26.82 ;
      RECT 152.33 26.62 153.71 26.76 ;
      RECT 153.495 33.035 153.785 33.265 ;
      RECT 153.57 32.06 153.71 33.265 ;
      RECT 152.33 32 152.65 32.26 ;
      RECT 152.33 32.06 153.71 32.2 ;
      RECT 152.33 11.26 152.65 11.52 ;
      RECT 153.265 11.275 153.555 11.505 ;
      RECT 152.33 11.32 153.555 11.46 ;
      RECT 152.33 19.08 152.65 19.34 ;
      RECT 152.805 19.095 153.095 19.325 ;
      RECT 152.33 19.14 153.095 19.28 ;
      RECT 152.33 27.58 152.65 27.84 ;
      RECT 152.805 27.595 153.095 27.825 ;
      RECT 152.33 27.64 153.095 27.78 ;
      RECT 152.33 33.02 152.65 33.28 ;
      RECT 152.805 33.035 153.095 33.265 ;
      RECT 152.33 33.08 153.095 33.22 ;
      RECT 142.3 13.7 146.12 13.84 ;
      RECT 145.98 13.36 146.12 13.84 ;
      RECT 142.3 13.36 142.44 13.84 ;
      RECT 145.98 13.36 151.64 13.5 ;
      RECT 151.5 13.02 151.64 13.5 ;
      RECT 139.54 13.36 142.44 13.5 ;
      RECT 139.54 13.19 139.68 13.5 ;
      RECT 136.78 13.19 139.68 13.33 ;
      RECT 152.33 12.96 152.65 13.22 ;
      RECT 135.77 12.96 136.09 13.22 ;
      RECT 136.78 13.02 136.92 13.33 ;
      RECT 151.5 13.02 152.65 13.16 ;
      RECT 135.77 13.02 136.92 13.16 ;
      RECT 152.33 29.62 152.65 29.88 ;
      RECT 152.27 29.635 152.65 29.865 ;
      RECT 152.335 16.375 152.625 16.605 ;
      RECT 149.815 16.375 150.105 16.605 ;
      RECT 148.625 16.375 148.915 16.605 ;
      RECT 148.625 16.42 152.625 16.56 ;
      RECT 151.9 16.035 152.19 16.265 ;
      RECT 150.33 16.035 150.62 16.265 ;
      RECT 148.23 16.035 148.52 16.265 ;
      RECT 148.23 16.08 152.19 16.22 ;
      RECT 124.73 35.4 125.05 35.66 ;
      RECT 151.425 35.415 151.715 35.645 ;
      RECT 124.285 35.415 124.575 35.645 ;
      RECT 124.285 35.46 151.715 35.6 ;
      RECT 149.57 18.4 149.89 18.66 ;
      RECT 150.965 18.415 151.255 18.645 ;
      RECT 149.57 18.46 151.255 18.6 ;
      RECT 138.53 29.96 138.85 30.22 ;
      RECT 150.965 29.975 151.255 30.205 ;
      RECT 138.53 30.02 151.255 30.16 ;
      RECT 149.57 19.76 149.89 20.02 ;
      RECT 149.57 19.82 150.49 19.96 ;
      RECT 150.35 19.095 150.49 19.96 ;
      RECT 150.275 19.095 150.565 19.325 ;
      RECT 149.57 17.04 149.89 17.3 ;
      RECT 149.05 17.055 149.34 17.285 ;
      RECT 149.05 17.1 149.89 17.24 ;
      RECT 149.57 21.46 149.89 21.72 ;
      RECT 148.665 21.475 148.955 21.705 ;
      RECT 148.665 21.52 149.89 21.66 ;
      RECT 149.57 22.82 149.89 23.08 ;
      RECT 148.665 22.835 148.955 23.065 ;
      RECT 148.665 22.88 149.89 23.02 ;
      RECT 130.25 20.1 130.57 20.36 ;
      RECT 139.925 20.115 140.215 20.345 ;
      RECT 130.25 20.16 141.06 20.3 ;
      RECT 140.92 19.82 141.06 20.3 ;
      RECT 140.92 19.82 146.58 19.96 ;
      RECT 146.44 18.8 146.58 19.96 ;
      RECT 149.125 18.755 149.415 18.985 ;
      RECT 146.44 18.8 149.415 18.94 ;
      RECT 146.81 19.08 147.13 19.34 ;
      RECT 147.745 19.095 148.035 19.325 ;
      RECT 146.81 19.14 148.035 19.28 ;
      RECT 142.3 18.8 145.66 18.94 ;
      RECT 145.52 18.46 145.66 18.94 ;
      RECT 142.3 18.46 142.44 18.94 ;
      RECT 146.81 18.4 147.13 18.66 ;
      RECT 141.29 18.4 141.61 18.66 ;
      RECT 145.52 18.46 147.13 18.6 ;
      RECT 141.29 18.46 142.44 18.6 ;
      RECT 137.395 22.155 137.685 22.385 ;
      RECT 137.47 21.86 137.61 22.385 ;
      RECT 146.81 21.8 147.13 22.06 ;
      RECT 141.29 21.8 141.61 22.06 ;
      RECT 137.47 21.86 147.13 22 ;
      RECT 143.22 21.475 143.36 22 ;
      RECT 143.145 21.475 143.435 21.705 ;
      RECT 146.81 24.86 147.13 25.12 ;
      RECT 143.535 24.92 147.13 25.06 ;
      RECT 143.535 24.535 143.675 25.06 ;
      RECT 143.46 24.535 143.75 24.765 ;
      RECT 146.81 25.54 147.13 25.8 ;
      RECT 145.98 25.6 147.13 25.74 ;
      RECT 145.98 25.43 146.12 25.74 ;
      RECT 142.3 25.43 146.12 25.57 ;
      RECT 142.3 24.58 142.44 25.57 ;
      RECT 142.685 24.535 142.975 24.765 ;
      RECT 142.3 24.58 142.975 24.72 ;
      RECT 146.81 26.56 147.13 26.82 ;
      RECT 145.445 26.575 145.735 26.805 ;
      RECT 145.445 26.62 147.13 26.76 ;
      RECT 144.05 22.82 144.37 23.08 ;
      RECT 144.985 22.835 145.275 23.065 ;
      RECT 142.76 22.88 145.275 23.02 ;
      RECT 138.16 22.88 139.22 23.02 ;
      RECT 139.08 22.71 139.22 23.02 ;
      RECT 142.76 22.71 142.9 23.02 ;
      RECT 138.16 22.155 138.3 23.02 ;
      RECT 139.08 22.71 142.9 22.85 ;
      RECT 138.085 22.155 138.375 22.385 ;
      RECT 144.05 26.56 144.37 26.82 ;
      RECT 130.25 26.56 130.57 26.82 ;
      RECT 130.25 26.62 144.37 26.76 ;
      RECT 143.135 27.255 143.425 27.485 ;
      RECT 140.615 27.255 140.905 27.485 ;
      RECT 139.425 27.255 139.715 27.485 ;
      RECT 139.425 27.3 143.425 27.44 ;
      RECT 142.7 26.915 142.99 27.145 ;
      RECT 141.13 26.915 141.42 27.145 ;
      RECT 139.03 26.915 139.32 27.145 ;
      RECT 139.03 26.96 142.99 27.1 ;
      RECT 141.29 24.52 141.61 24.78 ;
      RECT 141.29 24.535 141.825 24.765 ;
      RECT 141.29 17.38 141.61 17.64 ;
      RECT 139.925 17.395 140.215 17.625 ;
      RECT 139.925 17.44 141.61 17.58 ;
      RECT 141.29 25.54 141.61 25.8 ;
      RECT 140.845 25.555 141.135 25.785 ;
      RECT 140.845 25.6 141.61 25.74 ;
      RECT 141.29 27.92 141.61 28.18 ;
      RECT 139.85 27.935 140.14 28.165 ;
      RECT 139.85 27.98 141.61 28.12 ;
      RECT 138.53 15.68 138.85 15.94 ;
      RECT 139.925 15.695 140.215 15.925 ;
      RECT 138.53 15.74 140.215 15.88 ;
      RECT 138.53 14.66 138.85 14.92 ;
      RECT 138.62 13.655 138.76 14.92 ;
      RECT 134.02 14.04 137.84 14.18 ;
      RECT 137.7 13.7 137.84 14.18 ;
      RECT 134.02 13.36 134.16 14.18 ;
      RECT 138.545 13.655 138.835 13.885 ;
      RECT 137.7 13.7 138.835 13.84 ;
      RECT 117.92 13.7 121.28 13.84 ;
      RECT 121.14 13.36 121.28 13.84 ;
      RECT 117.92 13.36 118.06 13.84 ;
      RECT 116.005 13.315 116.295 13.545 ;
      RECT 130.8 13.36 134.16 13.5 ;
      RECT 121.14 13.36 122.2 13.5 ;
      RECT 122.06 13.19 122.2 13.5 ;
      RECT 116.005 13.36 118.06 13.5 ;
      RECT 130.8 13.19 130.94 13.5 ;
      RECT 122.06 13.19 130.94 13.33 ;
      RECT 138.53 19.08 138.85 19.34 ;
      RECT 133.025 19.095 133.315 19.325 ;
      RECT 133.025 19.14 138.85 19.28 ;
      RECT 113.69 25.2 114.01 25.46 ;
      RECT 126.66 25.26 127.72 25.4 ;
      RECT 127.58 24.52 127.72 25.4 ;
      RECT 113.69 25.26 115.3 25.4 ;
      RECT 115.16 24.58 115.3 25.4 ;
      RECT 126.66 24.92 126.8 25.4 ;
      RECT 130.25 24.86 130.57 25.12 ;
      RECT 127.58 24.92 130.57 25.06 ;
      RECT 119.76 24.92 126.8 25.06 ;
      RECT 119.76 24.58 119.9 25.06 ;
      RECT 130.34 24.24 130.48 25.12 ;
      RECT 127.49 24.52 127.81 24.78 ;
      RECT 137.625 24.535 137.915 24.765 ;
      RECT 115.16 24.58 119.9 24.72 ;
      RECT 137.7 23.9 137.84 24.765 ;
      RECT 130.34 24.24 135.54 24.38 ;
      RECT 135.4 23.9 135.54 24.38 ;
      RECT 135.4 23.9 137.84 24.04 ;
      RECT 137.615 16.375 137.905 16.605 ;
      RECT 135.095 16.375 135.385 16.605 ;
      RECT 133.905 16.375 134.195 16.605 ;
      RECT 133.905 16.42 137.905 16.56 ;
      RECT 137.615 19.435 137.905 19.665 ;
      RECT 135.095 19.435 135.385 19.665 ;
      RECT 133.905 19.435 134.195 19.665 ;
      RECT 133.905 19.48 137.905 19.62 ;
      RECT 137.18 16.035 137.47 16.265 ;
      RECT 135.61 16.035 135.9 16.265 ;
      RECT 133.51 16.035 133.8 16.265 ;
      RECT 133.51 16.08 137.47 16.22 ;
      RECT 137.18 19.775 137.47 20.005 ;
      RECT 135.61 19.775 135.9 20.005 ;
      RECT 133.51 19.775 133.8 20.005 ;
      RECT 133.51 19.82 137.47 19.96 ;
      RECT 135.77 25.54 136.09 25.8 ;
      RECT 135.77 25.6 137.15 25.74 ;
      RECT 137.01 24.535 137.15 25.74 ;
      RECT 136.935 24.535 137.225 24.765 ;
      RECT 135.77 22.82 136.09 23.08 ;
      RECT 135.86 22.54 136 23.08 ;
      RECT 136.705 22.495 136.995 22.725 ;
      RECT 135.86 22.54 136.995 22.68 ;
      RECT 133.01 24.86 133.33 25.12 ;
      RECT 133.01 24.92 136.46 25.06 ;
      RECT 136.32 24.535 136.46 25.06 ;
      RECT 136.245 24.535 136.535 24.765 ;
      RECT 135.77 16.7 136.09 16.96 ;
      RECT 134.33 16.715 134.62 16.945 ;
      RECT 134.33 16.76 136.09 16.9 ;
      RECT 135.77 21.46 136.09 21.72 ;
      RECT 134.865 21.475 135.155 21.705 ;
      RECT 134.865 21.52 136.09 21.66 ;
      RECT 129.575 27.595 129.865 27.825 ;
      RECT 129.65 26.96 129.79 27.825 ;
      RECT 135.77 26.9 136.09 27.16 ;
      RECT 133.01 26.9 133.33 27.16 ;
      RECT 121.97 26.9 122.29 27.16 ;
      RECT 128.96 26.96 136.09 27.1 ;
      RECT 121.97 26.96 125.88 27.1 ;
      RECT 125.74 26.79 125.88 27.1 ;
      RECT 128.96 26.79 129.1 27.1 ;
      RECT 125.74 26.79 129.1 26.93 ;
      RECT 135.77 27.92 136.09 28.18 ;
      RECT 128.885 27.935 129.175 28.165 ;
      RECT 128.885 27.98 136.09 28.12 ;
      RECT 133.01 22.14 133.33 22.4 ;
      RECT 135.555 22.155 135.845 22.385 ;
      RECT 130.955 22.155 131.245 22.385 ;
      RECT 130.955 22.2 135.845 22.34 ;
      RECT 133.01 25.54 133.33 25.8 ;
      RECT 127.49 25.54 127.81 25.8 ;
      RECT 131.72 25.6 133.33 25.74 ;
      RECT 127.49 25.6 128.64 25.74 ;
      RECT 128.5 25.43 128.64 25.74 ;
      RECT 132.64 24.58 132.78 25.74 ;
      RECT 131.72 25.43 131.86 25.74 ;
      RECT 128.5 25.43 131.86 25.57 ;
      RECT 135.095 24.535 135.385 24.765 ;
      RECT 132.64 24.58 135.385 24.72 ;
      RECT 130.25 23.84 130.57 24.1 ;
      RECT 134.405 23.855 134.695 24.085 ;
      RECT 130.25 23.9 134.695 24.04 ;
      RECT 130.25 19.08 130.57 19.34 ;
      RECT 130.34 18.8 130.48 19.34 ;
      RECT 134.33 18.755 134.62 18.985 ;
      RECT 130.34 18.8 134.62 18.94 ;
      RECT 133.01 14.32 133.33 14.58 ;
      RECT 130.25 14.32 130.57 14.58 ;
      RECT 130.25 14.38 133.33 14.52 ;
      RECT 129.115 22.155 129.405 22.385 ;
      RECT 129.19 21.86 129.33 22.385 ;
      RECT 129.19 21.86 133.24 22 ;
      RECT 133.1 21.12 133.24 22 ;
      RECT 133.01 21.12 133.33 21.38 ;
      RECT 133.01 22.82 133.33 23.08 ;
      RECT 132.105 22.835 132.395 23.065 ;
      RECT 132.105 22.88 133.33 23.02 ;
      RECT 127.49 21.12 127.81 21.38 ;
      RECT 132.105 21.135 132.395 21.365 ;
      RECT 127.965 21.135 128.255 21.365 ;
      RECT 127.49 21.18 132.395 21.32 ;
      RECT 131.645 22.835 131.935 23.065 ;
      RECT 122.445 22.88 131.935 23.02 ;
      RECT 122.445 22.495 122.585 23.02 ;
      RECT 122.37 22.495 122.66 22.725 ;
      RECT 130.25 34.72 130.57 34.98 ;
      RECT 131.185 34.735 131.475 34.965 ;
      RECT 130.25 34.78 131.475 34.92 ;
      RECT 130.25 28.26 130.57 28.52 ;
      RECT 127.045 28.275 127.335 28.505 ;
      RECT 128.5 28.32 130.57 28.46 ;
      RECT 128.5 27.98 128.64 28.46 ;
      RECT 127.12 27.98 127.26 28.505 ;
      RECT 127.12 27.98 128.64 28.12 ;
      RECT 130.25 29.28 130.57 29.54 ;
      RECT 127.49 29.28 127.81 29.54 ;
      RECT 127.49 29.34 130.57 29.48 ;
      RECT 111.02 22.71 115.76 22.85 ;
      RECT 115.62 22.54 115.76 22.85 ;
      RECT 119.21 22.48 119.53 22.74 ;
      RECT 129.805 22.495 130.095 22.725 ;
      RECT 110.025 22.495 110.315 22.725 ;
      RECT 111.02 22.54 111.16 22.85 ;
      RECT 126.2 22.54 130.095 22.68 ;
      RECT 115.62 22.54 120.82 22.68 ;
      RECT 120.68 21.18 120.82 22.68 ;
      RECT 110.025 22.54 111.16 22.68 ;
      RECT 126.2 21.18 126.34 22.68 ;
      RECT 120.68 21.18 126.34 21.32 ;
      RECT 128.875 35.755 129.165 35.985 ;
      RECT 126.355 35.755 126.645 35.985 ;
      RECT 125.165 35.755 125.455 35.985 ;
      RECT 125.165 35.8 129.165 35.94 ;
      RECT 128.44 36.095 128.73 36.325 ;
      RECT 126.87 36.095 127.16 36.325 ;
      RECT 124.77 36.095 125.06 36.325 ;
      RECT 124.77 36.14 128.73 36.28 ;
      RECT 127.49 22.14 127.81 22.4 ;
      RECT 128.425 22.155 128.715 22.385 ;
      RECT 127.49 22.2 128.715 22.34 ;
      RECT 102.65 28.26 102.97 28.52 ;
      RECT 109.64 28.32 112.08 28.46 ;
      RECT 111.94 28.15 112.08 28.46 ;
      RECT 102.65 28.32 103.8 28.46 ;
      RECT 103.66 27.98 103.8 28.46 ;
      RECT 109.64 27.98 109.78 28.46 ;
      RECT 111.94 28.15 117.6 28.29 ;
      RECT 117.46 27.64 117.6 28.29 ;
      RECT 121.14 27.98 125.88 28.12 ;
      RECT 125.74 27.3 125.88 28.12 ;
      RECT 103.66 27.98 109.78 28.12 ;
      RECT 121.14 27.64 121.28 28.12 ;
      RECT 128.425 27.595 128.715 27.825 ;
      RECT 117.46 27.64 121.28 27.78 ;
      RECT 128.5 27.3 128.64 27.825 ;
      RECT 125.74 27.3 128.64 27.44 ;
      RECT 127.49 27.58 127.81 27.84 ;
      RECT 127.49 27.595 128.025 27.825 ;
      RECT 125.59 35.075 125.88 35.305 ;
      RECT 125.665 34.78 125.805 35.305 ;
      RECT 127.49 34.72 127.81 34.98 ;
      RECT 125.665 34.78 127.81 34.92 ;
      RECT 125.655 21.815 125.945 22.045 ;
      RECT 123.135 21.815 123.425 22.045 ;
      RECT 121.945 21.815 122.235 22.045 ;
      RECT 121.945 21.86 125.945 22 ;
      RECT 125.22 21.475 125.51 21.705 ;
      RECT 123.65 21.475 123.94 21.705 ;
      RECT 121.55 21.475 121.84 21.705 ;
      RECT 121.55 21.52 125.51 21.66 ;
      RECT 124.73 15.68 125.05 15.94 ;
      RECT 125.205 15.695 125.495 15.925 ;
      RECT 124.73 15.74 125.495 15.88 ;
      RECT 125.205 17.395 125.495 17.625 ;
      RECT 124.36 17.44 125.495 17.58 ;
      RECT 118.38 17.44 120.36 17.58 ;
      RECT 120.22 17.27 120.36 17.58 ;
      RECT 124.36 17.27 124.5 17.58 ;
      RECT 118.38 17.1 118.52 17.58 ;
      RECT 120.22 17.27 124.5 17.41 ;
      RECT 114.625 17.055 114.915 17.285 ;
      RECT 114.625 17.1 118.52 17.24 ;
      RECT 124.73 22.14 125.05 22.4 ;
      RECT 121.065 22.155 121.355 22.385 ;
      RECT 121.065 22.2 125.05 22.34 ;
      RECT 121.97 19.08 122.29 19.34 ;
      RECT 124.745 19.095 125.035 19.325 ;
      RECT 120.605 19.095 120.895 19.325 ;
      RECT 120.605 19.14 125.035 19.28 ;
      RECT 119.64 16.715 119.93 16.945 ;
      RECT 119.64 16.76 123.58 16.9 ;
      RECT 123.44 15.74 123.58 16.9 ;
      RECT 119.21 15.68 119.53 15.94 ;
      RECT 119.21 15.74 123.58 15.88 ;
      RECT 122.895 16.375 123.185 16.605 ;
      RECT 120.375 16.375 120.665 16.605 ;
      RECT 119.185 16.375 119.475 16.605 ;
      RECT 119.185 16.42 123.185 16.56 ;
      RECT 122.46 16.035 122.75 16.265 ;
      RECT 120.89 16.035 121.18 16.265 ;
      RECT 118.79 16.035 119.08 16.265 ;
      RECT 118.79 16.08 122.75 16.22 ;
      RECT 119.21 14.66 119.53 14.92 ;
      RECT 117.385 14.675 117.675 14.905 ;
      RECT 117.385 14.72 119.53 14.86 ;
      RECT 119.21 17.04 119.53 17.3 ;
      RECT 119.3 16.76 119.44 17.3 ;
      RECT 118.305 16.715 118.595 16.945 ;
      RECT 118.305 16.76 119.44 16.9 ;
      RECT 116.005 22.155 116.295 22.385 ;
      RECT 116.08 21.86 116.22 22.385 ;
      RECT 119.21 21.8 119.53 22.06 ;
      RECT 116.08 21.86 119.53 22 ;
      RECT 119.21 25.54 119.53 25.8 ;
      RECT 113.32 25.6 119.53 25.74 ;
      RECT 113.32 24.535 113.46 25.74 ;
      RECT 113.245 24.535 113.535 24.765 ;
      RECT 119.21 26.56 119.53 26.82 ;
      RECT 117.385 26.575 117.675 26.805 ;
      RECT 117.385 26.62 119.53 26.76 ;
      RECT 116.45 22.82 116.77 23.08 ;
      RECT 117.385 22.835 117.675 23.065 ;
      RECT 116.45 22.88 117.675 23.02 ;
      RECT 116.45 20.1 116.77 20.36 ;
      RECT 116.925 20.115 117.215 20.345 ;
      RECT 105.04 20.16 117.215 20.3 ;
      RECT 105.04 19.48 105.18 20.3 ;
      RECT 105.04 19.48 106.56 19.62 ;
      RECT 106.42 19.095 106.56 19.62 ;
      RECT 106.345 19.095 106.635 19.325 ;
      RECT 108.17 14.32 108.49 14.58 ;
      RECT 105.41 14.32 105.73 14.58 ;
      RECT 105.41 14.38 116.91 14.52 ;
      RECT 116.77 13.655 116.91 14.52 ;
      RECT 116.695 13.655 116.985 13.885 ;
      RECT 116.45 22.14 116.77 22.4 ;
      RECT 116.45 22.155 116.985 22.385 ;
      RECT 116.45 11.26 116.77 11.52 ;
      RECT 115.085 11.275 115.375 11.505 ;
      RECT 115.085 11.32 116.77 11.46 ;
      RECT 115.545 13.315 115.835 13.545 ;
      RECT 115.62 13.02 115.76 13.545 ;
      RECT 116.45 12.96 116.77 13.22 ;
      RECT 115.62 13.02 116.77 13.16 ;
      RECT 116.45 16.7 116.77 16.96 ;
      RECT 115.315 16.715 115.605 16.945 ;
      RECT 115.315 16.76 116.77 16.9 ;
      RECT 116.45 17.38 116.77 17.64 ;
      RECT 116.005 17.395 116.295 17.625 ;
      RECT 116.005 17.44 116.77 17.58 ;
      RECT 116.45 19.08 116.77 19.34 ;
      RECT 111.36 19.095 111.65 19.325 ;
      RECT 115.62 19.14 116.77 19.28 ;
      RECT 111.36 19.14 112.54 19.28 ;
      RECT 112.4 18.97 112.54 19.28 ;
      RECT 115.62 18.97 115.76 19.28 ;
      RECT 112.4 18.97 115.76 19.11 ;
      RECT 116.45 27.58 116.77 27.84 ;
      RECT 111.79 27.595 112.08 27.825 ;
      RECT 111.79 27.64 116.77 27.78 ;
      RECT 115.545 22.155 115.835 22.385 ;
      RECT 115.62 21.18 115.76 22.385 ;
      RECT 111.02 21.35 114.84 21.49 ;
      RECT 114.7 21.18 114.84 21.49 ;
      RECT 105.41 21.12 105.73 21.38 ;
      RECT 111.02 21.18 111.16 21.49 ;
      RECT 114.7 21.18 115.76 21.32 ;
      RECT 105.41 21.18 111.16 21.32 ;
      RECT 115.075 27.255 115.365 27.485 ;
      RECT 112.555 27.255 112.845 27.485 ;
      RECT 111.365 27.255 111.655 27.485 ;
      RECT 111.365 27.3 115.365 27.44 ;
      RECT 105.41 13.64 105.73 13.9 ;
      RECT 114.855 13.655 115.145 13.885 ;
      RECT 105.41 13.7 106.1 13.84 ;
      RECT 105.96 13.36 106.1 13.84 ;
      RECT 114.93 13.36 115.07 13.885 ;
      RECT 110.93 13.3 111.25 13.56 ;
      RECT 105.96 13.36 115.07 13.5 ;
      RECT 111.315 22.14 111.635 22.4 ;
      RECT 114.855 22.155 115.145 22.385 ;
      RECT 114.93 21.86 115.07 22.385 ;
      RECT 111.405 21.86 111.545 22.4 ;
      RECT 111.405 21.86 115.07 22 ;
      RECT 114.64 26.915 114.93 27.145 ;
      RECT 113.07 26.915 113.36 27.145 ;
      RECT 110.97 26.915 111.26 27.145 ;
      RECT 110.97 26.96 114.93 27.1 ;
      RECT 114.615 19.435 114.905 19.665 ;
      RECT 112.095 19.435 112.385 19.665 ;
      RECT 110.905 19.435 111.195 19.665 ;
      RECT 110.905 19.48 114.905 19.62 ;
      RECT 114.18 19.775 114.47 20.005 ;
      RECT 112.61 19.775 112.9 20.005 ;
      RECT 110.51 19.775 110.8 20.005 ;
      RECT 110.51 19.82 114.47 19.96 ;
      RECT 113.69 13.64 114.01 13.9 ;
      RECT 114.165 13.655 114.455 13.885 ;
      RECT 113.69 13.7 114.455 13.84 ;
      RECT 114.165 16.715 114.455 16.945 ;
      RECT 114.24 15.74 114.38 16.945 ;
      RECT 98.6 16.08 101.5 16.22 ;
      RECT 101.36 15.74 101.5 16.22 ;
      RECT 98.6 15.74 98.74 16.22 ;
      RECT 97.13 15.68 97.45 15.94 ;
      RECT 110.485 15.695 110.775 15.925 ;
      RECT 101.36 15.74 114.38 15.88 ;
      RECT 97.13 15.74 98.74 15.88 ;
      RECT 113.69 22.14 114.01 22.4 ;
      RECT 114.165 22.155 114.455 22.385 ;
      RECT 111.865 22.155 112.155 22.385 ;
      RECT 111.865 22.2 114.455 22.34 ;
      RECT 100.9 30.02 106.56 30.16 ;
      RECT 106.42 29.34 106.56 30.16 ;
      RECT 100.9 29.34 101.04 30.16 ;
      RECT 99.89 29.28 100.21 29.54 ;
      RECT 114.165 29.295 114.455 29.525 ;
      RECT 106.42 29.34 114.455 29.48 ;
      RECT 99.89 29.34 101.04 29.48 ;
      RECT 113.69 17.38 114.01 17.64 ;
      RECT 112.86 17.44 114.01 17.58 ;
      RECT 112.86 16.715 113 17.58 ;
      RECT 112.785 16.715 113.075 16.945 ;
      RECT 108.185 19.095 108.475 19.325 ;
      RECT 108.185 19.14 109.78 19.28 ;
      RECT 109.64 18.46 109.78 19.28 ;
      RECT 113.69 18.4 114.01 18.66 ;
      RECT 109.64 18.46 114.01 18.6 ;
      RECT 89.86 27.3 109.78 27.44 ;
      RECT 109.64 26.62 109.78 27.44 ;
      RECT 89.86 26.62 90 27.44 ;
      RECT 113.69 26.56 114.01 26.82 ;
      RECT 88.85 26.56 89.17 26.82 ;
      RECT 109.64 26.62 114.01 26.76 ;
      RECT 88.85 26.62 90 26.76 ;
      RECT 113.475 16.715 113.765 16.945 ;
      RECT 113.55 16.42 113.69 16.945 ;
      RECT 110.93 16.36 111.25 16.62 ;
      RECT 110.93 16.42 113.69 16.56 ;
      RECT 111.855 30.315 112.145 30.545 ;
      RECT 109.335 30.315 109.625 30.545 ;
      RECT 108.145 30.315 108.435 30.545 ;
      RECT 108.145 30.36 112.145 30.5 ;
      RECT 111.42 30.655 111.71 30.885 ;
      RECT 109.85 30.655 110.14 30.885 ;
      RECT 107.75 30.655 108.04 30.885 ;
      RECT 107.75 30.7 111.71 30.84 ;
      RECT 110.025 19.095 110.315 19.325 ;
      RECT 110.025 19.14 111.16 19.28 ;
      RECT 111.02 18.74 111.16 19.28 ;
      RECT 110.93 18.74 111.25 19 ;
      RECT 110.93 27.58 111.25 27.84 ;
      RECT 110.485 27.595 110.775 27.825 ;
      RECT 110.485 27.64 111.25 27.78 ;
      RECT 110.93 29.96 111.25 30.22 ;
      RECT 107.265 29.975 107.555 30.205 ;
      RECT 107.265 30.02 111.25 30.16 ;
      RECT 110.485 22.155 110.775 22.385 ;
      RECT 110.1 22.2 110.775 22.34 ;
      RECT 103.66 22.2 107.48 22.34 ;
      RECT 107.34 21.52 107.48 22.34 ;
      RECT 110.1 21.52 110.24 22.34 ;
      RECT 103.66 21.52 103.8 22.34 ;
      RECT 107.34 21.52 110.24 21.66 ;
      RECT 100.44 21.52 103.8 21.66 ;
      RECT 100.44 21.135 100.58 21.66 ;
      RECT 97.13 21.12 97.45 21.38 ;
      RECT 100.365 21.135 100.655 21.365 ;
      RECT 97.13 21.18 100.655 21.32 ;
      RECT 108.17 22.14 108.49 22.4 ;
      RECT 109.335 22.155 109.625 22.385 ;
      RECT 108.17 22.2 109.625 22.34 ;
      RECT 108.17 22.82 108.49 23.08 ;
      RECT 108.645 22.835 108.935 23.065 ;
      RECT 108.17 22.88 108.935 23.02 ;
      RECT 108.17 17.38 108.49 17.64 ;
      RECT 108.26 16.76 108.4 17.64 ;
      RECT 104.89 16.715 105.18 16.945 ;
      RECT 104.89 16.76 108.4 16.9 ;
      RECT 108.17 18.4 108.49 18.66 ;
      RECT 104.965 18.415 105.255 18.645 ;
      RECT 104.965 18.46 108.49 18.6 ;
      RECT 108.175 16.375 108.465 16.605 ;
      RECT 105.655 16.375 105.945 16.605 ;
      RECT 104.465 16.375 104.755 16.605 ;
      RECT 104.465 16.42 108.465 16.56 ;
      RECT 107.74 16.035 108.03 16.265 ;
      RECT 106.17 16.035 106.46 16.265 ;
      RECT 104.07 16.035 104.36 16.265 ;
      RECT 104.07 16.08 108.03 16.22 ;
      RECT 105.41 19.76 105.73 20.02 ;
      RECT 105.41 19.82 107.02 19.96 ;
      RECT 106.88 19.14 107.02 19.96 ;
      RECT 107.495 19.095 107.785 19.325 ;
      RECT 106.88 19.14 107.785 19.28 ;
      RECT 99.89 18.74 100.21 19 ;
      RECT 106.805 18.755 107.095 18.985 ;
      RECT 99.89 18.8 107.095 18.94 ;
      RECT 91.61 20.1 91.93 20.36 ;
      RECT 84.11 20.16 97.82 20.3 ;
      RECT 97.68 19.48 97.82 20.3 ;
      RECT 84.11 19.095 84.25 20.3 ;
      RECT 98.6 19.48 104.26 19.62 ;
      RECT 104.12 19.14 104.26 19.62 ;
      RECT 97.45 19.48 97.82 19.62 ;
      RECT 98.6 19.14 98.74 19.62 ;
      RECT 97.45 19.095 97.59 19.62 ;
      RECT 105.41 19.08 105.73 19.34 ;
      RECT 105.41 19.095 105.945 19.325 ;
      RECT 97.375 19.095 97.665 19.325 ;
      RECT 84.035 19.095 84.325 19.325 ;
      RECT 104.12 19.14 105.945 19.28 ;
      RECT 97.375 19.14 98.74 19.28 ;
      RECT 105.41 25.54 105.73 25.8 ;
      RECT 104.58 25.6 105.73 25.74 ;
      RECT 104.58 25.26 104.72 25.74 ;
      RECT 96.3 25.43 101.04 25.57 ;
      RECT 100.9 25.26 101.04 25.57 ;
      RECT 86.09 25.2 86.41 25.46 ;
      RECT 96.3 25.26 96.44 25.57 ;
      RECT 100.9 25.26 104.72 25.4 ;
      RECT 85.26 25.26 96.44 25.4 ;
      RECT 95.61 24.535 95.75 25.4 ;
      RECT 85.26 24.92 85.4 25.4 ;
      RECT 84.57 24.92 85.4 25.06 ;
      RECT 84.57 24.535 84.71 25.06 ;
      RECT 95.535 24.535 95.825 24.765 ;
      RECT 84.495 24.535 84.785 24.765 ;
      RECT 99.89 11.6 100.21 11.86 ;
      RECT 99.89 11.66 100.58 11.8 ;
      RECT 100.44 11.32 100.58 11.8 ;
      RECT 103.585 11.275 103.875 11.505 ;
      RECT 100.44 11.32 103.875 11.46 ;
      RECT 102.65 16.7 102.97 16.96 ;
      RECT 103.585 16.715 103.875 16.945 ;
      RECT 102.65 16.76 103.875 16.9 ;
      RECT 93.54 22.88 97.82 23.02 ;
      RECT 97.68 22.2 97.82 23.02 ;
      RECT 93.54 22.54 93.68 23.02 ;
      RECT 88.85 22.48 89.17 22.74 ;
      RECT 83.33 22.48 83.65 22.74 ;
      RECT 83.33 22.54 93.68 22.68 ;
      RECT 86.64 22.155 86.78 22.68 ;
      RECT 102.65 22.14 102.97 22.4 ;
      RECT 86.565 22.155 86.855 22.385 ;
      RECT 97.68 22.2 102.97 22.34 ;
      RECT 102.65 24.18 102.97 24.44 ;
      RECT 96.225 24.195 96.515 24.425 ;
      RECT 96.225 24.24 102.97 24.38 ;
      RECT 80.2 35.46 90.92 35.6 ;
      RECT 90.78 34.78 90.92 35.6 ;
      RECT 48.46 35.46 79.42 35.6 ;
      RECT 79.28 34.78 79.42 35.6 ;
      RECT 80.2 34.78 80.34 35.6 ;
      RECT 48.46 35.12 48.6 35.6 ;
      RECT 47.54 35.12 48.6 35.26 ;
      RECT 47.54 34.72 47.68 35.26 ;
      RECT 102.65 34.72 102.97 34.98 ;
      RECT 47.45 34.72 47.77 34.98 ;
      RECT 99.905 34.735 100.195 34.965 ;
      RECT 90.78 34.78 102.97 34.92 ;
      RECT 79.28 34.78 80.34 34.92 ;
      RECT 99.89 17.38 100.21 17.64 ;
      RECT 100.825 17.395 101.115 17.625 ;
      RECT 99.89 17.44 101.115 17.58 ;
      RECT 83.33 13.98 83.65 14.24 ;
      RECT 65.48 14.04 84.48 14.18 ;
      RECT 84.34 13.7 84.48 14.18 ;
      RECT 65.48 13.655 65.62 14.18 ;
      RECT 99.89 13.64 100.21 13.9 ;
      RECT 65.405 13.655 65.695 13.885 ;
      RECT 84.34 13.7 100.21 13.84 ;
      RECT 99.89 24.86 100.21 25.12 ;
      RECT 96.76 24.92 100.21 25.06 ;
      RECT 96.76 24.535 96.9 25.06 ;
      RECT 96.685 24.535 96.975 24.765 ;
      RECT 96.685 33.035 96.975 33.265 ;
      RECT 96.76 32.74 96.9 33.265 ;
      RECT 99.89 32.68 100.21 32.94 ;
      RECT 96.76 32.74 100.21 32.88 ;
      RECT 98.515 16.375 98.805 16.605 ;
      RECT 95.995 16.375 96.285 16.605 ;
      RECT 94.805 16.375 95.095 16.605 ;
      RECT 94.805 16.42 98.805 16.56 ;
      RECT 98.08 16.035 98.37 16.265 ;
      RECT 96.51 16.035 96.8 16.265 ;
      RECT 94.41 16.035 94.7 16.265 ;
      RECT 94.41 16.08 98.37 16.22 ;
      RECT 97.13 18.4 97.45 18.66 ;
      RECT 98.065 18.415 98.355 18.645 ;
      RECT 97.13 18.46 98.355 18.6 ;
      RECT 97.13 23.84 97.45 24.1 ;
      RECT 98.065 23.855 98.355 24.085 ;
      RECT 97.13 23.9 98.355 24.04 ;
      RECT 97.13 33.7 97.45 33.96 ;
      RECT 98.065 33.715 98.355 33.945 ;
      RECT 97.13 33.76 98.355 33.9 ;
      RECT 98.055 21.815 98.345 22.045 ;
      RECT 95.535 21.815 95.825 22.045 ;
      RECT 94.345 21.815 94.635 22.045 ;
      RECT 94.345 21.86 98.345 22 ;
      RECT 97.62 21.475 97.91 21.705 ;
      RECT 96.05 21.475 96.34 21.705 ;
      RECT 93.95 21.475 94.24 21.705 ;
      RECT 93.95 21.52 97.91 21.66 ;
      RECT 97.595 35.755 97.885 35.985 ;
      RECT 95.075 35.755 95.365 35.985 ;
      RECT 93.885 35.755 94.175 35.985 ;
      RECT 93.885 35.8 97.885 35.94 ;
      RECT 97.13 24.52 97.45 24.78 ;
      RECT 97.13 24.535 97.665 24.765 ;
      RECT 97.13 33.02 97.45 33.28 ;
      RECT 97.13 33.035 97.665 33.265 ;
      RECT 97.13 16.7 97.45 16.96 ;
      RECT 95.23 16.715 95.52 16.945 ;
      RECT 95.23 16.76 97.45 16.9 ;
      RECT 97.13 19.76 97.45 20.02 ;
      RECT 96.76 19.82 97.45 19.96 ;
      RECT 96.76 19.095 96.9 19.96 ;
      RECT 96.685 19.095 96.975 19.325 ;
      RECT 97.13 22.14 97.45 22.4 ;
      RECT 94.8 22.155 95.09 22.385 ;
      RECT 94.8 22.2 97.45 22.34 ;
      RECT 97.13 35.06 97.45 35.32 ;
      RECT 94.34 35.075 94.63 35.305 ;
      RECT 94.34 35.12 97.45 35.26 ;
      RECT 97.16 36.095 97.45 36.325 ;
      RECT 95.59 36.095 95.88 36.325 ;
      RECT 93.49 36.095 93.78 36.325 ;
      RECT 93.49 36.14 97.45 36.28 ;
      RECT 96.225 18.755 96.515 18.985 ;
      RECT 95.38 18.8 96.515 18.94 ;
      RECT 95.38 18.63 95.52 18.94 ;
      RECT 89.4 18.63 95.52 18.77 ;
      RECT 86.09 18.4 86.41 18.66 ;
      RECT 89.4 18.46 89.54 18.77 ;
      RECT 86.09 18.46 89.54 18.6 ;
      RECT 89.86 19.65 95.06 19.79 ;
      RECT 94.92 19.48 95.06 19.79 ;
      RECT 89.86 19.48 90 19.79 ;
      RECT 94.92 19.48 95.75 19.62 ;
      RECT 95.61 19.095 95.75 19.62 ;
      RECT 86.18 19.48 90 19.62 ;
      RECT 86.18 19.08 86.32 19.62 ;
      RECT 86.09 19.08 86.41 19.34 ;
      RECT 95.535 19.095 95.825 19.325 ;
      RECT 85.96 19.095 86.41 19.325 ;
      RECT 86.64 33.42 95.75 33.56 ;
      RECT 95.61 33.035 95.75 33.56 ;
      RECT 86.64 32.06 86.78 33.56 ;
      RECT 95.535 33.035 95.825 33.265 ;
      RECT 86.09 32 86.41 32.26 ;
      RECT 86.09 32.06 86.78 32.2 ;
      RECT 88.85 19.08 89.17 19.34 ;
      RECT 94.845 19.095 95.135 19.325 ;
      RECT 86.565 19.095 86.855 19.325 ;
      RECT 86.565 19.14 95.135 19.28 ;
      RECT 88.85 24.86 89.17 25.12 ;
      RECT 87.1 24.92 90.46 25.06 ;
      RECT 90.32 24.58 90.46 25.06 ;
      RECT 87.1 24.58 87.24 25.06 ;
      RECT 94.845 24.535 95.135 24.765 ;
      RECT 85.185 24.535 85.475 24.765 ;
      RECT 78.745 24.535 79.035 24.765 ;
      RECT 70.465 24.535 70.755 24.765 ;
      RECT 90.32 24.58 95.135 24.72 ;
      RECT 85.185 24.58 87.24 24.72 ;
      RECT 85.26 23.9 85.4 24.765 ;
      RECT 78.82 23.9 78.96 24.765 ;
      RECT 70.54 23.9 70.68 24.765 ;
      RECT 72.29 23.84 72.61 24.1 ;
      RECT 70.54 23.9 85.4 24.04 ;
      RECT 94.845 33.035 95.135 33.265 ;
      RECT 94.92 32.06 95.06 33.265 ;
      RECT 89.86 32.4 94.14 32.54 ;
      RECT 94 32.06 94.14 32.54 ;
      RECT 89.86 32.06 90 32.54 ;
      RECT 88.85 32 89.17 32.26 ;
      RECT 94 32.06 95.06 32.2 ;
      RECT 88.85 32.06 90 32.2 ;
      RECT 94.37 16.7 94.69 16.96 ;
      RECT 93.925 16.715 94.215 16.945 ;
      RECT 93.925 16.76 94.69 16.9 ;
      RECT 94.37 22.48 94.69 22.74 ;
      RECT 94.46 22.2 94.6 22.74 ;
      RECT 93.465 22.155 93.755 22.385 ;
      RECT 93.465 22.2 94.6 22.34 ;
      RECT 91.61 35.4 91.93 35.66 ;
      RECT 93.005 35.415 93.295 35.645 ;
      RECT 91.61 35.46 93.295 35.6 ;
      RECT 67.475 22.155 67.765 22.385 ;
      RECT 69.16 22.2 74.36 22.34 ;
      RECT 74.22 21.86 74.36 22.34 ;
      RECT 66.86 22.2 67.765 22.34 ;
      RECT 69.16 21.86 69.3 22.34 ;
      RECT 66.86 21.8 67 22.34 ;
      RECT 66.77 21.8 67.09 22.06 ;
      RECT 74.22 21.86 79.88 22 ;
      RECT 79.74 21.52 79.88 22 ;
      RECT 66.77 21.86 69.3 22 ;
      RECT 91.61 21.46 91.93 21.72 ;
      RECT 86.64 21.52 91.93 21.66 ;
      RECT 79.74 21.52 80.8 21.66 ;
      RECT 80.66 21.35 80.8 21.66 ;
      RECT 86.64 21.35 86.78 21.66 ;
      RECT 80.66 21.35 86.78 21.49 ;
      RECT 91.61 25.54 91.93 25.8 ;
      RECT 82.5 25.6 91.93 25.74 ;
      RECT 82.5 25.26 82.64 25.74 ;
      RECT 68.24 25.43 74.82 25.57 ;
      RECT 74.68 25.26 74.82 25.57 ;
      RECT 66.77 25.2 67.09 25.46 ;
      RECT 68.24 25.26 68.38 25.57 ;
      RECT 74.68 25.26 82.64 25.4 ;
      RECT 66.77 25.26 68.38 25.4 ;
      RECT 82.04 24.58 82.18 25.4 ;
      RECT 76.445 24.535 76.585 25.4 ;
      RECT 82.655 24.535 82.945 24.765 ;
      RECT 76.37 24.535 76.66 24.765 ;
      RECT 82.04 24.58 82.945 24.72 ;
      RECT 88.85 15.68 89.17 15.94 ;
      RECT 87.945 15.695 88.235 15.925 ;
      RECT 87.945 15.74 89.17 15.88 ;
      RECT 88.85 19.76 89.17 20.02 ;
      RECT 85.26 19.82 89.17 19.96 ;
      RECT 85.26 19.14 85.4 19.96 ;
      RECT 84.725 19.095 85.015 19.325 ;
      RECT 84.725 19.14 85.4 19.28 ;
      RECT 86.09 17.38 86.41 17.64 ;
      RECT 80.2 17.44 86.41 17.58 ;
      RECT 80.2 16.76 80.34 17.58 ;
      RECT 75.05 16.7 75.37 16.96 ;
      RECT 73.685 16.715 73.975 16.945 ;
      RECT 73.685 16.76 80.34 16.9 ;
      RECT 28.13 33.36 28.45 33.62 ;
      RECT 28.13 33.42 41.7 33.56 ;
      RECT 41.56 33.08 41.7 33.56 ;
      RECT 36.5 33.035 36.64 33.56 ;
      RECT 86.09 33.02 86.41 33.28 ;
      RECT 36.425 33.035 36.715 33.265 ;
      RECT 74.22 33.08 86.41 33.22 ;
      RECT 41.56 33.08 69.3 33.22 ;
      RECT 69.16 32.74 69.3 33.22 ;
      RECT 74.22 32.74 74.36 33.22 ;
      RECT 69.16 32.74 74.36 32.88 ;
      RECT 85.635 16.375 85.925 16.605 ;
      RECT 83.115 16.375 83.405 16.605 ;
      RECT 81.925 16.375 82.215 16.605 ;
      RECT 81.925 16.42 85.925 16.56 ;
      RECT 85.2 16.035 85.49 16.265 ;
      RECT 83.63 16.035 83.92 16.265 ;
      RECT 81.53 16.035 81.82 16.265 ;
      RECT 81.53 16.08 85.49 16.22 ;
      RECT 80.57 19.76 80.89 20.02 ;
      RECT 80.57 19.82 83.1 19.96 ;
      RECT 82.96 18.8 83.1 19.96 ;
      RECT 85.185 18.755 85.475 18.985 ;
      RECT 82.96 18.8 85.475 18.94 ;
      RECT 83.33 26.56 83.65 26.82 ;
      RECT 84.725 26.575 85.015 26.805 ;
      RECT 83.33 26.62 85.015 26.76 ;
      RECT 80.57 24.18 80.89 24.44 ;
      RECT 83.805 24.195 84.095 24.425 ;
      RECT 80.57 24.24 84.095 24.38 ;
      RECT 83.33 17.04 83.65 17.3 ;
      RECT 82.35 17.055 82.64 17.285 ;
      RECT 82.35 17.1 83.65 17.24 ;
      RECT 83.33 21.8 83.65 22.06 ;
      RECT 80.57 21.8 80.89 22.06 ;
      RECT 80.57 21.86 83.65 22 ;
      RECT 82.415 27.255 82.705 27.485 ;
      RECT 79.895 27.255 80.185 27.485 ;
      RECT 78.705 27.255 78.995 27.485 ;
      RECT 78.705 27.3 82.705 27.44 ;
      RECT 81.98 26.915 82.27 27.145 ;
      RECT 80.41 26.915 80.7 27.145 ;
      RECT 78.31 26.915 78.6 27.145 ;
      RECT 78.31 26.96 82.27 27.1 ;
      RECT 80.57 25.54 80.89 25.8 ;
      RECT 81.965 25.555 82.255 25.785 ;
      RECT 80.57 25.6 82.255 25.74 ;
      RECT 80.57 33.7 80.89 33.96 ;
      RECT 69.53 33.7 69.85 33.96 ;
      RECT 81.965 33.715 82.255 33.945 ;
      RECT 73.3 33.76 82.255 33.9 ;
      RECT 69.53 33.76 70.68 33.9 ;
      RECT 70.54 33.42 70.68 33.9 ;
      RECT 73.3 33.42 73.44 33.9 ;
      RECT 70.54 33.42 73.44 33.56 ;
      RECT 80.57 16.7 80.89 16.96 ;
      RECT 81.045 16.715 81.335 16.945 ;
      RECT 80.57 16.76 81.335 16.9 ;
      RECT 77.81 18.4 78.13 18.66 ;
      RECT 81.045 18.415 81.335 18.645 ;
      RECT 77.81 18.46 81.335 18.6 ;
      RECT 80.57 11.6 80.89 11.86 ;
      RECT 78.36 11.66 80.89 11.8 ;
      RECT 78.36 11.275 78.5 11.8 ;
      RECT 78.285 11.275 78.575 11.505 ;
      RECT 80.57 18.74 80.89 19 ;
      RECT 75.05 18.74 75.37 19 ;
      RECT 69.53 18.74 69.85 19 ;
      RECT 73.225 18.755 73.515 18.985 ;
      RECT 69.53 18.8 80.89 18.94 ;
      RECT 80.57 24.86 80.89 25.12 ;
      RECT 77.44 24.92 80.89 25.06 ;
      RECT 77.44 24.58 77.58 25.06 ;
      RECT 76.905 24.535 77.195 24.765 ;
      RECT 76.905 24.58 77.58 24.72 ;
      RECT 80.57 27.58 80.89 27.84 ;
      RECT 79.13 27.595 79.42 27.825 ;
      RECT 79.13 27.64 80.89 27.78 ;
      RECT 79.655 32.695 79.945 32.925 ;
      RECT 77.135 32.695 77.425 32.925 ;
      RECT 75.945 32.695 76.235 32.925 ;
      RECT 75.945 32.74 79.945 32.88 ;
      RECT 79.22 32.355 79.51 32.585 ;
      RECT 77.65 32.355 77.94 32.585 ;
      RECT 75.55 32.355 75.84 32.585 ;
      RECT 75.55 32.4 79.51 32.54 ;
      RECT 78.735 19.435 79.025 19.665 ;
      RECT 76.215 19.435 76.505 19.665 ;
      RECT 75.025 19.435 75.315 19.665 ;
      RECT 75.025 19.48 79.025 19.62 ;
      RECT 78.3 19.775 78.59 20.005 ;
      RECT 76.73 19.775 77.02 20.005 ;
      RECT 74.63 19.775 74.92 20.005 ;
      RECT 74.63 19.82 78.59 19.96 ;
      RECT 77.81 24.52 78.13 24.78 ;
      RECT 77.81 24.535 78.345 24.765 ;
      RECT 77.81 25.54 78.13 25.8 ;
      RECT 75.525 25.555 75.815 25.785 ;
      RECT 75.525 25.6 78.13 25.74 ;
      RECT 77.81 33.36 78.13 33.62 ;
      RECT 76.37 33.375 76.66 33.605 ;
      RECT 76.37 33.42 78.13 33.56 ;
      RECT 75.05 27.24 75.37 27.5 ;
      RECT 77.825 27.255 78.115 27.485 ;
      RECT 75.05 27.3 78.115 27.44 ;
      RECT 72.29 24.52 72.61 24.78 ;
      RECT 72.29 24.58 72.98 24.72 ;
      RECT 72.84 24.41 72.98 24.72 ;
      RECT 72.84 24.41 75.74 24.55 ;
      RECT 75.6 24.24 75.74 24.55 ;
      RECT 77.365 24.195 77.655 24.425 ;
      RECT 75.6 24.24 77.655 24.38 ;
      RECT 67.705 20.115 67.995 20.345 ;
      RECT 67.705 20.16 74.36 20.3 ;
      RECT 74.22 19.15 74.36 20.3 ;
      RECT 75.48 19.105 75.77 19.335 ;
      RECT 74.22 19.15 75.77 19.29 ;
      RECT 75.435 24.86 75.755 25.12 ;
      RECT 69.935 24.92 75.755 25.06 ;
      RECT 69.935 24.535 70.075 25.06 ;
      RECT 69.86 24.535 70.15 24.765 ;
      RECT 69.53 15.68 69.85 15.94 ;
      RECT 73.225 15.695 73.515 15.925 ;
      RECT 69.53 15.74 73.515 15.88 ;
      RECT 72.29 19.76 72.61 20.02 ;
      RECT 71.46 19.82 72.61 19.96 ;
      RECT 66.4 19.82 67.46 19.96 ;
      RECT 67.32 19.65 67.46 19.96 ;
      RECT 71.46 19.65 71.6 19.96 ;
      RECT 66.4 19.095 66.54 19.96 ;
      RECT 67.32 19.65 71.6 19.79 ;
      RECT 66.325 19.095 66.615 19.325 ;
      RECT 65.02 21.35 71.6 21.49 ;
      RECT 71.46 21.18 71.6 21.49 ;
      RECT 72.29 21.12 72.61 21.38 ;
      RECT 64.01 21.12 64.33 21.38 ;
      RECT 65.02 21.18 65.16 21.49 ;
      RECT 71.46 21.18 72.61 21.32 ;
      RECT 64.01 21.18 65.16 21.32 ;
      RECT 72.29 26.56 72.61 26.82 ;
      RECT 61.25 26.56 61.57 26.82 ;
      RECT 70.925 26.575 71.215 26.805 ;
      RECT 61.25 26.62 72.61 26.76 ;
      RECT 70.915 16.375 71.205 16.605 ;
      RECT 68.395 16.375 68.685 16.605 ;
      RECT 67.205 16.375 67.495 16.605 ;
      RECT 67.205 16.42 71.205 16.56 ;
      RECT 70.48 16.035 70.77 16.265 ;
      RECT 68.91 16.035 69.2 16.265 ;
      RECT 66.81 16.035 67.1 16.265 ;
      RECT 66.81 16.08 70.77 16.22 ;
      RECT 69.53 11.26 69.85 11.52 ;
      RECT 69.085 11.275 69.375 11.505 ;
      RECT 69.085 11.32 69.85 11.46 ;
      RECT 69.53 16.7 69.85 16.96 ;
      RECT 66.325 16.715 66.615 16.945 ;
      RECT 66.325 16.76 69.85 16.9 ;
      RECT 69.53 27.58 69.85 27.84 ;
      RECT 64.025 27.595 64.315 27.825 ;
      RECT 51.605 27.595 51.895 27.825 ;
      RECT 51.605 27.64 69.85 27.78 ;
      RECT 69.53 29.28 69.85 29.54 ;
      RECT 66.77 29.28 67.09 29.54 ;
      RECT 66.77 29.34 69.85 29.48 ;
      RECT 69.53 38.46 69.85 38.72 ;
      RECT 66.785 38.475 67.075 38.705 ;
      RECT 66.785 38.52 69.85 38.66 ;
      RECT 52.97 24.86 53.29 25.12 ;
      RECT 60.42 24.92 68.84 25.06 ;
      RECT 68.7 24.58 68.84 25.06 ;
      RECT 52.97 24.92 54.12 25.06 ;
      RECT 53.98 24.58 54.12 25.06 ;
      RECT 60.42 24.58 60.56 25.06 ;
      RECT 69.085 24.535 69.375 24.765 ;
      RECT 68.7 24.58 69.375 24.72 ;
      RECT 53.98 24.58 60.56 24.72 ;
      RECT 68.625 24.195 68.915 24.425 ;
      RECT 62.26 24.24 68.915 24.38 ;
      RECT 62.26 23.9 62.4 24.38 ;
      RECT 61.25 23.84 61.57 24.1 ;
      RECT 61.25 23.9 62.4 24.04 ;
      RECT 68.615 27.255 68.905 27.485 ;
      RECT 66.095 27.255 66.385 27.485 ;
      RECT 64.905 27.255 65.195 27.485 ;
      RECT 64.905 27.3 68.905 27.44 ;
      RECT 68.18 26.915 68.47 27.145 ;
      RECT 66.61 26.915 66.9 27.145 ;
      RECT 64.51 26.915 64.8 27.145 ;
      RECT 64.51 26.96 68.47 27.1 ;
      RECT 64.01 22.82 64.33 23.08 ;
      RECT 68.165 22.835 68.455 23.065 ;
      RECT 64.01 22.88 68.455 23.02 ;
      RECT 66.77 24.52 67.09 24.78 ;
      RECT 67.935 24.535 68.225 24.765 ;
      RECT 66.77 24.58 68.225 24.72 ;
      RECT 66.77 17.04 67.09 17.3 ;
      RECT 67.63 17.055 67.92 17.285 ;
      RECT 66.77 17.1 67.92 17.24 ;
      RECT 52.97 25.54 53.29 25.8 ;
      RECT 67.245 25.555 67.535 25.785 ;
      RECT 65.94 25.6 67.535 25.74 ;
      RECT 52.97 25.6 55.04 25.74 ;
      RECT 54.9 25.26 55.04 25.74 ;
      RECT 65.94 25.43 66.08 25.74 ;
      RECT 59.5 25.43 66.08 25.57 ;
      RECT 59.5 25.26 59.64 25.57 ;
      RECT 54.9 25.26 59.64 25.4 ;
      RECT 66.77 19.08 67.09 19.34 ;
      RECT 66.77 19.095 67.1 19.325 ;
      RECT 66.77 13.64 67.09 13.9 ;
      RECT 66.095 13.655 66.385 13.885 ;
      RECT 66.095 13.7 67.09 13.84 ;
      RECT 58.49 22.48 58.81 22.74 ;
      RECT 66.325 22.495 66.615 22.725 ;
      RECT 58.49 22.54 66.615 22.68 ;
      RECT 65.865 19.095 66.155 19.325 ;
      RECT 65.48 19.14 66.155 19.28 ;
      RECT 65.48 18.46 65.62 19.28 ;
      RECT 58.49 18.4 58.81 18.66 ;
      RECT 58.49 18.46 65.62 18.6 ;
      RECT 65.635 22.155 65.925 22.385 ;
      RECT 65.71 21.86 65.85 22.385 ;
      RECT 58.49 21.8 58.81 22.06 ;
      RECT 55.73 21.8 56.05 22.06 ;
      RECT 47.45 21.8 47.77 22.06 ;
      RECT 47.45 21.86 65.85 22 ;
      RECT 64.01 28.26 64.33 28.52 ;
      RECT 64.01 28.32 65.545 28.46 ;
      RECT 65.405 27.935 65.545 28.46 ;
      RECT 65.33 27.935 65.62 28.165 ;
      RECT 55.73 19.76 56.05 20.02 ;
      RECT 55.73 19.82 65.165 19.96 ;
      RECT 65.025 19.105 65.165 19.96 ;
      RECT 64.95 19.105 65.24 19.335 ;
      RECT 61.25 13.3 61.57 13.56 ;
      RECT 58.49 13.3 58.81 13.56 ;
      RECT 64.945 13.315 65.235 13.545 ;
      RECT 53.905 13.315 54.195 13.545 ;
      RECT 53.905 13.36 65.235 13.5 ;
      RECT 61.25 17.38 61.57 17.64 ;
      RECT 61.25 17.44 65.16 17.58 ;
      RECT 65.02 16.715 65.16 17.58 ;
      RECT 64.945 16.715 65.235 16.945 ;
      RECT 64.01 22.14 64.33 22.4 ;
      RECT 64.945 22.155 65.235 22.385 ;
      RECT 64.01 22.2 65.235 22.34 ;
      RECT 64.485 19.095 64.775 19.325 ;
      RECT 64.56 18.8 64.7 19.325 ;
      RECT 64.01 18.74 64.33 19 ;
      RECT 64.01 18.8 64.7 18.94 ;
      RECT 63.18 14.72 64.7 14.86 ;
      RECT 64.56 14.04 64.7 14.86 ;
      RECT 53.06 14.72 56.42 14.86 ;
      RECT 56.28 14.04 56.42 14.86 ;
      RECT 63.18 14.38 63.32 14.86 ;
      RECT 53.06 14.38 53.2 14.86 ;
      RECT 58.49 14.32 58.81 14.58 ;
      RECT 47.45 14.32 47.77 14.58 ;
      RECT 56.28 14.38 63.32 14.52 ;
      RECT 46.76 14.38 53.2 14.52 ;
      RECT 46.76 13.655 46.9 14.52 ;
      RECT 64.33 14.04 64.7 14.18 ;
      RECT 55.13 14.04 56.42 14.18 ;
      RECT 64.33 13.655 64.47 14.18 ;
      RECT 55.13 13.655 55.27 14.18 ;
      RECT 64.255 13.655 64.545 13.885 ;
      RECT 55.055 13.655 55.345 13.885 ;
      RECT 46.685 13.655 46.975 13.885 ;
      RECT 64.01 14.32 64.33 14.58 ;
      RECT 63.64 14.38 64.33 14.52 ;
      RECT 63.64 13.655 63.78 14.52 ;
      RECT 57.2 13.87 62.86 14.01 ;
      RECT 62.72 13.7 62.86 14.01 ;
      RECT 55.73 13.64 56.05 13.9 ;
      RECT 63.565 13.655 63.855 13.885 ;
      RECT 57.2 13.7 57.34 14.01 ;
      RECT 62.72 13.7 63.855 13.84 ;
      RECT 55.73 13.7 57.34 13.84 ;
      RECT 58.49 11.94 58.81 12.2 ;
      RECT 59.885 11.955 60.175 12.185 ;
      RECT 58.49 12 60.175 12.14 ;
      RECT 58.49 19.08 58.81 19.34 ;
      RECT 59.425 19.095 59.715 19.325 ;
      RECT 58.49 19.14 59.715 19.28 ;
      RECT 58.49 26.56 58.81 26.82 ;
      RECT 50.21 26.56 50.53 26.82 ;
      RECT 50.21 26.62 58.81 26.76 ;
      RECT 47.45 15.68 47.77 15.94 ;
      RECT 58.505 15.695 58.795 15.925 ;
      RECT 47.45 15.74 58.795 15.88 ;
      RECT 56.195 16.375 56.485 16.605 ;
      RECT 53.675 16.375 53.965 16.605 ;
      RECT 52.485 16.375 52.775 16.605 ;
      RECT 52.485 16.42 56.485 16.56 ;
      RECT 56.195 27.255 56.485 27.485 ;
      RECT 53.675 27.255 53.965 27.485 ;
      RECT 52.485 27.255 52.775 27.485 ;
      RECT 52.485 27.3 56.485 27.44 ;
      RECT 55.73 11.94 56.05 12.2 ;
      RECT 54.9 12 56.05 12.14 ;
      RECT 54.9 11.66 55.04 12.14 ;
      RECT 47.08 11.83 52.28 11.97 ;
      RECT 52.14 11.66 52.28 11.97 ;
      RECT 37.42 11.83 42.62 11.97 ;
      RECT 42.48 11.66 42.62 11.97 ;
      RECT 44.69 11.6 45.01 11.86 ;
      RECT 35.965 11.615 36.255 11.845 ;
      RECT 47.08 11.66 47.22 11.97 ;
      RECT 37.42 11.66 37.56 11.97 ;
      RECT 52.14 11.66 55.04 11.8 ;
      RECT 42.48 11.66 47.22 11.8 ;
      RECT 35.965 11.66 37.56 11.8 ;
      RECT 55.73 14.32 56.05 14.58 ;
      RECT 54.44 14.38 56.05 14.52 ;
      RECT 54.44 13.655 54.58 14.52 ;
      RECT 50.21 13.98 50.53 14.24 ;
      RECT 50.21 14.04 54.58 14.18 ;
      RECT 54.365 13.655 54.655 13.885 ;
      RECT 55.76 16.035 56.05 16.265 ;
      RECT 54.19 16.035 54.48 16.265 ;
      RECT 52.09 16.035 52.38 16.265 ;
      RECT 52.09 16.08 56.05 16.22 ;
      RECT 55.73 18.4 56.05 18.66 ;
      RECT 53.905 18.415 54.195 18.645 ;
      RECT 53.905 18.46 56.05 18.6 ;
      RECT 55.76 26.915 56.05 27.145 ;
      RECT 54.19 26.915 54.48 27.145 ;
      RECT 52.09 26.915 52.38 27.145 ;
      RECT 52.09 26.96 56.05 27.1 ;
      RECT 52.97 13.64 53.29 13.9 ;
      RECT 52.97 13.655 53.505 13.885 ;
      RECT 48.615 13.655 48.905 13.885 ;
      RECT 52.14 13.7 53.505 13.84 ;
      RECT 48.615 13.7 49.98 13.84 ;
      RECT 49.84 13.36 49.98 13.84 ;
      RECT 52.14 13.36 52.28 13.84 ;
      RECT 49.84 13.36 52.28 13.5 ;
      RECT 52.97 9.22 53.29 9.48 ;
      RECT 39.63 9.22 39.95 9.48 ;
      RECT 52.14 9.28 53.29 9.42 ;
      RECT 39.63 9.28 40.78 9.42 ;
      RECT 40.64 8.6 40.78 9.42 ;
      RECT 52.14 8.6 52.28 9.42 ;
      RECT 40.64 8.6 52.28 8.74 ;
      RECT 52.97 27.92 53.29 28.18 ;
      RECT 52.91 27.935 53.29 28.165 ;
      RECT 50.21 17.04 50.53 17.3 ;
      RECT 52.83 17.055 53.12 17.285 ;
      RECT 50.21 17.1 53.12 17.24 ;
      RECT 50.21 14.66 50.53 14.92 ;
      RECT 52.525 14.675 52.815 14.905 ;
      RECT 50.21 14.72 52.815 14.86 ;
      RECT 47.45 16.7 47.77 16.96 ;
      RECT 51.605 16.715 51.895 16.945 ;
      RECT 47.45 16.76 51.895 16.9 ;
      RECT 51.595 19.435 51.885 19.665 ;
      RECT 49.075 19.435 49.365 19.665 ;
      RECT 47.885 19.435 48.175 19.665 ;
      RECT 47.885 19.48 51.885 19.62 ;
      RECT 51.16 19.775 51.45 20.005 ;
      RECT 49.59 19.775 49.88 20.005 ;
      RECT 47.49 19.775 47.78 20.005 ;
      RECT 47.49 19.82 51.45 19.96 ;
      RECT 50.21 25.2 50.53 25.46 ;
      RECT 44.32 25.26 50.53 25.4 ;
      RECT 49.38 24.535 49.52 25.4 ;
      RECT 44.32 24.58 44.46 25.4 ;
      RECT 49.305 24.535 49.595 24.765 ;
      RECT 40.18 24.58 44.46 24.72 ;
      RECT 40.18 24.24 40.32 24.72 ;
      RECT 36.885 24.195 37.175 24.425 ;
      RECT 36.885 24.24 40.32 24.38 ;
      RECT 44.69 14.66 45.01 14.92 ;
      RECT 49.305 14.675 49.595 14.905 ;
      RECT 44.69 14.72 49.595 14.86 ;
      RECT 48.31 18.755 48.6 18.985 ;
      RECT 48.385 18.46 48.525 18.985 ;
      RECT 44.69 18.4 45.01 18.66 ;
      RECT 44.69 18.46 48.525 18.6 ;
      RECT 47.925 13.315 48.215 13.545 ;
      RECT 48 13.02 48.14 13.545 ;
      RECT 47.45 12.96 47.77 13.22 ;
      RECT 47.45 13.02 48.14 13.16 ;
      RECT 35.045 10.935 35.335 11.165 ;
      RECT 35.12 10.47 35.26 11.165 ;
      RECT 33.65 10.58 33.97 10.84 ;
      RECT 40.18 10.64 46.76 10.78 ;
      RECT 46.62 10.3 46.76 10.78 ;
      RECT 33.65 10.64 35.26 10.78 ;
      RECT 40.18 10.47 40.32 10.78 ;
      RECT 35.12 10.47 40.32 10.61 ;
      RECT 47.45 10.24 47.77 10.5 ;
      RECT 46.62 10.3 47.77 10.44 ;
      RECT 47.45 19.08 47.77 19.34 ;
      RECT 47.005 19.095 47.295 19.325 ;
      RECT 47.005 19.14 47.77 19.28 ;
      RECT 47.45 26.56 47.77 26.82 ;
      RECT 36.41 26.56 36.73 26.82 ;
      RECT 36.41 26.62 47.77 26.76 ;
      RECT 19.85 28.26 20.17 28.52 ;
      RECT 19.85 28.32 39.86 28.46 ;
      RECT 39.72 27.98 39.86 28.46 ;
      RECT 47.45 27.92 47.77 28.18 ;
      RECT 39.72 27.98 47.77 28.12 ;
      RECT 47.465 13.655 47.755 13.885 ;
      RECT 47.54 13.36 47.68 13.885 ;
      RECT 41.93 13.3 42.25 13.56 ;
      RECT 41.93 13.36 47.68 13.5 ;
      RECT 46.085 13.655 46.375 13.885 ;
      RECT 41.56 13.7 46.375 13.84 ;
      RECT 41.56 13.02 41.7 13.84 ;
      RECT 44.69 12.96 45.01 13.22 ;
      RECT 41.56 13.02 45.01 13.16 ;
      RECT 41.1 14.38 44 14.52 ;
      RECT 43.86 14.04 44 14.52 ;
      RECT 41.1 14.04 41.24 14.52 ;
      RECT 44.69 13.98 45.01 14.24 ;
      RECT 36.41 13.98 36.73 14.24 ;
      RECT 43.86 14.04 45.01 14.18 ;
      RECT 36.41 14.04 41.24 14.18 ;
      RECT 36.96 13.655 37.1 14.18 ;
      RECT 36.885 13.655 37.175 13.885 ;
      RECT 44.69 22.82 45.01 23.08 ;
      RECT 43.785 22.835 44.075 23.065 ;
      RECT 43.785 22.88 45.01 23.02 ;
      RECT 44.69 26.9 45.01 27.16 ;
      RECT 43.785 26.915 44.075 27.145 ;
      RECT 43.785 26.96 45.01 27.1 ;
      RECT 36.885 33.035 37.175 33.265 ;
      RECT 36.96 32.4 37.1 33.265 ;
      RECT 44.69 32.34 45.01 32.6 ;
      RECT 36.96 32.4 45.01 32.54 ;
      RECT 41.93 11.26 42.25 11.52 ;
      RECT 35.505 11.275 35.795 11.505 ;
      RECT 24.925 11.275 25.215 11.505 ;
      RECT 24.925 11.32 42.25 11.46 ;
      RECT 41.93 15.68 42.25 15.94 ;
      RECT 40.105 15.695 40.395 15.925 ;
      RECT 40.105 15.74 42.25 15.88 ;
      RECT 41.93 17.38 42.25 17.64 ;
      RECT 28.13 17.38 28.45 17.64 ;
      RECT 41.1 17.44 42.25 17.58 ;
      RECT 32.36 17.44 34.8 17.58 ;
      RECT 34.66 17.27 34.8 17.58 ;
      RECT 28.13 17.44 29.28 17.58 ;
      RECT 29.14 17.1 29.28 17.58 ;
      RECT 41.1 17.1 41.24 17.58 ;
      RECT 32.36 17.1 32.5 17.58 ;
      RECT 34.66 17.27 38.94 17.41 ;
      RECT 38.8 17.1 38.94 17.41 ;
      RECT 38.8 17.1 41.24 17.24 ;
      RECT 29.14 17.1 32.5 17.24 ;
      RECT 41.93 18.4 42.25 18.66 ;
      RECT 40.565 18.415 40.855 18.645 ;
      RECT 40.565 18.46 42.25 18.6 ;
      RECT 41.93 29.62 42.25 29.88 ;
      RECT 36.885 29.635 37.175 29.865 ;
      RECT 36.885 29.68 42.25 29.82 ;
      RECT 41.93 34.72 42.25 34.98 ;
      RECT 40.105 34.735 40.395 34.965 ;
      RECT 40.105 34.78 42.25 34.92 ;
      RECT 41.475 27.255 41.765 27.485 ;
      RECT 38.955 27.255 39.245 27.485 ;
      RECT 37.765 27.255 38.055 27.485 ;
      RECT 37.765 27.3 41.765 27.44 ;
      RECT 41.04 26.915 41.33 27.145 ;
      RECT 39.47 26.915 39.76 27.145 ;
      RECT 37.37 26.915 37.66 27.145 ;
      RECT 37.37 26.96 41.33 27.1 ;
      RECT 37.575 13.655 37.865 13.885 ;
      RECT 37.65 13.02 37.79 13.885 ;
      RECT 39.17 12.96 39.49 13.22 ;
      RECT 37.65 13.02 39.49 13.16 ;
      RECT 39.17 24.52 39.49 24.78 ;
      RECT 37.575 24.535 37.865 24.765 ;
      RECT 37.575 24.58 39.49 24.72 ;
      RECT 39.17 25.54 39.49 25.8 ;
      RECT 38.265 25.555 38.555 25.785 ;
      RECT 38.265 25.6 39.49 25.74 ;
      RECT 39.17 27.92 39.49 28.18 ;
      RECT 38.19 27.935 38.48 28.165 ;
      RECT 38.19 27.98 39.49 28.12 ;
      RECT 39.17 29.96 39.49 30.22 ;
      RECT 37.575 29.975 37.865 30.205 ;
      RECT 37.575 30.02 39.49 30.16 ;
      RECT 39.17 33.02 39.49 33.28 ;
      RECT 37.575 33.035 37.865 33.265 ;
      RECT 37.575 33.08 39.49 33.22 ;
      RECT 36.41 14.66 36.73 14.92 ;
      RECT 38.265 14.675 38.555 14.905 ;
      RECT 36.41 14.72 38.555 14.86 ;
      RECT 26.38 29.68 29.28 29.82 ;
      RECT 29.14 29.34 29.28 29.82 ;
      RECT 26.38 29.34 26.52 29.82 ;
      RECT 25.37 29.28 25.69 29.54 ;
      RECT 38.265 29.295 38.555 29.525 ;
      RECT 29.14 29.34 38.555 29.48 ;
      RECT 25.37 29.34 26.52 29.48 ;
      RECT 36.41 33.7 36.73 33.96 ;
      RECT 38.265 33.715 38.555 33.945 ;
      RECT 36.41 33.76 38.555 33.9 ;
      RECT 38.255 19.435 38.545 19.665 ;
      RECT 35.735 19.435 36.025 19.665 ;
      RECT 34.545 19.435 34.835 19.665 ;
      RECT 34.545 19.48 38.545 19.62 ;
      RECT 37.82 19.775 38.11 20.005 ;
      RECT 36.25 19.775 36.54 20.005 ;
      RECT 34.15 19.775 34.44 20.005 ;
      RECT 34.15 19.82 38.11 19.96 ;
      RECT 37.795 16.375 38.085 16.605 ;
      RECT 35.275 16.375 35.565 16.605 ;
      RECT 34.085 16.375 34.375 16.605 ;
      RECT 34.085 16.42 38.085 16.56 ;
      RECT 37.795 35.755 38.085 35.985 ;
      RECT 35.275 35.755 35.565 35.985 ;
      RECT 34.085 35.755 34.375 35.985 ;
      RECT 34.085 35.8 38.085 35.94 ;
      RECT 37.36 16.035 37.65 16.265 ;
      RECT 35.79 16.035 36.08 16.265 ;
      RECT 33.69 16.035 33.98 16.265 ;
      RECT 33.69 16.08 37.65 16.22 ;
      RECT 37.36 36.095 37.65 36.325 ;
      RECT 35.79 36.095 36.08 36.325 ;
      RECT 33.69 36.095 33.98 36.325 ;
      RECT 33.69 36.14 37.65 36.28 ;
      RECT 33.65 27.58 33.97 27.84 ;
      RECT 36.885 27.595 37.175 27.825 ;
      RECT 22.165 27.595 22.455 27.825 ;
      RECT 22.165 27.64 37.175 27.78 ;
      RECT 36.41 11.94 36.73 12.2 ;
      RECT 33.665 11.955 33.955 12.185 ;
      RECT 33.665 12 36.73 12.14 ;
      RECT 36.41 16.7 36.73 16.96 ;
      RECT 34.51 16.715 34.8 16.945 ;
      RECT 34.51 16.76 36.73 16.9 ;
      RECT 36.41 18.74 36.73 19 ;
      RECT 34.97 18.755 35.26 18.985 ;
      RECT 34.97 18.8 36.73 18.94 ;
      RECT 36.41 22.82 36.73 23.08 ;
      RECT 36.5 22.2 36.64 23.08 ;
      RECT 35.045 22.155 35.335 22.385 ;
      RECT 35.045 22.2 36.64 22.34 ;
      RECT 36.41 24.86 36.73 25.12 ;
      RECT 36.5 24.58 36.64 25.12 ;
      RECT 35.735 24.535 36.025 24.765 ;
      RECT 35.735 24.58 36.64 24.72 ;
      RECT 36.41 30.98 36.73 31.24 ;
      RECT 35.81 31.04 36.73 31.18 ;
      RECT 35.81 29.975 35.95 31.18 ;
      RECT 35.735 29.975 36.025 30.205 ;
      RECT 35.735 33.035 36.025 33.265 ;
      RECT 35.81 32.06 35.95 33.265 ;
      RECT 36.41 32 36.73 32.26 ;
      RECT 35.81 32.06 36.73 32.2 ;
      RECT 36.41 35.06 36.73 35.32 ;
      RECT 34.51 35.075 34.8 35.305 ;
      RECT 34.51 35.12 36.73 35.26 ;
      RECT 36.425 13.315 36.715 13.545 ;
      RECT 35.12 13.36 36.715 13.5 ;
      RECT 35.12 13.19 35.26 13.5 ;
      RECT 29.14 13.19 35.26 13.33 ;
      RECT 28.13 12.96 28.45 13.22 ;
      RECT 29.14 13.02 29.28 13.33 ;
      RECT 28.13 13.02 29.28 13.16 ;
      RECT 25 30.36 30.2 30.5 ;
      RECT 30.06 29.68 30.2 30.5 ;
      RECT 25 30.02 25.14 30.5 ;
      RECT 20.86 30.02 25.14 30.16 ;
      RECT 20.86 29.68 21 30.16 ;
      RECT 19.85 29.62 20.17 29.88 ;
      RECT 36.425 29.635 36.715 29.865 ;
      RECT 30.06 29.68 36.715 29.82 ;
      RECT 19.85 29.68 21 29.82 ;
      RECT 33.65 13.98 33.97 14.24 ;
      RECT 33.65 14.04 35.95 14.18 ;
      RECT 35.81 13.655 35.95 14.18 ;
      RECT 35.735 13.655 36.025 13.885 ;
      RECT 30.89 13.64 31.21 13.9 ;
      RECT 35.045 13.655 35.335 13.885 ;
      RECT 30.89 13.7 35.335 13.84 ;
      RECT 30.89 24.52 31.21 24.78 ;
      RECT 35.045 24.535 35.335 24.765 ;
      RECT 30.89 24.58 35.335 24.72 ;
      RECT 31.9 30.36 34.34 30.5 ;
      RECT 34.2 30.02 34.34 30.5 ;
      RECT 31.9 30.02 32.04 30.5 ;
      RECT 30.89 29.96 31.21 30.22 ;
      RECT 35.045 29.975 35.335 30.205 ;
      RECT 34.2 30.02 35.335 30.16 ;
      RECT 30.89 30.02 32.04 30.16 ;
      RECT 35.045 33.035 35.335 33.265 ;
      RECT 35.12 32.74 35.26 33.265 ;
      RECT 30.89 32.68 31.21 32.94 ;
      RECT 30.89 32.74 35.26 32.88 ;
      RECT 30.89 10.24 31.21 10.5 ;
      RECT 34.585 10.255 34.875 10.485 ;
      RECT 30.89 10.3 34.875 10.44 ;
      RECT 33.65 16.7 33.97 16.96 ;
      RECT 33.205 16.715 33.495 16.945 ;
      RECT 33.205 16.76 33.97 16.9 ;
      RECT 33.65 35.4 33.97 35.66 ;
      RECT 33.205 35.415 33.495 35.645 ;
      RECT 33.205 35.46 33.97 35.6 ;
      RECT 28.13 26.56 28.45 26.82 ;
      RECT 29.065 26.575 29.355 26.805 ;
      RECT 28.13 26.62 29.355 26.76 ;
      RECT 28.13 11.94 28.45 12.2 ;
      RECT 27.3 12 28.45 12.14 ;
      RECT 16.72 12 18.7 12.14 ;
      RECT 18.56 11.32 18.7 12.14 ;
      RECT 27.3 11.83 27.44 12.14 ;
      RECT 16.72 11.275 16.86 12.14 ;
      RECT 24.08 11.83 27.44 11.97 ;
      RECT 24.08 11.32 24.22 11.97 ;
      RECT 16.645 11.275 16.935 11.505 ;
      RECT 18.56 11.32 24.22 11.46 ;
      RECT 28.13 19.08 28.45 19.34 ;
      RECT 21.245 19.095 21.535 19.325 ;
      RECT 21.245 19.14 28.45 19.28 ;
      RECT 26.755 27.255 27.045 27.485 ;
      RECT 24.235 27.255 24.525 27.485 ;
      RECT 23.045 27.255 23.335 27.485 ;
      RECT 23.045 27.3 27.045 27.44 ;
      RECT 26.32 26.915 26.61 27.145 ;
      RECT 24.75 26.915 25.04 27.145 ;
      RECT 22.65 26.915 22.94 27.145 ;
      RECT 22.65 26.96 26.61 27.1 ;
      RECT 25.37 27.92 25.69 28.18 ;
      RECT 23.47 27.935 23.76 28.165 ;
      RECT 23.47 27.98 25.69 28.12 ;
      RECT 19.85 22.14 20.17 22.4 ;
      RECT 18.485 22.155 18.775 22.385 ;
      RECT 18.485 22.2 20.17 22.34 ;
      RECT 10.12 9.62 189.98 10.1 ;
      RECT 10.12 12.34 189.98 12.82 ;
      RECT 10.12 15.06 189.98 15.54 ;
      RECT 10.12 17.78 189.98 18.26 ;
      RECT 10.12 20.5 189.98 20.98 ;
      RECT 10.12 23.22 189.98 23.7 ;
      RECT 10.12 25.94 189.98 26.42 ;
      RECT 10.12 28.66 189.98 29.14 ;
      RECT 10.12 31.38 189.98 31.86 ;
      RECT 10.12 34.1 189.98 34.58 ;
      RECT 10.12 36.82 189.98 37.3 ;
      RECT 10.12 39.54 189.98 40.02 ;
      RECT 10.12 42.26 189.98 42.74 ;
      RECT 10.12 44.98 189.98 45.46 ;
      RECT 10.12 47.7 189.98 48.18 ;
      RECT 10.12 50.42 189.98 50.9 ;
      RECT 10.12 53.14 189.98 53.62 ;
      RECT 10.12 55.86 189.98 56.34 ;
      RECT 10.12 58.58 189.98 59.06 ;
      RECT 177.17 11.26 177.49 11.52 ;
      RECT 171.65 14.66 171.97 14.92 ;
      RECT 171.65 19.08 171.97 19.34 ;
      RECT 168.89 11.26 169.21 11.52 ;
      RECT 149.57 19.08 149.89 19.34 ;
      RECT 144.05 24.52 144.37 24.78 ;
      RECT 138.53 27.24 138.85 27.5 ;
      RECT 135.77 24.52 136.09 24.78 ;
      RECT 133.01 11.26 133.33 11.52 ;
      RECT 133.01 16.7 133.33 16.96 ;
      RECT 130.25 22.14 130.57 22.4 ;
      RECT 130.25 27.24 130.57 27.825 ;
      RECT 124.73 11.26 125.05 11.52 ;
      RECT 124.73 20.1 125.05 20.36 ;
      RECT 121.97 14.66 122.29 14.92 ;
      RECT 119.21 11.26 119.53 11.52 ;
      RECT 119.21 18.4 119.53 18.66 ;
      RECT 108.17 29.62 108.86 29.88 ;
      RECT 97.13 11.26 97.45 11.52 ;
      RECT 91.61 11.26 91.93 11.52 ;
      RECT 83.33 11.26 83.65 11.52 ;
      RECT 83.33 19.76 83.65 20.02 ;
      RECT 83.33 24.52 83.65 24.78 ;
      RECT 75.05 32.68 75.37 32.94 ;
      RECT 72.29 19.08 72.61 19.34 ;
      RECT 66.77 14.66 67.09 14.92 ;
      RECT 66.77 22.48 67.09 22.74 ;
      RECT 61.25 19.08 61.57 19.34 ;
      RECT 58.49 17.38 58.81 17.64 ;
      RECT 47.45 11.26 47.77 11.52 ;
      RECT 36.41 10.92 36.73 11.18 ;
      RECT 36.41 24.18 36.73 24.44 ;
      RECT 33.65 19.08 33.97 19.34 ;
    LAYER via ;
      RECT 189.215 12.505 189.365 12.655 ;
      RECT 189.215 17.945 189.365 18.095 ;
      RECT 189.215 23.385 189.365 23.535 ;
      RECT 189.215 28.825 189.365 28.975 ;
      RECT 189.215 34.265 189.365 34.415 ;
      RECT 189.215 39.705 189.365 39.855 ;
      RECT 189.215 45.145 189.365 45.295 ;
      RECT 189.215 50.585 189.365 50.735 ;
      RECT 189.215 56.025 189.365 56.175 ;
      RECT 187.375 9.895 187.525 10.045 ;
      RECT 187.375 15.225 187.525 15.375 ;
      RECT 187.375 20.665 187.525 20.815 ;
      RECT 187.375 26.105 187.525 26.255 ;
      RECT 187.375 31.545 187.525 31.695 ;
      RECT 187.375 36.985 187.525 37.135 ;
      RECT 187.375 42.425 187.525 42.575 ;
      RECT 187.375 47.865 187.525 48.015 ;
      RECT 187.375 53.305 187.525 53.455 ;
      RECT 187.375 58.745 187.525 58.895 ;
      RECT 186.455 12.505 186.605 12.655 ;
      RECT 186.455 17.945 186.605 18.095 ;
      RECT 186.455 23.385 186.605 23.535 ;
      RECT 186.455 28.825 186.605 28.975 ;
      RECT 186.455 34.265 186.605 34.415 ;
      RECT 186.455 39.705 186.605 39.855 ;
      RECT 186.455 45.145 186.605 45.295 ;
      RECT 186.455 50.585 186.605 50.735 ;
      RECT 186.455 56.025 186.605 56.175 ;
      RECT 184.615 9.895 184.765 10.045 ;
      RECT 184.615 15.225 184.765 15.375 ;
      RECT 184.615 20.665 184.765 20.815 ;
      RECT 184.615 26.105 184.765 26.255 ;
      RECT 184.615 31.545 184.765 31.695 ;
      RECT 184.615 36.985 184.765 37.135 ;
      RECT 184.615 42.425 184.765 42.575 ;
      RECT 184.615 47.865 184.765 48.015 ;
      RECT 184.615 53.305 184.765 53.455 ;
      RECT 184.615 58.745 184.765 58.895 ;
      RECT 183.695 12.505 183.845 12.655 ;
      RECT 183.695 17.945 183.845 18.095 ;
      RECT 183.695 23.385 183.845 23.535 ;
      RECT 183.695 28.825 183.845 28.975 ;
      RECT 183.695 34.265 183.845 34.415 ;
      RECT 183.695 39.705 183.845 39.855 ;
      RECT 183.695 45.145 183.845 45.295 ;
      RECT 183.695 50.585 183.845 50.735 ;
      RECT 183.695 56.025 183.845 56.175 ;
      RECT 181.855 9.895 182.005 10.045 ;
      RECT 181.855 15.225 182.005 15.375 ;
      RECT 181.855 20.665 182.005 20.815 ;
      RECT 181.855 26.105 182.005 26.255 ;
      RECT 181.855 31.545 182.005 31.695 ;
      RECT 181.855 36.985 182.005 37.135 ;
      RECT 181.855 42.425 182.005 42.575 ;
      RECT 181.855 47.865 182.005 48.015 ;
      RECT 181.855 53.305 182.005 53.455 ;
      RECT 181.855 58.745 182.005 58.895 ;
      RECT 180.935 12.505 181.085 12.655 ;
      RECT 180.935 17.945 181.085 18.095 ;
      RECT 180.935 23.385 181.085 23.535 ;
      RECT 180.935 28.825 181.085 28.975 ;
      RECT 180.935 34.265 181.085 34.415 ;
      RECT 180.935 39.705 181.085 39.855 ;
      RECT 180.935 45.145 181.085 45.295 ;
      RECT 180.935 50.585 181.085 50.735 ;
      RECT 180.935 56.025 181.085 56.175 ;
      RECT 180.015 11.995 180.165 12.145 ;
      RECT 180.015 16.755 180.165 16.905 ;
      RECT 179.095 9.895 179.245 10.045 ;
      RECT 179.095 15.225 179.245 15.375 ;
      RECT 179.095 20.665 179.245 20.815 ;
      RECT 179.095 26.105 179.245 26.255 ;
      RECT 179.095 31.545 179.245 31.695 ;
      RECT 179.095 36.985 179.245 37.135 ;
      RECT 179.095 42.425 179.245 42.575 ;
      RECT 179.095 47.865 179.245 48.015 ;
      RECT 179.095 53.305 179.245 53.455 ;
      RECT 179.095 58.745 179.245 58.895 ;
      RECT 178.175 12.505 178.325 12.655 ;
      RECT 178.175 17.945 178.325 18.095 ;
      RECT 178.175 23.385 178.325 23.535 ;
      RECT 178.175 28.825 178.325 28.975 ;
      RECT 178.175 34.265 178.325 34.415 ;
      RECT 178.175 39.705 178.325 39.855 ;
      RECT 178.175 45.145 178.325 45.295 ;
      RECT 178.175 50.585 178.325 50.735 ;
      RECT 178.175 56.025 178.325 56.175 ;
      RECT 177.255 11.315 177.405 11.465 ;
      RECT 177.255 15.735 177.405 15.885 ;
      RECT 177.255 17.435 177.405 17.585 ;
      RECT 177.255 19.475 177.405 19.625 ;
      RECT 176.335 9.895 176.485 10.045 ;
      RECT 176.335 15.225 176.485 15.375 ;
      RECT 176.335 20.665 176.485 20.815 ;
      RECT 176.335 26.105 176.485 26.255 ;
      RECT 176.335 31.545 176.485 31.695 ;
      RECT 176.335 36.985 176.485 37.135 ;
      RECT 176.335 42.425 176.485 42.575 ;
      RECT 176.335 47.865 176.485 48.015 ;
      RECT 176.335 53.305 176.485 53.455 ;
      RECT 176.335 58.745 176.485 58.895 ;
      RECT 175.415 12.505 175.565 12.655 ;
      RECT 175.415 17.945 175.565 18.095 ;
      RECT 175.415 23.385 175.565 23.535 ;
      RECT 175.415 28.825 175.565 28.975 ;
      RECT 175.415 34.265 175.565 34.415 ;
      RECT 175.415 39.705 175.565 39.855 ;
      RECT 175.415 45.145 175.565 45.295 ;
      RECT 175.415 50.585 175.565 50.735 ;
      RECT 175.415 56.025 175.565 56.175 ;
      RECT 173.575 9.895 173.725 10.045 ;
      RECT 173.575 15.225 173.725 15.375 ;
      RECT 173.575 20.665 173.725 20.815 ;
      RECT 173.575 26.105 173.725 26.255 ;
      RECT 173.575 31.545 173.725 31.695 ;
      RECT 173.575 36.985 173.725 37.135 ;
      RECT 173.575 42.425 173.725 42.575 ;
      RECT 173.575 47.865 173.725 48.015 ;
      RECT 173.575 53.305 173.725 53.455 ;
      RECT 173.575 58.745 173.725 58.895 ;
      RECT 172.655 12.505 172.805 12.655 ;
      RECT 172.655 17.945 172.805 18.095 ;
      RECT 172.655 23.385 172.805 23.535 ;
      RECT 172.655 28.825 172.805 28.975 ;
      RECT 172.655 34.265 172.805 34.415 ;
      RECT 172.655 39.705 172.805 39.855 ;
      RECT 172.655 45.145 172.805 45.295 ;
      RECT 172.655 50.585 172.805 50.735 ;
      RECT 172.655 56.025 172.805 56.175 ;
      RECT 171.735 14.715 171.885 14.865 ;
      RECT 171.735 17.435 171.885 17.585 ;
      RECT 171.735 18.455 171.885 18.605 ;
      RECT 171.735 19.135 171.885 19.285 ;
      RECT 171.735 20.155 171.885 20.305 ;
      RECT 170.815 9.895 170.965 10.045 ;
      RECT 170.815 15.225 170.965 15.375 ;
      RECT 170.815 20.665 170.965 20.815 ;
      RECT 170.815 26.105 170.965 26.255 ;
      RECT 170.815 31.545 170.965 31.695 ;
      RECT 170.815 36.985 170.965 37.135 ;
      RECT 170.815 42.425 170.965 42.575 ;
      RECT 170.815 47.865 170.965 48.015 ;
      RECT 170.815 53.305 170.965 53.455 ;
      RECT 170.815 58.745 170.965 58.895 ;
      RECT 169.895 12.505 170.045 12.655 ;
      RECT 169.895 17.945 170.045 18.095 ;
      RECT 169.895 23.385 170.045 23.535 ;
      RECT 169.895 28.825 170.045 28.975 ;
      RECT 169.895 34.265 170.045 34.415 ;
      RECT 169.895 39.705 170.045 39.855 ;
      RECT 169.895 45.145 170.045 45.295 ;
      RECT 169.895 50.585 170.045 50.735 ;
      RECT 169.895 56.025 170.045 56.175 ;
      RECT 168.975 11.315 169.125 11.465 ;
      RECT 168.975 15.735 169.125 15.885 ;
      RECT 168.975 18.455 169.125 18.605 ;
      RECT 168.975 22.195 169.125 22.345 ;
      RECT 168.975 26.955 169.125 27.105 ;
      RECT 168.055 9.895 168.205 10.045 ;
      RECT 168.055 15.225 168.205 15.375 ;
      RECT 168.055 20.665 168.205 20.815 ;
      RECT 168.055 26.105 168.205 26.255 ;
      RECT 168.055 31.545 168.205 31.695 ;
      RECT 168.055 36.985 168.205 37.135 ;
      RECT 168.055 42.425 168.205 42.575 ;
      RECT 168.055 47.865 168.205 48.015 ;
      RECT 168.055 53.305 168.205 53.455 ;
      RECT 168.055 58.745 168.205 58.895 ;
      RECT 167.135 12.505 167.285 12.655 ;
      RECT 167.135 17.945 167.285 18.095 ;
      RECT 167.135 23.385 167.285 23.535 ;
      RECT 167.135 28.825 167.285 28.975 ;
      RECT 167.135 34.265 167.285 34.415 ;
      RECT 167.135 39.705 167.285 39.855 ;
      RECT 167.135 45.145 167.285 45.295 ;
      RECT 167.135 50.585 167.285 50.735 ;
      RECT 167.135 56.025 167.285 56.175 ;
      RECT 165.295 9.895 165.445 10.045 ;
      RECT 165.295 15.225 165.445 15.375 ;
      RECT 165.295 20.665 165.445 20.815 ;
      RECT 165.295 26.105 165.445 26.255 ;
      RECT 165.295 31.545 165.445 31.695 ;
      RECT 165.295 36.985 165.445 37.135 ;
      RECT 165.295 42.425 165.445 42.575 ;
      RECT 165.295 47.865 165.445 48.015 ;
      RECT 165.295 53.305 165.445 53.455 ;
      RECT 165.295 58.745 165.445 58.895 ;
      RECT 164.375 12.505 164.525 12.655 ;
      RECT 164.375 17.945 164.525 18.095 ;
      RECT 164.375 23.385 164.525 23.535 ;
      RECT 164.375 28.825 164.525 28.975 ;
      RECT 164.375 34.265 164.525 34.415 ;
      RECT 164.375 39.705 164.525 39.855 ;
      RECT 164.375 45.145 164.525 45.295 ;
      RECT 164.375 50.585 164.525 50.735 ;
      RECT 164.375 56.025 164.525 56.175 ;
      RECT 163.455 14.375 163.605 14.525 ;
      RECT 163.455 15.735 163.605 15.885 ;
      RECT 163.455 23.895 163.605 24.045 ;
      RECT 162.535 9.895 162.685 10.045 ;
      RECT 162.535 15.225 162.685 15.375 ;
      RECT 162.535 20.665 162.685 20.815 ;
      RECT 162.535 26.105 162.685 26.255 ;
      RECT 162.535 31.545 162.685 31.695 ;
      RECT 162.535 36.985 162.685 37.135 ;
      RECT 162.535 42.425 162.685 42.575 ;
      RECT 162.535 47.865 162.685 48.015 ;
      RECT 162.535 53.305 162.685 53.455 ;
      RECT 162.535 58.745 162.685 58.895 ;
      RECT 161.615 12.505 161.765 12.655 ;
      RECT 161.615 17.945 161.765 18.095 ;
      RECT 161.615 23.385 161.765 23.535 ;
      RECT 161.615 28.825 161.765 28.975 ;
      RECT 161.615 34.265 161.765 34.415 ;
      RECT 161.615 39.705 161.765 39.855 ;
      RECT 161.615 45.145 161.765 45.295 ;
      RECT 161.615 50.585 161.765 50.735 ;
      RECT 161.615 56.025 161.765 56.175 ;
      RECT 160.695 16.755 160.845 16.905 ;
      RECT 160.695 19.475 160.845 19.625 ;
      RECT 160.695 30.015 160.845 30.165 ;
      RECT 160.695 33.415 160.845 33.565 ;
      RECT 159.775 9.895 159.925 10.045 ;
      RECT 159.775 15.225 159.925 15.375 ;
      RECT 159.775 20.665 159.925 20.815 ;
      RECT 159.775 26.105 159.925 26.255 ;
      RECT 159.775 31.545 159.925 31.695 ;
      RECT 159.775 36.985 159.925 37.135 ;
      RECT 159.775 42.425 159.925 42.575 ;
      RECT 159.775 47.865 159.925 48.015 ;
      RECT 159.775 53.305 159.925 53.455 ;
      RECT 159.775 58.745 159.925 58.895 ;
      RECT 158.855 12.505 159.005 12.655 ;
      RECT 158.855 17.945 159.005 18.095 ;
      RECT 158.855 23.385 159.005 23.535 ;
      RECT 158.855 28.825 159.005 28.975 ;
      RECT 158.855 34.265 159.005 34.415 ;
      RECT 158.855 39.705 159.005 39.855 ;
      RECT 158.855 45.145 159.005 45.295 ;
      RECT 158.855 50.585 159.005 50.735 ;
      RECT 158.855 56.025 159.005 56.175 ;
      RECT 157.935 17.435 158.085 17.585 ;
      RECT 157.935 18.455 158.085 18.605 ;
      RECT 157.935 19.135 158.085 19.285 ;
      RECT 157.935 25.255 158.085 25.405 ;
      RECT 157.935 27.295 158.085 27.445 ;
      RECT 157.935 27.975 158.085 28.125 ;
      RECT 157.935 32.735 158.085 32.885 ;
      RECT 157.935 34.775 158.085 34.925 ;
      RECT 157.015 9.895 157.165 10.045 ;
      RECT 157.015 15.225 157.165 15.375 ;
      RECT 157.015 20.665 157.165 20.815 ;
      RECT 157.015 26.105 157.165 26.255 ;
      RECT 157.015 31.545 157.165 31.695 ;
      RECT 157.015 36.985 157.165 37.135 ;
      RECT 157.015 42.425 157.165 42.575 ;
      RECT 157.015 47.865 157.165 48.015 ;
      RECT 157.015 53.305 157.165 53.455 ;
      RECT 157.015 58.745 157.165 58.895 ;
      RECT 156.095 12.505 156.245 12.655 ;
      RECT 156.095 17.945 156.245 18.095 ;
      RECT 156.095 23.385 156.245 23.535 ;
      RECT 156.095 28.825 156.245 28.975 ;
      RECT 156.095 34.265 156.245 34.415 ;
      RECT 156.095 39.705 156.245 39.855 ;
      RECT 156.095 45.145 156.245 45.295 ;
      RECT 156.095 50.585 156.245 50.735 ;
      RECT 156.095 56.025 156.245 56.175 ;
      RECT 155.175 11.315 155.325 11.465 ;
      RECT 155.175 24.575 155.325 24.725 ;
      RECT 155.175 29.335 155.325 29.485 ;
      RECT 155.175 32.395 155.325 32.545 ;
      RECT 155.175 33.755 155.325 33.905 ;
      RECT 155.175 35.115 155.325 35.265 ;
      RECT 154.255 9.895 154.405 10.045 ;
      RECT 154.255 15.225 154.405 15.375 ;
      RECT 154.255 20.665 154.405 20.815 ;
      RECT 154.255 26.105 154.405 26.255 ;
      RECT 154.255 31.545 154.405 31.695 ;
      RECT 154.255 36.985 154.405 37.135 ;
      RECT 154.255 42.425 154.405 42.575 ;
      RECT 154.255 47.865 154.405 48.015 ;
      RECT 154.255 53.305 154.405 53.455 ;
      RECT 154.255 58.745 154.405 58.895 ;
      RECT 153.335 12.505 153.485 12.655 ;
      RECT 153.335 17.945 153.485 18.095 ;
      RECT 153.335 23.385 153.485 23.535 ;
      RECT 153.335 28.825 153.485 28.975 ;
      RECT 153.335 34.265 153.485 34.415 ;
      RECT 153.335 39.705 153.485 39.855 ;
      RECT 153.335 45.145 153.485 45.295 ;
      RECT 153.335 50.585 153.485 50.735 ;
      RECT 153.335 56.025 153.485 56.175 ;
      RECT 152.415 11.315 152.565 11.465 ;
      RECT 152.415 13.015 152.565 13.165 ;
      RECT 152.415 15.735 152.565 15.885 ;
      RECT 152.415 18.455 152.565 18.605 ;
      RECT 152.415 19.135 152.565 19.285 ;
      RECT 152.415 19.815 152.565 19.965 ;
      RECT 152.415 23.895 152.565 24.045 ;
      RECT 152.415 26.615 152.565 26.765 ;
      RECT 152.415 27.635 152.565 27.785 ;
      RECT 152.415 28.315 152.565 28.465 ;
      RECT 152.415 29.675 152.565 29.825 ;
      RECT 152.415 32.055 152.565 32.205 ;
      RECT 152.415 33.075 152.565 33.225 ;
      RECT 151.495 9.895 151.645 10.045 ;
      RECT 151.495 15.225 151.645 15.375 ;
      RECT 151.495 20.665 151.645 20.815 ;
      RECT 151.495 26.105 151.645 26.255 ;
      RECT 151.495 31.545 151.645 31.695 ;
      RECT 151.495 36.985 151.645 37.135 ;
      RECT 151.495 42.425 151.645 42.575 ;
      RECT 151.495 47.865 151.645 48.015 ;
      RECT 151.495 53.305 151.645 53.455 ;
      RECT 151.495 58.745 151.645 58.895 ;
      RECT 150.575 12.505 150.725 12.655 ;
      RECT 150.575 17.945 150.725 18.095 ;
      RECT 150.575 23.385 150.725 23.535 ;
      RECT 150.575 28.825 150.725 28.975 ;
      RECT 150.575 34.265 150.725 34.415 ;
      RECT 150.575 39.705 150.725 39.855 ;
      RECT 150.575 45.145 150.725 45.295 ;
      RECT 150.575 50.585 150.725 50.735 ;
      RECT 150.575 56.025 150.725 56.175 ;
      RECT 149.655 17.095 149.805 17.245 ;
      RECT 149.655 18.455 149.805 18.605 ;
      RECT 149.655 19.135 149.805 19.285 ;
      RECT 149.655 19.815 149.805 19.965 ;
      RECT 149.655 21.515 149.805 21.665 ;
      RECT 149.655 22.875 149.805 23.025 ;
      RECT 149.655 25.255 149.805 25.405 ;
      RECT 148.735 9.895 148.885 10.045 ;
      RECT 148.735 15.225 148.885 15.375 ;
      RECT 148.735 20.665 148.885 20.815 ;
      RECT 148.735 26.105 148.885 26.255 ;
      RECT 148.735 31.545 148.885 31.695 ;
      RECT 148.735 36.985 148.885 37.135 ;
      RECT 148.735 42.425 148.885 42.575 ;
      RECT 148.735 47.865 148.885 48.015 ;
      RECT 148.735 53.305 148.885 53.455 ;
      RECT 148.735 58.745 148.885 58.895 ;
      RECT 147.815 12.505 147.965 12.655 ;
      RECT 147.815 17.945 147.965 18.095 ;
      RECT 147.815 23.385 147.965 23.535 ;
      RECT 147.815 28.825 147.965 28.975 ;
      RECT 147.815 34.265 147.965 34.415 ;
      RECT 147.815 39.705 147.965 39.855 ;
      RECT 147.815 45.145 147.965 45.295 ;
      RECT 147.815 50.585 147.965 50.735 ;
      RECT 147.815 56.025 147.965 56.175 ;
      RECT 146.895 14.375 147.045 14.525 ;
      RECT 146.895 18.455 147.045 18.605 ;
      RECT 146.895 19.135 147.045 19.285 ;
      RECT 146.895 21.175 147.045 21.325 ;
      RECT 146.895 21.855 147.045 22.005 ;
      RECT 146.895 24.915 147.045 25.065 ;
      RECT 146.895 25.595 147.045 25.745 ;
      RECT 146.895 26.615 147.045 26.765 ;
      RECT 145.975 9.895 146.125 10.045 ;
      RECT 145.975 15.225 146.125 15.375 ;
      RECT 145.975 20.665 146.125 20.815 ;
      RECT 145.975 26.105 146.125 26.255 ;
      RECT 145.975 31.545 146.125 31.695 ;
      RECT 145.975 36.985 146.125 37.135 ;
      RECT 145.975 42.425 146.125 42.575 ;
      RECT 145.975 47.865 146.125 48.015 ;
      RECT 145.975 53.305 146.125 53.455 ;
      RECT 145.975 58.745 146.125 58.895 ;
      RECT 145.055 12.505 145.205 12.655 ;
      RECT 145.055 17.945 145.205 18.095 ;
      RECT 145.055 23.385 145.205 23.535 ;
      RECT 145.055 28.825 145.205 28.975 ;
      RECT 145.055 34.265 145.205 34.415 ;
      RECT 145.055 39.705 145.205 39.855 ;
      RECT 145.055 45.145 145.205 45.295 ;
      RECT 145.055 50.585 145.205 50.735 ;
      RECT 145.055 56.025 145.205 56.175 ;
      RECT 144.135 22.875 144.285 23.025 ;
      RECT 144.135 24.575 144.285 24.725 ;
      RECT 144.135 26.615 144.285 26.765 ;
      RECT 143.215 9.895 143.365 10.045 ;
      RECT 143.215 15.225 143.365 15.375 ;
      RECT 143.215 20.665 143.365 20.815 ;
      RECT 143.215 26.105 143.365 26.255 ;
      RECT 143.215 31.545 143.365 31.695 ;
      RECT 143.215 36.985 143.365 37.135 ;
      RECT 143.215 42.425 143.365 42.575 ;
      RECT 143.215 47.865 143.365 48.015 ;
      RECT 143.215 53.305 143.365 53.455 ;
      RECT 143.215 58.745 143.365 58.895 ;
      RECT 142.295 12.505 142.445 12.655 ;
      RECT 142.295 17.945 142.445 18.095 ;
      RECT 142.295 23.385 142.445 23.535 ;
      RECT 142.295 28.825 142.445 28.975 ;
      RECT 142.295 34.265 142.445 34.415 ;
      RECT 142.295 39.705 142.445 39.855 ;
      RECT 142.295 45.145 142.445 45.295 ;
      RECT 142.295 50.585 142.445 50.735 ;
      RECT 142.295 56.025 142.445 56.175 ;
      RECT 141.375 17.435 141.525 17.585 ;
      RECT 141.375 18.455 141.525 18.605 ;
      RECT 141.375 21.855 141.525 22.005 ;
      RECT 141.375 24.575 141.525 24.725 ;
      RECT 141.375 25.595 141.525 25.745 ;
      RECT 141.375 27.975 141.525 28.125 ;
      RECT 140.455 9.895 140.605 10.045 ;
      RECT 140.455 15.225 140.605 15.375 ;
      RECT 140.455 20.665 140.605 20.815 ;
      RECT 140.455 26.105 140.605 26.255 ;
      RECT 140.455 31.545 140.605 31.695 ;
      RECT 140.455 36.985 140.605 37.135 ;
      RECT 140.455 42.425 140.605 42.575 ;
      RECT 140.455 47.865 140.605 48.015 ;
      RECT 140.455 53.305 140.605 53.455 ;
      RECT 140.455 58.745 140.605 58.895 ;
      RECT 139.535 12.505 139.685 12.655 ;
      RECT 139.535 17.945 139.685 18.095 ;
      RECT 139.535 23.385 139.685 23.535 ;
      RECT 139.535 28.825 139.685 28.975 ;
      RECT 139.535 34.265 139.685 34.415 ;
      RECT 139.535 39.705 139.685 39.855 ;
      RECT 139.535 45.145 139.685 45.295 ;
      RECT 139.535 50.585 139.685 50.735 ;
      RECT 139.535 56.025 139.685 56.175 ;
      RECT 138.615 14.715 138.765 14.865 ;
      RECT 138.615 15.735 138.765 15.885 ;
      RECT 138.615 19.135 138.765 19.285 ;
      RECT 138.615 27.295 138.765 27.445 ;
      RECT 138.615 30.015 138.765 30.165 ;
      RECT 137.695 9.895 137.845 10.045 ;
      RECT 137.695 15.225 137.845 15.375 ;
      RECT 137.695 20.665 137.845 20.815 ;
      RECT 137.695 26.105 137.845 26.255 ;
      RECT 137.695 31.545 137.845 31.695 ;
      RECT 137.695 36.985 137.845 37.135 ;
      RECT 137.695 42.425 137.845 42.575 ;
      RECT 137.695 47.865 137.845 48.015 ;
      RECT 137.695 53.305 137.845 53.455 ;
      RECT 137.695 58.745 137.845 58.895 ;
      RECT 136.775 12.505 136.925 12.655 ;
      RECT 136.775 17.945 136.925 18.095 ;
      RECT 136.775 23.385 136.925 23.535 ;
      RECT 136.775 28.825 136.925 28.975 ;
      RECT 136.775 34.265 136.925 34.415 ;
      RECT 136.775 39.705 136.925 39.855 ;
      RECT 136.775 45.145 136.925 45.295 ;
      RECT 136.775 50.585 136.925 50.735 ;
      RECT 136.775 56.025 136.925 56.175 ;
      RECT 135.855 13.015 136.005 13.165 ;
      RECT 135.855 16.755 136.005 16.905 ;
      RECT 135.855 21.515 136.005 21.665 ;
      RECT 135.855 22.875 136.005 23.025 ;
      RECT 135.855 24.575 136.005 24.725 ;
      RECT 135.855 25.595 136.005 25.745 ;
      RECT 135.855 26.955 136.005 27.105 ;
      RECT 135.855 27.975 136.005 28.125 ;
      RECT 135.855 34.775 136.005 34.925 ;
      RECT 134.935 9.895 135.085 10.045 ;
      RECT 134.935 15.225 135.085 15.375 ;
      RECT 134.935 20.665 135.085 20.815 ;
      RECT 134.935 26.105 135.085 26.255 ;
      RECT 134.935 31.545 135.085 31.695 ;
      RECT 134.935 36.985 135.085 37.135 ;
      RECT 134.935 42.425 135.085 42.575 ;
      RECT 134.935 47.865 135.085 48.015 ;
      RECT 134.935 53.305 135.085 53.455 ;
      RECT 134.935 58.745 135.085 58.895 ;
      RECT 134.015 12.505 134.165 12.655 ;
      RECT 134.015 17.945 134.165 18.095 ;
      RECT 134.015 23.385 134.165 23.535 ;
      RECT 134.015 28.825 134.165 28.975 ;
      RECT 134.015 34.265 134.165 34.415 ;
      RECT 134.015 39.705 134.165 39.855 ;
      RECT 134.015 45.145 134.165 45.295 ;
      RECT 134.015 50.585 134.165 50.735 ;
      RECT 134.015 56.025 134.165 56.175 ;
      RECT 133.095 11.315 133.245 11.465 ;
      RECT 133.095 14.375 133.245 14.525 ;
      RECT 133.095 16.755 133.245 16.905 ;
      RECT 133.095 21.175 133.245 21.325 ;
      RECT 133.095 22.195 133.245 22.345 ;
      RECT 133.095 22.875 133.245 23.025 ;
      RECT 133.095 24.915 133.245 25.065 ;
      RECT 133.095 25.595 133.245 25.745 ;
      RECT 133.095 26.955 133.245 27.105 ;
      RECT 132.175 9.895 132.325 10.045 ;
      RECT 132.175 15.225 132.325 15.375 ;
      RECT 132.175 20.665 132.325 20.815 ;
      RECT 132.175 26.105 132.325 26.255 ;
      RECT 132.175 31.545 132.325 31.695 ;
      RECT 132.175 36.985 132.325 37.135 ;
      RECT 132.175 42.425 132.325 42.575 ;
      RECT 132.175 47.865 132.325 48.015 ;
      RECT 132.175 53.305 132.325 53.455 ;
      RECT 132.175 58.745 132.325 58.895 ;
      RECT 131.255 12.505 131.405 12.655 ;
      RECT 131.255 17.945 131.405 18.095 ;
      RECT 131.255 23.385 131.405 23.535 ;
      RECT 131.255 28.825 131.405 28.975 ;
      RECT 131.255 34.265 131.405 34.415 ;
      RECT 131.255 39.705 131.405 39.855 ;
      RECT 131.255 45.145 131.405 45.295 ;
      RECT 131.255 50.585 131.405 50.735 ;
      RECT 131.255 56.025 131.405 56.175 ;
      RECT 130.335 14.375 130.485 14.525 ;
      RECT 130.335 19.135 130.485 19.285 ;
      RECT 130.335 20.155 130.485 20.305 ;
      RECT 130.335 22.195 130.485 22.345 ;
      RECT 130.335 23.895 130.485 24.045 ;
      RECT 130.335 24.915 130.485 25.065 ;
      RECT 130.335 26.615 130.485 26.765 ;
      RECT 130.335 27.295 130.485 27.445 ;
      RECT 130.335 28.315 130.485 28.465 ;
      RECT 130.335 29.335 130.485 29.485 ;
      RECT 130.335 33.415 130.485 33.565 ;
      RECT 130.335 34.775 130.485 34.925 ;
      RECT 129.415 9.895 129.565 10.045 ;
      RECT 129.415 15.225 129.565 15.375 ;
      RECT 129.415 20.665 129.565 20.815 ;
      RECT 129.415 26.105 129.565 26.255 ;
      RECT 129.415 31.545 129.565 31.695 ;
      RECT 129.415 36.985 129.565 37.135 ;
      RECT 129.415 42.425 129.565 42.575 ;
      RECT 129.415 47.865 129.565 48.015 ;
      RECT 129.415 53.305 129.565 53.455 ;
      RECT 129.415 58.745 129.565 58.895 ;
      RECT 128.495 12.505 128.645 12.655 ;
      RECT 128.495 17.945 128.645 18.095 ;
      RECT 128.495 23.385 128.645 23.535 ;
      RECT 128.495 28.825 128.645 28.975 ;
      RECT 128.495 34.265 128.645 34.415 ;
      RECT 128.495 39.705 128.645 39.855 ;
      RECT 128.495 45.145 128.645 45.295 ;
      RECT 128.495 50.585 128.645 50.735 ;
      RECT 128.495 56.025 128.645 56.175 ;
      RECT 127.575 21.175 127.725 21.325 ;
      RECT 127.575 22.195 127.725 22.345 ;
      RECT 127.575 24.575 127.725 24.725 ;
      RECT 127.575 25.595 127.725 25.745 ;
      RECT 127.575 27.635 127.725 27.785 ;
      RECT 127.575 29.335 127.725 29.485 ;
      RECT 127.575 34.775 127.725 34.925 ;
      RECT 126.655 9.895 126.805 10.045 ;
      RECT 126.655 15.225 126.805 15.375 ;
      RECT 126.655 20.665 126.805 20.815 ;
      RECT 126.655 26.105 126.805 26.255 ;
      RECT 126.655 31.545 126.805 31.695 ;
      RECT 126.655 36.985 126.805 37.135 ;
      RECT 126.655 42.425 126.805 42.575 ;
      RECT 126.655 47.865 126.805 48.015 ;
      RECT 126.655 53.305 126.805 53.455 ;
      RECT 126.655 58.745 126.805 58.895 ;
      RECT 125.735 12.505 125.885 12.655 ;
      RECT 125.735 17.945 125.885 18.095 ;
      RECT 125.735 23.385 125.885 23.535 ;
      RECT 125.735 28.825 125.885 28.975 ;
      RECT 125.735 34.265 125.885 34.415 ;
      RECT 125.735 39.705 125.885 39.855 ;
      RECT 125.735 45.145 125.885 45.295 ;
      RECT 125.735 50.585 125.885 50.735 ;
      RECT 125.735 56.025 125.885 56.175 ;
      RECT 124.815 11.315 124.965 11.465 ;
      RECT 124.815 15.735 124.965 15.885 ;
      RECT 124.815 20.155 124.965 20.305 ;
      RECT 124.815 22.195 124.965 22.345 ;
      RECT 124.815 35.455 124.965 35.605 ;
      RECT 123.895 9.895 124.045 10.045 ;
      RECT 123.895 15.225 124.045 15.375 ;
      RECT 123.895 20.665 124.045 20.815 ;
      RECT 123.895 26.105 124.045 26.255 ;
      RECT 123.895 31.545 124.045 31.695 ;
      RECT 123.895 36.985 124.045 37.135 ;
      RECT 123.895 42.425 124.045 42.575 ;
      RECT 123.895 47.865 124.045 48.015 ;
      RECT 123.895 53.305 124.045 53.455 ;
      RECT 123.895 58.745 124.045 58.895 ;
      RECT 122.975 12.505 123.125 12.655 ;
      RECT 122.975 17.945 123.125 18.095 ;
      RECT 122.975 23.385 123.125 23.535 ;
      RECT 122.975 28.825 123.125 28.975 ;
      RECT 122.975 34.265 123.125 34.415 ;
      RECT 122.975 39.705 123.125 39.855 ;
      RECT 122.975 45.145 123.125 45.295 ;
      RECT 122.975 50.585 123.125 50.735 ;
      RECT 122.975 56.025 123.125 56.175 ;
      RECT 122.055 14.715 122.205 14.865 ;
      RECT 122.055 19.135 122.205 19.285 ;
      RECT 122.055 26.955 122.205 27.105 ;
      RECT 121.135 9.895 121.285 10.045 ;
      RECT 121.135 15.225 121.285 15.375 ;
      RECT 121.135 20.665 121.285 20.815 ;
      RECT 121.135 26.105 121.285 26.255 ;
      RECT 121.135 31.545 121.285 31.695 ;
      RECT 121.135 36.985 121.285 37.135 ;
      RECT 121.135 42.425 121.285 42.575 ;
      RECT 121.135 47.865 121.285 48.015 ;
      RECT 121.135 53.305 121.285 53.455 ;
      RECT 121.135 58.745 121.285 58.895 ;
      RECT 120.215 12.505 120.365 12.655 ;
      RECT 120.215 17.945 120.365 18.095 ;
      RECT 120.215 23.385 120.365 23.535 ;
      RECT 120.215 28.825 120.365 28.975 ;
      RECT 120.215 34.265 120.365 34.415 ;
      RECT 120.215 39.705 120.365 39.855 ;
      RECT 120.215 45.145 120.365 45.295 ;
      RECT 120.215 50.585 120.365 50.735 ;
      RECT 120.215 56.025 120.365 56.175 ;
      RECT 119.295 11.315 119.445 11.465 ;
      RECT 119.295 14.715 119.445 14.865 ;
      RECT 119.295 15.735 119.445 15.885 ;
      RECT 119.295 17.095 119.445 17.245 ;
      RECT 119.295 18.455 119.445 18.605 ;
      RECT 119.295 21.855 119.445 22.005 ;
      RECT 119.295 22.535 119.445 22.685 ;
      RECT 119.295 25.595 119.445 25.745 ;
      RECT 119.295 26.615 119.445 26.765 ;
      RECT 118.375 9.895 118.525 10.045 ;
      RECT 118.375 15.225 118.525 15.375 ;
      RECT 118.375 20.665 118.525 20.815 ;
      RECT 118.375 26.105 118.525 26.255 ;
      RECT 118.375 31.545 118.525 31.695 ;
      RECT 118.375 36.985 118.525 37.135 ;
      RECT 118.375 42.425 118.525 42.575 ;
      RECT 118.375 47.865 118.525 48.015 ;
      RECT 118.375 53.305 118.525 53.455 ;
      RECT 118.375 58.745 118.525 58.895 ;
      RECT 117.455 12.505 117.605 12.655 ;
      RECT 117.455 17.945 117.605 18.095 ;
      RECT 117.455 23.385 117.605 23.535 ;
      RECT 117.455 28.825 117.605 28.975 ;
      RECT 117.455 34.265 117.605 34.415 ;
      RECT 117.455 39.705 117.605 39.855 ;
      RECT 117.455 45.145 117.605 45.295 ;
      RECT 117.455 50.585 117.605 50.735 ;
      RECT 117.455 56.025 117.605 56.175 ;
      RECT 116.535 11.315 116.685 11.465 ;
      RECT 116.535 13.015 116.685 13.165 ;
      RECT 116.535 16.755 116.685 16.905 ;
      RECT 116.535 17.435 116.685 17.585 ;
      RECT 116.535 19.135 116.685 19.285 ;
      RECT 116.535 20.155 116.685 20.305 ;
      RECT 116.535 22.195 116.685 22.345 ;
      RECT 116.535 22.875 116.685 23.025 ;
      RECT 116.535 27.635 116.685 27.785 ;
      RECT 115.615 9.895 115.765 10.045 ;
      RECT 115.615 15.225 115.765 15.375 ;
      RECT 115.615 20.665 115.765 20.815 ;
      RECT 115.615 26.105 115.765 26.255 ;
      RECT 115.615 31.545 115.765 31.695 ;
      RECT 115.615 36.985 115.765 37.135 ;
      RECT 115.615 42.425 115.765 42.575 ;
      RECT 115.615 47.865 115.765 48.015 ;
      RECT 115.615 53.305 115.765 53.455 ;
      RECT 115.615 58.745 115.765 58.895 ;
      RECT 114.695 12.505 114.845 12.655 ;
      RECT 114.695 17.945 114.845 18.095 ;
      RECT 114.695 23.385 114.845 23.535 ;
      RECT 114.695 28.825 114.845 28.975 ;
      RECT 114.695 34.265 114.845 34.415 ;
      RECT 114.695 39.705 114.845 39.855 ;
      RECT 114.695 45.145 114.845 45.295 ;
      RECT 114.695 50.585 114.845 50.735 ;
      RECT 114.695 56.025 114.845 56.175 ;
      RECT 113.775 13.695 113.925 13.845 ;
      RECT 113.775 17.435 113.925 17.585 ;
      RECT 113.775 18.455 113.925 18.605 ;
      RECT 113.775 22.195 113.925 22.345 ;
      RECT 113.775 25.255 113.925 25.405 ;
      RECT 113.775 26.615 113.925 26.765 ;
      RECT 112.855 9.895 113.005 10.045 ;
      RECT 112.855 15.225 113.005 15.375 ;
      RECT 112.855 20.665 113.005 20.815 ;
      RECT 112.855 26.105 113.005 26.255 ;
      RECT 112.855 31.545 113.005 31.695 ;
      RECT 112.855 36.985 113.005 37.135 ;
      RECT 112.855 42.425 113.005 42.575 ;
      RECT 112.855 47.865 113.005 48.015 ;
      RECT 112.855 53.305 113.005 53.455 ;
      RECT 112.855 58.745 113.005 58.895 ;
      RECT 111.935 12.505 112.085 12.655 ;
      RECT 111.935 17.945 112.085 18.095 ;
      RECT 111.935 23.385 112.085 23.535 ;
      RECT 111.935 28.825 112.085 28.975 ;
      RECT 111.935 34.265 112.085 34.415 ;
      RECT 111.935 39.705 112.085 39.855 ;
      RECT 111.935 45.145 112.085 45.295 ;
      RECT 111.935 50.585 112.085 50.735 ;
      RECT 111.935 56.025 112.085 56.175 ;
      RECT 111.4 22.195 111.55 22.345 ;
      RECT 111.015 13.355 111.165 13.505 ;
      RECT 111.015 16.415 111.165 16.565 ;
      RECT 111.015 18.795 111.165 18.945 ;
      RECT 111.015 27.635 111.165 27.785 ;
      RECT 111.015 30.015 111.165 30.165 ;
      RECT 110.095 9.895 110.245 10.045 ;
      RECT 110.095 15.225 110.245 15.375 ;
      RECT 110.095 20.665 110.245 20.815 ;
      RECT 110.095 26.105 110.245 26.255 ;
      RECT 110.095 31.545 110.245 31.695 ;
      RECT 110.095 36.985 110.245 37.135 ;
      RECT 110.095 42.425 110.245 42.575 ;
      RECT 110.095 47.865 110.245 48.015 ;
      RECT 110.095 53.305 110.245 53.455 ;
      RECT 110.095 58.745 110.245 58.895 ;
      RECT 109.175 12.505 109.325 12.655 ;
      RECT 109.175 17.945 109.325 18.095 ;
      RECT 109.175 23.385 109.325 23.535 ;
      RECT 109.175 28.825 109.325 28.975 ;
      RECT 109.175 34.265 109.325 34.415 ;
      RECT 109.175 39.705 109.325 39.855 ;
      RECT 109.175 45.145 109.325 45.295 ;
      RECT 109.175 50.585 109.325 50.735 ;
      RECT 109.175 56.025 109.325 56.175 ;
      RECT 108.255 14.375 108.405 14.525 ;
      RECT 108.255 17.435 108.405 17.585 ;
      RECT 108.255 18.455 108.405 18.605 ;
      RECT 108.255 22.195 108.405 22.345 ;
      RECT 108.255 22.875 108.405 23.025 ;
      RECT 108.255 29.675 108.405 29.825 ;
      RECT 107.335 9.895 107.485 10.045 ;
      RECT 107.335 15.225 107.485 15.375 ;
      RECT 107.335 20.665 107.485 20.815 ;
      RECT 107.335 26.105 107.485 26.255 ;
      RECT 107.335 31.545 107.485 31.695 ;
      RECT 107.335 36.985 107.485 37.135 ;
      RECT 107.335 42.425 107.485 42.575 ;
      RECT 107.335 47.865 107.485 48.015 ;
      RECT 107.335 53.305 107.485 53.455 ;
      RECT 107.335 58.745 107.485 58.895 ;
      RECT 106.415 12.505 106.565 12.655 ;
      RECT 106.415 17.945 106.565 18.095 ;
      RECT 106.415 23.385 106.565 23.535 ;
      RECT 106.415 28.825 106.565 28.975 ;
      RECT 106.415 34.265 106.565 34.415 ;
      RECT 106.415 39.705 106.565 39.855 ;
      RECT 106.415 45.145 106.565 45.295 ;
      RECT 106.415 50.585 106.565 50.735 ;
      RECT 106.415 56.025 106.565 56.175 ;
      RECT 105.495 13.695 105.645 13.845 ;
      RECT 105.495 14.375 105.645 14.525 ;
      RECT 105.495 19.135 105.645 19.285 ;
      RECT 105.495 19.815 105.645 19.965 ;
      RECT 105.495 21.175 105.645 21.325 ;
      RECT 105.495 25.595 105.645 25.745 ;
      RECT 104.575 9.895 104.725 10.045 ;
      RECT 104.575 15.225 104.725 15.375 ;
      RECT 104.575 20.665 104.725 20.815 ;
      RECT 104.575 26.105 104.725 26.255 ;
      RECT 104.575 31.545 104.725 31.695 ;
      RECT 104.575 36.985 104.725 37.135 ;
      RECT 104.575 42.425 104.725 42.575 ;
      RECT 104.575 47.865 104.725 48.015 ;
      RECT 104.575 53.305 104.725 53.455 ;
      RECT 104.575 58.745 104.725 58.895 ;
      RECT 103.655 12.505 103.805 12.655 ;
      RECT 103.655 17.945 103.805 18.095 ;
      RECT 103.655 23.385 103.805 23.535 ;
      RECT 103.655 28.825 103.805 28.975 ;
      RECT 103.655 34.265 103.805 34.415 ;
      RECT 103.655 39.705 103.805 39.855 ;
      RECT 103.655 45.145 103.805 45.295 ;
      RECT 103.655 50.585 103.805 50.735 ;
      RECT 103.655 56.025 103.805 56.175 ;
      RECT 102.735 16.755 102.885 16.905 ;
      RECT 102.735 22.195 102.885 22.345 ;
      RECT 102.735 24.235 102.885 24.385 ;
      RECT 102.735 28.315 102.885 28.465 ;
      RECT 102.735 34.775 102.885 34.925 ;
      RECT 101.815 9.895 101.965 10.045 ;
      RECT 101.815 15.225 101.965 15.375 ;
      RECT 101.815 20.665 101.965 20.815 ;
      RECT 101.815 26.105 101.965 26.255 ;
      RECT 101.815 31.545 101.965 31.695 ;
      RECT 101.815 36.985 101.965 37.135 ;
      RECT 101.815 42.425 101.965 42.575 ;
      RECT 101.815 47.865 101.965 48.015 ;
      RECT 101.815 53.305 101.965 53.455 ;
      RECT 101.815 58.745 101.965 58.895 ;
      RECT 100.895 12.505 101.045 12.655 ;
      RECT 100.895 17.945 101.045 18.095 ;
      RECT 100.895 23.385 101.045 23.535 ;
      RECT 100.895 28.825 101.045 28.975 ;
      RECT 100.895 34.265 101.045 34.415 ;
      RECT 100.895 39.705 101.045 39.855 ;
      RECT 100.895 45.145 101.045 45.295 ;
      RECT 100.895 50.585 101.045 50.735 ;
      RECT 100.895 56.025 101.045 56.175 ;
      RECT 99.975 11.655 100.125 11.805 ;
      RECT 99.975 13.695 100.125 13.845 ;
      RECT 99.975 17.435 100.125 17.585 ;
      RECT 99.975 18.795 100.125 18.945 ;
      RECT 99.975 24.915 100.125 25.065 ;
      RECT 99.975 29.335 100.125 29.485 ;
      RECT 99.975 32.735 100.125 32.885 ;
      RECT 99.055 9.895 99.205 10.045 ;
      RECT 99.055 15.225 99.205 15.375 ;
      RECT 99.055 20.665 99.205 20.815 ;
      RECT 99.055 26.105 99.205 26.255 ;
      RECT 99.055 31.545 99.205 31.695 ;
      RECT 99.055 36.985 99.205 37.135 ;
      RECT 99.055 42.425 99.205 42.575 ;
      RECT 99.055 47.865 99.205 48.015 ;
      RECT 99.055 53.305 99.205 53.455 ;
      RECT 99.055 58.745 99.205 58.895 ;
      RECT 98.135 12.505 98.285 12.655 ;
      RECT 98.135 17.945 98.285 18.095 ;
      RECT 98.135 23.385 98.285 23.535 ;
      RECT 98.135 28.825 98.285 28.975 ;
      RECT 98.135 34.265 98.285 34.415 ;
      RECT 98.135 39.705 98.285 39.855 ;
      RECT 98.135 45.145 98.285 45.295 ;
      RECT 98.135 50.585 98.285 50.735 ;
      RECT 98.135 56.025 98.285 56.175 ;
      RECT 97.215 11.315 97.365 11.465 ;
      RECT 97.215 15.735 97.365 15.885 ;
      RECT 97.215 16.755 97.365 16.905 ;
      RECT 97.215 18.455 97.365 18.605 ;
      RECT 97.215 19.815 97.365 19.965 ;
      RECT 97.215 21.175 97.365 21.325 ;
      RECT 97.215 22.195 97.365 22.345 ;
      RECT 97.215 23.895 97.365 24.045 ;
      RECT 97.215 24.575 97.365 24.725 ;
      RECT 97.215 33.075 97.365 33.225 ;
      RECT 97.215 33.755 97.365 33.905 ;
      RECT 97.215 35.115 97.365 35.265 ;
      RECT 96.295 9.895 96.445 10.045 ;
      RECT 96.295 15.225 96.445 15.375 ;
      RECT 96.295 20.665 96.445 20.815 ;
      RECT 96.295 26.105 96.445 26.255 ;
      RECT 96.295 31.545 96.445 31.695 ;
      RECT 96.295 36.985 96.445 37.135 ;
      RECT 96.295 42.425 96.445 42.575 ;
      RECT 96.295 47.865 96.445 48.015 ;
      RECT 96.295 53.305 96.445 53.455 ;
      RECT 96.295 58.745 96.445 58.895 ;
      RECT 95.375 12.505 95.525 12.655 ;
      RECT 95.375 17.945 95.525 18.095 ;
      RECT 95.375 23.385 95.525 23.535 ;
      RECT 95.375 28.825 95.525 28.975 ;
      RECT 95.375 34.265 95.525 34.415 ;
      RECT 95.375 39.705 95.525 39.855 ;
      RECT 95.375 45.145 95.525 45.295 ;
      RECT 95.375 50.585 95.525 50.735 ;
      RECT 95.375 56.025 95.525 56.175 ;
      RECT 94.455 16.755 94.605 16.905 ;
      RECT 94.455 22.535 94.605 22.685 ;
      RECT 93.535 9.895 93.685 10.045 ;
      RECT 93.535 15.225 93.685 15.375 ;
      RECT 93.535 20.665 93.685 20.815 ;
      RECT 93.535 26.105 93.685 26.255 ;
      RECT 93.535 31.545 93.685 31.695 ;
      RECT 93.535 36.985 93.685 37.135 ;
      RECT 93.535 42.425 93.685 42.575 ;
      RECT 93.535 47.865 93.685 48.015 ;
      RECT 93.535 53.305 93.685 53.455 ;
      RECT 93.535 58.745 93.685 58.895 ;
      RECT 92.615 12.505 92.765 12.655 ;
      RECT 92.615 17.945 92.765 18.095 ;
      RECT 92.615 23.385 92.765 23.535 ;
      RECT 92.615 28.825 92.765 28.975 ;
      RECT 92.615 34.265 92.765 34.415 ;
      RECT 92.615 39.705 92.765 39.855 ;
      RECT 92.615 45.145 92.765 45.295 ;
      RECT 92.615 50.585 92.765 50.735 ;
      RECT 92.615 56.025 92.765 56.175 ;
      RECT 91.695 11.315 91.845 11.465 ;
      RECT 91.695 20.155 91.845 20.305 ;
      RECT 91.695 21.515 91.845 21.665 ;
      RECT 91.695 25.595 91.845 25.745 ;
      RECT 91.695 35.455 91.845 35.605 ;
      RECT 90.775 9.895 90.925 10.045 ;
      RECT 90.775 15.225 90.925 15.375 ;
      RECT 90.775 20.665 90.925 20.815 ;
      RECT 90.775 26.105 90.925 26.255 ;
      RECT 90.775 31.545 90.925 31.695 ;
      RECT 90.775 36.985 90.925 37.135 ;
      RECT 90.775 42.425 90.925 42.575 ;
      RECT 90.775 47.865 90.925 48.015 ;
      RECT 90.775 53.305 90.925 53.455 ;
      RECT 90.775 58.745 90.925 58.895 ;
      RECT 89.855 12.505 90.005 12.655 ;
      RECT 89.855 17.945 90.005 18.095 ;
      RECT 89.855 23.385 90.005 23.535 ;
      RECT 89.855 28.825 90.005 28.975 ;
      RECT 89.855 34.265 90.005 34.415 ;
      RECT 89.855 39.705 90.005 39.855 ;
      RECT 89.855 45.145 90.005 45.295 ;
      RECT 89.855 50.585 90.005 50.735 ;
      RECT 89.855 56.025 90.005 56.175 ;
      RECT 88.935 15.735 89.085 15.885 ;
      RECT 88.935 19.135 89.085 19.285 ;
      RECT 88.935 19.815 89.085 19.965 ;
      RECT 88.935 22.535 89.085 22.685 ;
      RECT 88.935 24.915 89.085 25.065 ;
      RECT 88.935 26.615 89.085 26.765 ;
      RECT 88.935 32.055 89.085 32.205 ;
      RECT 88.015 9.895 88.165 10.045 ;
      RECT 88.015 15.225 88.165 15.375 ;
      RECT 88.015 20.665 88.165 20.815 ;
      RECT 88.015 26.105 88.165 26.255 ;
      RECT 88.015 31.545 88.165 31.695 ;
      RECT 88.015 36.985 88.165 37.135 ;
      RECT 88.015 42.425 88.165 42.575 ;
      RECT 88.015 47.865 88.165 48.015 ;
      RECT 88.015 53.305 88.165 53.455 ;
      RECT 88.015 58.745 88.165 58.895 ;
      RECT 87.095 12.505 87.245 12.655 ;
      RECT 87.095 17.945 87.245 18.095 ;
      RECT 87.095 23.385 87.245 23.535 ;
      RECT 87.095 28.825 87.245 28.975 ;
      RECT 87.095 34.265 87.245 34.415 ;
      RECT 87.095 39.705 87.245 39.855 ;
      RECT 87.095 45.145 87.245 45.295 ;
      RECT 87.095 50.585 87.245 50.735 ;
      RECT 87.095 56.025 87.245 56.175 ;
      RECT 86.175 17.435 86.325 17.585 ;
      RECT 86.175 18.455 86.325 18.605 ;
      RECT 86.175 19.135 86.325 19.285 ;
      RECT 86.175 25.255 86.325 25.405 ;
      RECT 86.175 32.055 86.325 32.205 ;
      RECT 86.175 33.075 86.325 33.225 ;
      RECT 85.255 9.895 85.405 10.045 ;
      RECT 85.255 15.225 85.405 15.375 ;
      RECT 85.255 20.665 85.405 20.815 ;
      RECT 85.255 26.105 85.405 26.255 ;
      RECT 85.255 31.545 85.405 31.695 ;
      RECT 85.255 36.985 85.405 37.135 ;
      RECT 85.255 42.425 85.405 42.575 ;
      RECT 85.255 47.865 85.405 48.015 ;
      RECT 85.255 53.305 85.405 53.455 ;
      RECT 85.255 58.745 85.405 58.895 ;
      RECT 84.335 12.505 84.485 12.655 ;
      RECT 84.335 17.945 84.485 18.095 ;
      RECT 84.335 23.385 84.485 23.535 ;
      RECT 84.335 28.825 84.485 28.975 ;
      RECT 84.335 34.265 84.485 34.415 ;
      RECT 84.335 39.705 84.485 39.855 ;
      RECT 84.335 45.145 84.485 45.295 ;
      RECT 84.335 50.585 84.485 50.735 ;
      RECT 84.335 56.025 84.485 56.175 ;
      RECT 83.415 11.315 83.565 11.465 ;
      RECT 83.415 14.035 83.565 14.185 ;
      RECT 83.415 17.095 83.565 17.245 ;
      RECT 83.415 19.815 83.565 19.965 ;
      RECT 83.415 21.855 83.565 22.005 ;
      RECT 83.415 22.535 83.565 22.685 ;
      RECT 83.415 24.575 83.565 24.725 ;
      RECT 83.415 26.615 83.565 26.765 ;
      RECT 82.495 9.895 82.645 10.045 ;
      RECT 82.495 15.225 82.645 15.375 ;
      RECT 82.495 20.665 82.645 20.815 ;
      RECT 82.495 26.105 82.645 26.255 ;
      RECT 82.495 31.545 82.645 31.695 ;
      RECT 82.495 36.985 82.645 37.135 ;
      RECT 82.495 42.425 82.645 42.575 ;
      RECT 82.495 47.865 82.645 48.015 ;
      RECT 82.495 53.305 82.645 53.455 ;
      RECT 82.495 58.745 82.645 58.895 ;
      RECT 81.575 12.505 81.725 12.655 ;
      RECT 81.575 17.945 81.725 18.095 ;
      RECT 81.575 23.385 81.725 23.535 ;
      RECT 81.575 28.825 81.725 28.975 ;
      RECT 81.575 34.265 81.725 34.415 ;
      RECT 81.575 39.705 81.725 39.855 ;
      RECT 81.575 45.145 81.725 45.295 ;
      RECT 81.575 50.585 81.725 50.735 ;
      RECT 81.575 56.025 81.725 56.175 ;
      RECT 80.655 11.655 80.805 11.805 ;
      RECT 80.655 16.755 80.805 16.905 ;
      RECT 80.655 18.795 80.805 18.945 ;
      RECT 80.655 19.815 80.805 19.965 ;
      RECT 80.655 21.855 80.805 22.005 ;
      RECT 80.655 24.235 80.805 24.385 ;
      RECT 80.655 24.915 80.805 25.065 ;
      RECT 80.655 25.595 80.805 25.745 ;
      RECT 80.655 27.635 80.805 27.785 ;
      RECT 80.655 33.755 80.805 33.905 ;
      RECT 79.735 9.895 79.885 10.045 ;
      RECT 79.735 15.225 79.885 15.375 ;
      RECT 79.735 20.665 79.885 20.815 ;
      RECT 79.735 26.105 79.885 26.255 ;
      RECT 79.735 31.545 79.885 31.695 ;
      RECT 79.735 36.985 79.885 37.135 ;
      RECT 79.735 42.425 79.885 42.575 ;
      RECT 79.735 47.865 79.885 48.015 ;
      RECT 79.735 53.305 79.885 53.455 ;
      RECT 79.735 58.745 79.885 58.895 ;
      RECT 78.815 12.505 78.965 12.655 ;
      RECT 78.815 17.945 78.965 18.095 ;
      RECT 78.815 23.385 78.965 23.535 ;
      RECT 78.815 28.825 78.965 28.975 ;
      RECT 78.815 34.265 78.965 34.415 ;
      RECT 78.815 39.705 78.965 39.855 ;
      RECT 78.815 45.145 78.965 45.295 ;
      RECT 78.815 50.585 78.965 50.735 ;
      RECT 78.815 56.025 78.965 56.175 ;
      RECT 77.895 18.455 78.045 18.605 ;
      RECT 77.895 24.575 78.045 24.725 ;
      RECT 77.895 25.595 78.045 25.745 ;
      RECT 77.895 33.415 78.045 33.565 ;
      RECT 76.975 9.895 77.125 10.045 ;
      RECT 76.975 15.225 77.125 15.375 ;
      RECT 76.975 20.665 77.125 20.815 ;
      RECT 76.975 26.105 77.125 26.255 ;
      RECT 76.975 31.545 77.125 31.695 ;
      RECT 76.975 36.985 77.125 37.135 ;
      RECT 76.975 42.425 77.125 42.575 ;
      RECT 76.975 47.865 77.125 48.015 ;
      RECT 76.975 53.305 77.125 53.455 ;
      RECT 76.975 58.745 77.125 58.895 ;
      RECT 76.055 12.505 76.205 12.655 ;
      RECT 76.055 17.945 76.205 18.095 ;
      RECT 76.055 23.385 76.205 23.535 ;
      RECT 76.055 28.825 76.205 28.975 ;
      RECT 76.055 34.265 76.205 34.415 ;
      RECT 76.055 39.705 76.205 39.855 ;
      RECT 76.055 45.145 76.205 45.295 ;
      RECT 76.055 50.585 76.205 50.735 ;
      RECT 76.055 56.025 76.205 56.175 ;
      RECT 75.52 24.915 75.67 25.065 ;
      RECT 75.135 16.755 75.285 16.905 ;
      RECT 75.135 18.795 75.285 18.945 ;
      RECT 75.135 27.295 75.285 27.445 ;
      RECT 75.135 32.735 75.285 32.885 ;
      RECT 74.215 9.895 74.365 10.045 ;
      RECT 74.215 15.225 74.365 15.375 ;
      RECT 74.215 20.665 74.365 20.815 ;
      RECT 74.215 26.105 74.365 26.255 ;
      RECT 74.215 31.545 74.365 31.695 ;
      RECT 74.215 36.985 74.365 37.135 ;
      RECT 74.215 42.425 74.365 42.575 ;
      RECT 74.215 47.865 74.365 48.015 ;
      RECT 74.215 53.305 74.365 53.455 ;
      RECT 74.215 58.745 74.365 58.895 ;
      RECT 73.295 12.505 73.445 12.655 ;
      RECT 73.295 17.945 73.445 18.095 ;
      RECT 73.295 23.385 73.445 23.535 ;
      RECT 73.295 28.825 73.445 28.975 ;
      RECT 73.295 34.265 73.445 34.415 ;
      RECT 73.295 39.705 73.445 39.855 ;
      RECT 73.295 45.145 73.445 45.295 ;
      RECT 73.295 50.585 73.445 50.735 ;
      RECT 73.295 56.025 73.445 56.175 ;
      RECT 72.375 19.135 72.525 19.285 ;
      RECT 72.375 19.815 72.525 19.965 ;
      RECT 72.375 21.175 72.525 21.325 ;
      RECT 72.375 23.895 72.525 24.045 ;
      RECT 72.375 24.575 72.525 24.725 ;
      RECT 72.375 26.615 72.525 26.765 ;
      RECT 71.455 9.895 71.605 10.045 ;
      RECT 71.455 15.225 71.605 15.375 ;
      RECT 71.455 20.665 71.605 20.815 ;
      RECT 71.455 26.105 71.605 26.255 ;
      RECT 71.455 31.545 71.605 31.695 ;
      RECT 71.455 36.985 71.605 37.135 ;
      RECT 71.455 42.425 71.605 42.575 ;
      RECT 71.455 47.865 71.605 48.015 ;
      RECT 71.455 53.305 71.605 53.455 ;
      RECT 71.455 58.745 71.605 58.895 ;
      RECT 70.535 12.505 70.685 12.655 ;
      RECT 70.535 17.945 70.685 18.095 ;
      RECT 70.535 23.385 70.685 23.535 ;
      RECT 70.535 28.825 70.685 28.975 ;
      RECT 70.535 34.265 70.685 34.415 ;
      RECT 70.535 39.705 70.685 39.855 ;
      RECT 70.535 45.145 70.685 45.295 ;
      RECT 70.535 50.585 70.685 50.735 ;
      RECT 70.535 56.025 70.685 56.175 ;
      RECT 69.615 11.315 69.765 11.465 ;
      RECT 69.615 15.735 69.765 15.885 ;
      RECT 69.615 16.755 69.765 16.905 ;
      RECT 69.615 18.795 69.765 18.945 ;
      RECT 69.615 27.635 69.765 27.785 ;
      RECT 69.615 29.335 69.765 29.485 ;
      RECT 69.615 33.755 69.765 33.905 ;
      RECT 69.615 38.515 69.765 38.665 ;
      RECT 68.695 9.895 68.845 10.045 ;
      RECT 68.695 15.225 68.845 15.375 ;
      RECT 68.695 20.665 68.845 20.815 ;
      RECT 68.695 26.105 68.845 26.255 ;
      RECT 68.695 31.545 68.845 31.695 ;
      RECT 68.695 36.985 68.845 37.135 ;
      RECT 68.695 42.425 68.845 42.575 ;
      RECT 68.695 47.865 68.845 48.015 ;
      RECT 68.695 53.305 68.845 53.455 ;
      RECT 68.695 58.745 68.845 58.895 ;
      RECT 67.775 12.505 67.925 12.655 ;
      RECT 67.775 17.945 67.925 18.095 ;
      RECT 67.775 23.385 67.925 23.535 ;
      RECT 67.775 28.825 67.925 28.975 ;
      RECT 67.775 34.265 67.925 34.415 ;
      RECT 67.775 39.705 67.925 39.855 ;
      RECT 67.775 45.145 67.925 45.295 ;
      RECT 67.775 50.585 67.925 50.735 ;
      RECT 67.775 56.025 67.925 56.175 ;
      RECT 66.855 13.695 67.005 13.845 ;
      RECT 66.855 14.715 67.005 14.865 ;
      RECT 66.855 17.095 67.005 17.245 ;
      RECT 66.855 19.135 67.005 19.285 ;
      RECT 66.855 21.855 67.005 22.005 ;
      RECT 66.855 22.535 67.005 22.685 ;
      RECT 66.855 24.575 67.005 24.725 ;
      RECT 66.855 25.255 67.005 25.405 ;
      RECT 66.855 29.335 67.005 29.485 ;
      RECT 65.935 9.895 66.085 10.045 ;
      RECT 65.935 15.225 66.085 15.375 ;
      RECT 65.935 20.665 66.085 20.815 ;
      RECT 65.935 26.105 66.085 26.255 ;
      RECT 65.935 31.545 66.085 31.695 ;
      RECT 65.935 36.985 66.085 37.135 ;
      RECT 65.935 42.425 66.085 42.575 ;
      RECT 65.935 47.865 66.085 48.015 ;
      RECT 65.935 53.305 66.085 53.455 ;
      RECT 65.935 58.745 66.085 58.895 ;
      RECT 65.015 12.505 65.165 12.655 ;
      RECT 65.015 17.945 65.165 18.095 ;
      RECT 65.015 23.385 65.165 23.535 ;
      RECT 65.015 28.825 65.165 28.975 ;
      RECT 65.015 34.265 65.165 34.415 ;
      RECT 65.015 39.705 65.165 39.855 ;
      RECT 65.015 45.145 65.165 45.295 ;
      RECT 65.015 50.585 65.165 50.735 ;
      RECT 65.015 56.025 65.165 56.175 ;
      RECT 64.095 14.375 64.245 14.525 ;
      RECT 64.095 18.795 64.245 18.945 ;
      RECT 64.095 21.175 64.245 21.325 ;
      RECT 64.095 22.195 64.245 22.345 ;
      RECT 64.095 22.875 64.245 23.025 ;
      RECT 64.095 28.315 64.245 28.465 ;
      RECT 63.175 9.895 63.325 10.045 ;
      RECT 63.175 15.225 63.325 15.375 ;
      RECT 63.175 20.665 63.325 20.815 ;
      RECT 63.175 26.105 63.325 26.255 ;
      RECT 63.175 31.545 63.325 31.695 ;
      RECT 63.175 36.985 63.325 37.135 ;
      RECT 63.175 42.425 63.325 42.575 ;
      RECT 63.175 47.865 63.325 48.015 ;
      RECT 63.175 53.305 63.325 53.455 ;
      RECT 63.175 58.745 63.325 58.895 ;
      RECT 62.255 12.505 62.405 12.655 ;
      RECT 62.255 17.945 62.405 18.095 ;
      RECT 62.255 23.385 62.405 23.535 ;
      RECT 62.255 28.825 62.405 28.975 ;
      RECT 62.255 34.265 62.405 34.415 ;
      RECT 62.255 39.705 62.405 39.855 ;
      RECT 62.255 45.145 62.405 45.295 ;
      RECT 62.255 50.585 62.405 50.735 ;
      RECT 62.255 56.025 62.405 56.175 ;
      RECT 61.335 13.355 61.485 13.505 ;
      RECT 61.335 17.435 61.485 17.585 ;
      RECT 61.335 19.135 61.485 19.285 ;
      RECT 61.335 23.895 61.485 24.045 ;
      RECT 61.335 26.615 61.485 26.765 ;
      RECT 60.415 9.895 60.565 10.045 ;
      RECT 60.415 15.225 60.565 15.375 ;
      RECT 60.415 20.665 60.565 20.815 ;
      RECT 60.415 26.105 60.565 26.255 ;
      RECT 60.415 31.545 60.565 31.695 ;
      RECT 60.415 36.985 60.565 37.135 ;
      RECT 60.415 42.425 60.565 42.575 ;
      RECT 60.415 47.865 60.565 48.015 ;
      RECT 60.415 53.305 60.565 53.455 ;
      RECT 60.415 58.745 60.565 58.895 ;
      RECT 59.495 12.505 59.645 12.655 ;
      RECT 59.495 17.945 59.645 18.095 ;
      RECT 59.495 23.385 59.645 23.535 ;
      RECT 59.495 28.825 59.645 28.975 ;
      RECT 59.495 34.265 59.645 34.415 ;
      RECT 59.495 39.705 59.645 39.855 ;
      RECT 59.495 45.145 59.645 45.295 ;
      RECT 59.495 50.585 59.645 50.735 ;
      RECT 59.495 56.025 59.645 56.175 ;
      RECT 58.575 11.995 58.725 12.145 ;
      RECT 58.575 13.355 58.725 13.505 ;
      RECT 58.575 14.375 58.725 14.525 ;
      RECT 58.575 17.435 58.725 17.585 ;
      RECT 58.575 18.455 58.725 18.605 ;
      RECT 58.575 19.135 58.725 19.285 ;
      RECT 58.575 21.855 58.725 22.005 ;
      RECT 58.575 22.535 58.725 22.685 ;
      RECT 58.575 26.615 58.725 26.765 ;
      RECT 57.655 9.895 57.805 10.045 ;
      RECT 57.655 15.225 57.805 15.375 ;
      RECT 57.655 20.665 57.805 20.815 ;
      RECT 57.655 26.105 57.805 26.255 ;
      RECT 57.655 31.545 57.805 31.695 ;
      RECT 57.655 36.985 57.805 37.135 ;
      RECT 57.655 42.425 57.805 42.575 ;
      RECT 57.655 47.865 57.805 48.015 ;
      RECT 57.655 53.305 57.805 53.455 ;
      RECT 57.655 58.745 57.805 58.895 ;
      RECT 56.735 12.505 56.885 12.655 ;
      RECT 56.735 17.945 56.885 18.095 ;
      RECT 56.735 23.385 56.885 23.535 ;
      RECT 56.735 28.825 56.885 28.975 ;
      RECT 56.735 34.265 56.885 34.415 ;
      RECT 56.735 39.705 56.885 39.855 ;
      RECT 56.735 45.145 56.885 45.295 ;
      RECT 56.735 50.585 56.885 50.735 ;
      RECT 56.735 56.025 56.885 56.175 ;
      RECT 55.815 11.995 55.965 12.145 ;
      RECT 55.815 13.695 55.965 13.845 ;
      RECT 55.815 14.375 55.965 14.525 ;
      RECT 55.815 18.455 55.965 18.605 ;
      RECT 55.815 19.815 55.965 19.965 ;
      RECT 55.815 21.855 55.965 22.005 ;
      RECT 54.895 9.895 55.045 10.045 ;
      RECT 54.895 15.225 55.045 15.375 ;
      RECT 54.895 20.665 55.045 20.815 ;
      RECT 54.895 26.105 55.045 26.255 ;
      RECT 54.895 31.545 55.045 31.695 ;
      RECT 54.895 36.985 55.045 37.135 ;
      RECT 54.895 42.425 55.045 42.575 ;
      RECT 54.895 47.865 55.045 48.015 ;
      RECT 54.895 53.305 55.045 53.455 ;
      RECT 54.895 58.745 55.045 58.895 ;
      RECT 53.975 12.505 54.125 12.655 ;
      RECT 53.975 17.945 54.125 18.095 ;
      RECT 53.975 23.385 54.125 23.535 ;
      RECT 53.975 28.825 54.125 28.975 ;
      RECT 53.975 34.265 54.125 34.415 ;
      RECT 53.975 39.705 54.125 39.855 ;
      RECT 53.975 45.145 54.125 45.295 ;
      RECT 53.975 50.585 54.125 50.735 ;
      RECT 53.975 56.025 54.125 56.175 ;
      RECT 53.055 9.275 53.205 9.425 ;
      RECT 53.055 13.695 53.205 13.845 ;
      RECT 53.055 24.915 53.205 25.065 ;
      RECT 53.055 25.595 53.205 25.745 ;
      RECT 53.055 27.975 53.205 28.125 ;
      RECT 52.135 9.895 52.285 10.045 ;
      RECT 52.135 15.225 52.285 15.375 ;
      RECT 52.135 20.665 52.285 20.815 ;
      RECT 52.135 26.105 52.285 26.255 ;
      RECT 52.135 31.545 52.285 31.695 ;
      RECT 52.135 36.985 52.285 37.135 ;
      RECT 52.135 42.425 52.285 42.575 ;
      RECT 52.135 47.865 52.285 48.015 ;
      RECT 52.135 53.305 52.285 53.455 ;
      RECT 52.135 58.745 52.285 58.895 ;
      RECT 51.215 12.505 51.365 12.655 ;
      RECT 51.215 17.945 51.365 18.095 ;
      RECT 51.215 23.385 51.365 23.535 ;
      RECT 51.215 28.825 51.365 28.975 ;
      RECT 51.215 34.265 51.365 34.415 ;
      RECT 51.215 39.705 51.365 39.855 ;
      RECT 51.215 45.145 51.365 45.295 ;
      RECT 51.215 50.585 51.365 50.735 ;
      RECT 51.215 56.025 51.365 56.175 ;
      RECT 50.295 14.035 50.445 14.185 ;
      RECT 50.295 14.715 50.445 14.865 ;
      RECT 50.295 17.095 50.445 17.245 ;
      RECT 50.295 25.255 50.445 25.405 ;
      RECT 50.295 26.615 50.445 26.765 ;
      RECT 49.375 9.895 49.525 10.045 ;
      RECT 49.375 15.225 49.525 15.375 ;
      RECT 49.375 20.665 49.525 20.815 ;
      RECT 49.375 26.105 49.525 26.255 ;
      RECT 49.375 31.545 49.525 31.695 ;
      RECT 49.375 36.985 49.525 37.135 ;
      RECT 49.375 42.425 49.525 42.575 ;
      RECT 49.375 47.865 49.525 48.015 ;
      RECT 49.375 53.305 49.525 53.455 ;
      RECT 49.375 58.745 49.525 58.895 ;
      RECT 48.455 12.505 48.605 12.655 ;
      RECT 48.455 17.945 48.605 18.095 ;
      RECT 48.455 23.385 48.605 23.535 ;
      RECT 48.455 28.825 48.605 28.975 ;
      RECT 48.455 34.265 48.605 34.415 ;
      RECT 48.455 39.705 48.605 39.855 ;
      RECT 48.455 45.145 48.605 45.295 ;
      RECT 48.455 50.585 48.605 50.735 ;
      RECT 48.455 56.025 48.605 56.175 ;
      RECT 47.535 10.295 47.685 10.445 ;
      RECT 47.535 11.315 47.685 11.465 ;
      RECT 47.535 13.015 47.685 13.165 ;
      RECT 47.535 14.375 47.685 14.525 ;
      RECT 47.535 15.735 47.685 15.885 ;
      RECT 47.535 16.755 47.685 16.905 ;
      RECT 47.535 19.135 47.685 19.285 ;
      RECT 47.535 21.855 47.685 22.005 ;
      RECT 47.535 26.615 47.685 26.765 ;
      RECT 47.535 27.975 47.685 28.125 ;
      RECT 47.535 34.775 47.685 34.925 ;
      RECT 46.615 9.895 46.765 10.045 ;
      RECT 46.615 15.225 46.765 15.375 ;
      RECT 46.615 20.665 46.765 20.815 ;
      RECT 46.615 26.105 46.765 26.255 ;
      RECT 46.615 31.545 46.765 31.695 ;
      RECT 46.615 36.985 46.765 37.135 ;
      RECT 46.615 42.425 46.765 42.575 ;
      RECT 46.615 47.865 46.765 48.015 ;
      RECT 46.615 53.305 46.765 53.455 ;
      RECT 46.615 58.745 46.765 58.895 ;
      RECT 45.695 12.505 45.845 12.655 ;
      RECT 45.695 17.945 45.845 18.095 ;
      RECT 45.695 23.385 45.845 23.535 ;
      RECT 45.695 28.825 45.845 28.975 ;
      RECT 45.695 34.265 45.845 34.415 ;
      RECT 45.695 39.705 45.845 39.855 ;
      RECT 45.695 45.145 45.845 45.295 ;
      RECT 45.695 50.585 45.845 50.735 ;
      RECT 45.695 56.025 45.845 56.175 ;
      RECT 44.775 11.655 44.925 11.805 ;
      RECT 44.775 13.015 44.925 13.165 ;
      RECT 44.775 14.035 44.925 14.185 ;
      RECT 44.775 14.715 44.925 14.865 ;
      RECT 44.775 18.455 44.925 18.605 ;
      RECT 44.775 22.875 44.925 23.025 ;
      RECT 44.775 26.955 44.925 27.105 ;
      RECT 44.775 32.395 44.925 32.545 ;
      RECT 43.855 9.895 44.005 10.045 ;
      RECT 43.855 15.225 44.005 15.375 ;
      RECT 43.855 20.665 44.005 20.815 ;
      RECT 43.855 26.105 44.005 26.255 ;
      RECT 43.855 31.545 44.005 31.695 ;
      RECT 43.855 36.985 44.005 37.135 ;
      RECT 43.855 42.425 44.005 42.575 ;
      RECT 43.855 47.865 44.005 48.015 ;
      RECT 43.855 53.305 44.005 53.455 ;
      RECT 43.855 58.745 44.005 58.895 ;
      RECT 42.935 12.505 43.085 12.655 ;
      RECT 42.935 17.945 43.085 18.095 ;
      RECT 42.935 23.385 43.085 23.535 ;
      RECT 42.935 28.825 43.085 28.975 ;
      RECT 42.935 34.265 43.085 34.415 ;
      RECT 42.935 39.705 43.085 39.855 ;
      RECT 42.935 45.145 43.085 45.295 ;
      RECT 42.935 50.585 43.085 50.735 ;
      RECT 42.935 56.025 43.085 56.175 ;
      RECT 42.015 11.315 42.165 11.465 ;
      RECT 42.015 13.355 42.165 13.505 ;
      RECT 42.015 15.735 42.165 15.885 ;
      RECT 42.015 17.435 42.165 17.585 ;
      RECT 42.015 18.455 42.165 18.605 ;
      RECT 42.015 29.675 42.165 29.825 ;
      RECT 42.015 34.775 42.165 34.925 ;
      RECT 41.095 9.895 41.245 10.045 ;
      RECT 41.095 15.225 41.245 15.375 ;
      RECT 41.095 20.665 41.245 20.815 ;
      RECT 41.095 26.105 41.245 26.255 ;
      RECT 41.095 31.545 41.245 31.695 ;
      RECT 41.095 36.985 41.245 37.135 ;
      RECT 41.095 42.425 41.245 42.575 ;
      RECT 41.095 47.865 41.245 48.015 ;
      RECT 41.095 53.305 41.245 53.455 ;
      RECT 41.095 58.745 41.245 58.895 ;
      RECT 40.175 12.505 40.325 12.655 ;
      RECT 40.175 17.945 40.325 18.095 ;
      RECT 40.175 23.385 40.325 23.535 ;
      RECT 40.175 28.825 40.325 28.975 ;
      RECT 40.175 34.265 40.325 34.415 ;
      RECT 40.175 39.705 40.325 39.855 ;
      RECT 40.175 45.145 40.325 45.295 ;
      RECT 40.175 50.585 40.325 50.735 ;
      RECT 40.175 56.025 40.325 56.175 ;
      RECT 39.715 9.275 39.865 9.425 ;
      RECT 39.255 13.015 39.405 13.165 ;
      RECT 39.255 24.575 39.405 24.725 ;
      RECT 39.255 25.595 39.405 25.745 ;
      RECT 39.255 27.975 39.405 28.125 ;
      RECT 39.255 30.015 39.405 30.165 ;
      RECT 39.255 33.075 39.405 33.225 ;
      RECT 38.335 9.895 38.485 10.045 ;
      RECT 38.335 15.225 38.485 15.375 ;
      RECT 38.335 20.665 38.485 20.815 ;
      RECT 38.335 26.105 38.485 26.255 ;
      RECT 38.335 31.545 38.485 31.695 ;
      RECT 38.335 36.985 38.485 37.135 ;
      RECT 38.335 42.425 38.485 42.575 ;
      RECT 38.335 47.865 38.485 48.015 ;
      RECT 38.335 53.305 38.485 53.455 ;
      RECT 38.335 58.745 38.485 58.895 ;
      RECT 37.415 12.505 37.565 12.655 ;
      RECT 37.415 17.945 37.565 18.095 ;
      RECT 37.415 23.385 37.565 23.535 ;
      RECT 37.415 28.825 37.565 28.975 ;
      RECT 37.415 34.265 37.565 34.415 ;
      RECT 37.415 39.705 37.565 39.855 ;
      RECT 37.415 45.145 37.565 45.295 ;
      RECT 37.415 50.585 37.565 50.735 ;
      RECT 37.415 56.025 37.565 56.175 ;
      RECT 36.495 10.975 36.645 11.125 ;
      RECT 36.495 11.995 36.645 12.145 ;
      RECT 36.495 14.035 36.645 14.185 ;
      RECT 36.495 14.715 36.645 14.865 ;
      RECT 36.495 16.755 36.645 16.905 ;
      RECT 36.495 18.795 36.645 18.945 ;
      RECT 36.495 22.875 36.645 23.025 ;
      RECT 36.495 24.235 36.645 24.385 ;
      RECT 36.495 24.915 36.645 25.065 ;
      RECT 36.495 26.615 36.645 26.765 ;
      RECT 36.495 31.035 36.645 31.185 ;
      RECT 36.495 32.055 36.645 32.205 ;
      RECT 36.495 33.755 36.645 33.905 ;
      RECT 36.495 35.115 36.645 35.265 ;
      RECT 35.575 9.895 35.725 10.045 ;
      RECT 35.575 15.225 35.725 15.375 ;
      RECT 35.575 20.665 35.725 20.815 ;
      RECT 35.575 26.105 35.725 26.255 ;
      RECT 35.575 31.545 35.725 31.695 ;
      RECT 35.575 36.985 35.725 37.135 ;
      RECT 35.575 42.425 35.725 42.575 ;
      RECT 35.575 47.865 35.725 48.015 ;
      RECT 35.575 53.305 35.725 53.455 ;
      RECT 35.575 58.745 35.725 58.895 ;
      RECT 34.655 12.505 34.805 12.655 ;
      RECT 34.655 17.945 34.805 18.095 ;
      RECT 34.655 23.385 34.805 23.535 ;
      RECT 34.655 28.825 34.805 28.975 ;
      RECT 34.655 34.265 34.805 34.415 ;
      RECT 34.655 39.705 34.805 39.855 ;
      RECT 34.655 45.145 34.805 45.295 ;
      RECT 34.655 50.585 34.805 50.735 ;
      RECT 34.655 56.025 34.805 56.175 ;
      RECT 33.735 10.635 33.885 10.785 ;
      RECT 33.735 14.035 33.885 14.185 ;
      RECT 33.735 16.755 33.885 16.905 ;
      RECT 33.735 19.135 33.885 19.285 ;
      RECT 33.735 27.635 33.885 27.785 ;
      RECT 33.735 35.455 33.885 35.605 ;
      RECT 32.815 9.895 32.965 10.045 ;
      RECT 32.815 15.225 32.965 15.375 ;
      RECT 32.815 20.665 32.965 20.815 ;
      RECT 32.815 26.105 32.965 26.255 ;
      RECT 32.815 31.545 32.965 31.695 ;
      RECT 32.815 36.985 32.965 37.135 ;
      RECT 32.815 42.425 32.965 42.575 ;
      RECT 32.815 47.865 32.965 48.015 ;
      RECT 32.815 53.305 32.965 53.455 ;
      RECT 32.815 58.745 32.965 58.895 ;
      RECT 31.895 12.505 32.045 12.655 ;
      RECT 31.895 17.945 32.045 18.095 ;
      RECT 31.895 23.385 32.045 23.535 ;
      RECT 31.895 28.825 32.045 28.975 ;
      RECT 31.895 34.265 32.045 34.415 ;
      RECT 31.895 39.705 32.045 39.855 ;
      RECT 31.895 45.145 32.045 45.295 ;
      RECT 31.895 50.585 32.045 50.735 ;
      RECT 31.895 56.025 32.045 56.175 ;
      RECT 30.975 10.295 31.125 10.445 ;
      RECT 30.975 13.695 31.125 13.845 ;
      RECT 30.975 24.575 31.125 24.725 ;
      RECT 30.975 30.015 31.125 30.165 ;
      RECT 30.975 32.735 31.125 32.885 ;
      RECT 30.055 9.895 30.205 10.045 ;
      RECT 30.055 15.225 30.205 15.375 ;
      RECT 30.055 20.665 30.205 20.815 ;
      RECT 30.055 26.105 30.205 26.255 ;
      RECT 30.055 31.545 30.205 31.695 ;
      RECT 30.055 36.985 30.205 37.135 ;
      RECT 30.055 42.425 30.205 42.575 ;
      RECT 30.055 47.865 30.205 48.015 ;
      RECT 30.055 53.305 30.205 53.455 ;
      RECT 30.055 58.745 30.205 58.895 ;
      RECT 29.135 12.505 29.285 12.655 ;
      RECT 29.135 17.945 29.285 18.095 ;
      RECT 29.135 23.385 29.285 23.535 ;
      RECT 29.135 28.825 29.285 28.975 ;
      RECT 29.135 34.265 29.285 34.415 ;
      RECT 29.135 39.705 29.285 39.855 ;
      RECT 29.135 45.145 29.285 45.295 ;
      RECT 29.135 50.585 29.285 50.735 ;
      RECT 29.135 56.025 29.285 56.175 ;
      RECT 28.215 11.995 28.365 12.145 ;
      RECT 28.215 13.015 28.365 13.165 ;
      RECT 28.215 17.435 28.365 17.585 ;
      RECT 28.215 19.135 28.365 19.285 ;
      RECT 28.215 26.615 28.365 26.765 ;
      RECT 28.215 33.415 28.365 33.565 ;
      RECT 27.295 9.895 27.445 10.045 ;
      RECT 27.295 15.225 27.445 15.375 ;
      RECT 27.295 20.665 27.445 20.815 ;
      RECT 27.295 26.105 27.445 26.255 ;
      RECT 27.295 31.545 27.445 31.695 ;
      RECT 27.295 36.985 27.445 37.135 ;
      RECT 27.295 42.425 27.445 42.575 ;
      RECT 27.295 47.865 27.445 48.015 ;
      RECT 27.295 53.305 27.445 53.455 ;
      RECT 27.295 58.745 27.445 58.895 ;
      RECT 26.375 12.505 26.525 12.655 ;
      RECT 26.375 17.945 26.525 18.095 ;
      RECT 26.375 23.385 26.525 23.535 ;
      RECT 26.375 28.825 26.525 28.975 ;
      RECT 26.375 34.265 26.525 34.415 ;
      RECT 26.375 39.705 26.525 39.855 ;
      RECT 26.375 45.145 26.525 45.295 ;
      RECT 26.375 50.585 26.525 50.735 ;
      RECT 26.375 56.025 26.525 56.175 ;
      RECT 25.455 27.975 25.605 28.125 ;
      RECT 25.455 29.335 25.605 29.485 ;
      RECT 24.535 9.895 24.685 10.045 ;
      RECT 24.535 15.225 24.685 15.375 ;
      RECT 24.535 20.665 24.685 20.815 ;
      RECT 24.535 26.105 24.685 26.255 ;
      RECT 24.535 31.545 24.685 31.695 ;
      RECT 24.535 36.985 24.685 37.135 ;
      RECT 24.535 42.425 24.685 42.575 ;
      RECT 24.535 47.865 24.685 48.015 ;
      RECT 24.535 53.305 24.685 53.455 ;
      RECT 24.535 58.745 24.685 58.895 ;
      RECT 23.615 12.505 23.765 12.655 ;
      RECT 23.615 17.945 23.765 18.095 ;
      RECT 23.615 23.385 23.765 23.535 ;
      RECT 23.615 28.825 23.765 28.975 ;
      RECT 23.615 34.265 23.765 34.415 ;
      RECT 23.615 39.705 23.765 39.855 ;
      RECT 23.615 45.145 23.765 45.295 ;
      RECT 23.615 50.585 23.765 50.735 ;
      RECT 23.615 56.025 23.765 56.175 ;
      RECT 21.775 9.895 21.925 10.045 ;
      RECT 21.775 15.225 21.925 15.375 ;
      RECT 21.775 20.665 21.925 20.815 ;
      RECT 21.775 26.105 21.925 26.255 ;
      RECT 21.775 31.545 21.925 31.695 ;
      RECT 21.775 36.985 21.925 37.135 ;
      RECT 21.775 42.425 21.925 42.575 ;
      RECT 21.775 47.865 21.925 48.015 ;
      RECT 21.775 53.305 21.925 53.455 ;
      RECT 21.775 58.745 21.925 58.895 ;
      RECT 20.855 12.505 21.005 12.655 ;
      RECT 20.855 17.945 21.005 18.095 ;
      RECT 20.855 23.385 21.005 23.535 ;
      RECT 20.855 28.825 21.005 28.975 ;
      RECT 20.855 34.265 21.005 34.415 ;
      RECT 20.855 39.705 21.005 39.855 ;
      RECT 20.855 45.145 21.005 45.295 ;
      RECT 20.855 50.585 21.005 50.735 ;
      RECT 20.855 56.025 21.005 56.175 ;
      RECT 19.935 22.195 20.085 22.345 ;
      RECT 19.935 28.315 20.085 28.465 ;
      RECT 19.935 29.675 20.085 29.825 ;
      RECT 19.015 9.895 19.165 10.045 ;
      RECT 19.015 15.225 19.165 15.375 ;
      RECT 19.015 20.665 19.165 20.815 ;
      RECT 19.015 26.105 19.165 26.255 ;
      RECT 19.015 31.545 19.165 31.695 ;
      RECT 19.015 36.985 19.165 37.135 ;
      RECT 19.015 42.425 19.165 42.575 ;
      RECT 19.015 47.865 19.165 48.015 ;
      RECT 19.015 53.305 19.165 53.455 ;
      RECT 19.015 58.745 19.165 58.895 ;
      RECT 18.095 12.505 18.245 12.655 ;
      RECT 18.095 17.945 18.245 18.095 ;
      RECT 18.095 23.385 18.245 23.535 ;
      RECT 18.095 28.825 18.245 28.975 ;
      RECT 18.095 34.265 18.245 34.415 ;
      RECT 18.095 39.705 18.245 39.855 ;
      RECT 18.095 45.145 18.245 45.295 ;
      RECT 18.095 50.585 18.245 50.735 ;
      RECT 18.095 56.025 18.245 56.175 ;
      RECT 16.255 9.895 16.405 10.045 ;
      RECT 16.255 15.225 16.405 15.375 ;
      RECT 16.255 20.665 16.405 20.815 ;
      RECT 16.255 26.105 16.405 26.255 ;
      RECT 16.255 31.545 16.405 31.695 ;
      RECT 16.255 36.985 16.405 37.135 ;
      RECT 16.255 42.425 16.405 42.575 ;
      RECT 16.255 47.865 16.405 48.015 ;
      RECT 16.255 53.305 16.405 53.455 ;
      RECT 16.255 58.745 16.405 58.895 ;
      RECT 15.335 12.505 15.485 12.655 ;
      RECT 15.335 17.945 15.485 18.095 ;
      RECT 15.335 23.385 15.485 23.535 ;
      RECT 15.335 28.825 15.485 28.975 ;
      RECT 15.335 34.265 15.485 34.415 ;
      RECT 15.335 39.705 15.485 39.855 ;
      RECT 15.335 45.145 15.485 45.295 ;
      RECT 15.335 50.585 15.485 50.735 ;
      RECT 15.335 56.025 15.485 56.175 ;
    LAYER met2 ;
      RECT 179.96 16.67 180.22 16.99 ;
      RECT 180.02 11.91 180.16 16.99 ;
      RECT 179.96 11.91 180.22 12.23 ;
      RECT 177.2 15.335 177.46 15.97 ;
      RECT 177.19 15.335 177.47 15.705 ;
      RECT 177.26 11.23 177.4 15.97 ;
      RECT 177.2 11.23 177.46 11.55 ;
      RECT 177.2 19.39 177.46 19.71 ;
      RECT 177.26 17.35 177.4 19.71 ;
      RECT 177.2 17.35 177.46 17.67 ;
      RECT 171.68 20.07 171.94 20.39 ;
      RECT 171.74 19.05 171.88 20.39 ;
      RECT 171.68 19.05 171.94 19.37 ;
      RECT 171.28 19.14 171.94 19.28 ;
      RECT 171.28 16.42 171.42 19.28 ;
      RECT 171.28 16.42 171.88 16.56 ;
      RECT 171.74 14.63 171.88 16.56 ;
      RECT 171.68 14.63 171.94 14.95 ;
      RECT 171.68 18.37 171.94 18.69 ;
      RECT 171.74 17.35 171.88 18.69 ;
      RECT 171.68 17.35 171.94 17.67 ;
      RECT 168.92 18.37 169.18 18.69 ;
      RECT 168.98 9.235 169.12 18.69 ;
      RECT 168.92 15.65 169.18 15.97 ;
      RECT 168.92 11.23 169.18 11.55 ;
      RECT 168.91 9.235 169.19 9.605 ;
      RECT 168.92 26.87 169.18 27.19 ;
      RECT 168.98 22.11 169.12 27.19 ;
      RECT 168.92 22.11 169.18 22.43 ;
      RECT 163.4 23.81 163.66 24.13 ;
      RECT 163.46 14.29 163.6 24.13 ;
      RECT 163.4 15.65 163.66 15.97 ;
      RECT 163.4 14.29 163.66 14.61 ;
      RECT 160.64 16.555 160.9 16.99 ;
      RECT 160.63 16.555 160.91 16.925 ;
      RECT 160.63 19.605 160.91 19.975 ;
      RECT 160.64 19.39 160.9 19.975 ;
      RECT 160.64 33.33 160.9 33.65 ;
      RECT 160.7 29.93 160.84 33.65 ;
      RECT 160.64 29.93 160.9 30.25 ;
      RECT 157.88 19.05 158.14 19.37 ;
      RECT 157.88 19.14 158.54 19.28 ;
      RECT 158.4 16.42 158.54 19.28 ;
      RECT 157.94 16.42 158.54 16.56 ;
      RECT 157.94 15.335 158.08 16.56 ;
      RECT 157.87 15.335 158.15 15.705 ;
      RECT 157.88 34.69 158.14 35.01 ;
      RECT 157.94 33.42 158.08 35.01 ;
      RECT 157.94 33.42 158.54 33.56 ;
      RECT 158.4 27.3 158.54 33.56 ;
      RECT 157.88 27.21 158.14 27.53 ;
      RECT 157.88 27.3 158.54 27.44 ;
      RECT 157.88 18.37 158.14 18.69 ;
      RECT 157.94 17.35 158.08 18.69 ;
      RECT 157.88 17.35 158.14 17.67 ;
      RECT 157.88 32.65 158.14 32.97 ;
      RECT 157.48 32.74 158.14 32.88 ;
      RECT 157.48 25.26 157.62 32.88 ;
      RECT 157.88 27.89 158.14 28.21 ;
      RECT 157.48 27.98 158.14 28.12 ;
      RECT 157.88 25.17 158.14 25.49 ;
      RECT 157.48 25.26 158.14 25.4 ;
      RECT 155.12 32.31 155.38 32.63 ;
      RECT 155.18 11.23 155.32 32.63 ;
      RECT 155.12 29.25 155.38 29.57 ;
      RECT 155.12 24.49 155.38 24.81 ;
      RECT 155.12 11.23 155.38 11.55 ;
      RECT 155.12 35.03 155.38 35.35 ;
      RECT 155.18 33.67 155.32 35.35 ;
      RECT 155.12 33.67 155.38 33.99 ;
      RECT 152.36 31.97 152.62 32.29 ;
      RECT 152.36 32.06 153.02 32.2 ;
      RECT 152.88 19.82 153.02 32.2 ;
      RECT 152.36 26.53 152.62 26.85 ;
      RECT 152.36 26.62 153.02 26.76 ;
      RECT 152.36 19.73 152.62 20.05 ;
      RECT 152.36 19.82 153.02 19.96 ;
      RECT 152.36 18.37 152.62 18.69 ;
      RECT 152.42 11.23 152.56 18.69 ;
      RECT 152.36 15.65 152.62 15.97 ;
      RECT 152.36 12.93 152.62 13.25 ;
      RECT 152.36 11.23 152.62 11.55 ;
      RECT 151.96 34.1 152.56 34.24 ;
      RECT 152.42 32.99 152.56 34.24 ;
      RECT 151.96 19.14 152.1 34.24 ;
      RECT 152.36 32.99 152.62 33.31 ;
      RECT 152.36 27.55 152.62 27.87 ;
      RECT 151.96 27.64 152.62 27.78 ;
      RECT 152.36 23.81 152.62 24.13 ;
      RECT 151.96 23.9 152.62 24.04 ;
      RECT 152.36 19.05 152.62 19.37 ;
      RECT 151.96 19.14 152.62 19.28 ;
      RECT 152.36 29.59 152.62 29.91 ;
      RECT 152.42 28.23 152.56 29.91 ;
      RECT 152.36 28.23 152.62 28.55 ;
      RECT 149.6 19.05 149.86 19.37 ;
      RECT 149.6 19.14 150.26 19.28 ;
      RECT 150.12 16.08 150.26 19.28 ;
      RECT 149.66 16.08 150.26 16.22 ;
      RECT 149.66 10.3 149.8 16.22 ;
      RECT 149.66 10.3 150.26 10.44 ;
      RECT 150.12 9.235 150.26 10.44 ;
      RECT 150.05 9.235 150.33 9.605 ;
      RECT 149.6 25.17 149.86 25.49 ;
      RECT 149.66 22.79 149.8 25.49 ;
      RECT 149.59 24.485 149.87 24.855 ;
      RECT 149.6 22.79 149.86 23.11 ;
      RECT 149.6 18.37 149.86 18.69 ;
      RECT 149.66 17.01 149.8 18.69 ;
      RECT 149.6 17.01 149.86 17.33 ;
      RECT 149.6 21.43 149.86 21.75 ;
      RECT 149.66 19.73 149.8 21.75 ;
      RECT 149.6 19.73 149.86 20.05 ;
      RECT 146.84 25.51 147.1 25.83 ;
      RECT 146.84 25.6 147.5 25.74 ;
      RECT 147.36 18.46 147.5 25.74 ;
      RECT 146.84 18.37 147.1 18.69 ;
      RECT 146.84 18.46 147.5 18.6 ;
      RECT 146.81 24.86 147.13 25.12 ;
      RECT 146.9 21.77 147.04 25.12 ;
      RECT 146.84 21.77 147.1 22.09 ;
      RECT 146.84 19.05 147.1 19.37 ;
      RECT 146.44 19.14 147.1 19.28 ;
      RECT 146.44 14.38 146.58 19.28 ;
      RECT 146.84 14.29 147.1 14.61 ;
      RECT 146.44 14.38 147.1 14.52 ;
      RECT 146.84 26.53 147.1 26.85 ;
      RECT 146.44 26.62 147.1 26.76 ;
      RECT 146.44 21.18 146.58 26.76 ;
      RECT 146.84 21.09 147.1 21.41 ;
      RECT 146.44 21.18 147.1 21.32 ;
      RECT 144.08 26.53 144.34 26.85 ;
      RECT 144.14 22.79 144.28 26.85 ;
      RECT 144.08 24.49 144.34 24.81 ;
      RECT 144.08 22.79 144.34 23.11 ;
      RECT 141.32 21.77 141.58 22.09 ;
      RECT 141.38 20.825 141.52 22.09 ;
      RECT 141.31 20.825 141.59 21.195 ;
      RECT 141.32 18.37 141.58 18.69 ;
      RECT 141.38 17.35 141.52 18.69 ;
      RECT 141.32 17.35 141.58 17.67 ;
      RECT 141.32 27.89 141.58 28.21 ;
      RECT 141.38 25.51 141.52 28.21 ;
      RECT 141.32 25.51 141.58 25.83 ;
      RECT 138.56 29.93 138.82 30.25 ;
      RECT 138.62 16.555 138.76 30.25 ;
      RECT 138.56 27.21 138.82 27.53 ;
      RECT 138.56 19.05 138.82 19.37 ;
      RECT 138.55 16.555 138.83 16.925 ;
      RECT 138.56 15.65 138.82 15.97 ;
      RECT 138.62 14.63 138.76 15.97 ;
      RECT 138.56 14.63 138.82 14.95 ;
      RECT 135.79 23.875 136.07 24.245 ;
      RECT 135.86 22.79 136 24.245 ;
      RECT 135.8 22.79 136.06 23.11 ;
      RECT 135.8 24.49 136.06 24.81 ;
      RECT 135.4 24.58 136.06 24.72 ;
      RECT 135.4 13.02 135.54 24.72 ;
      RECT 135.8 12.93 136.06 13.25 ;
      RECT 135.4 13.02 136.06 13.16 ;
      RECT 135.8 21.43 136.06 21.75 ;
      RECT 135.86 16.67 136 21.75 ;
      RECT 135.8 16.67 136.06 16.99 ;
      RECT 135.8 26.87 136.06 27.19 ;
      RECT 135.86 25.51 136 27.19 ;
      RECT 135.8 25.51 136.06 25.83 ;
      RECT 135.8 34.69 136.06 35.01 ;
      RECT 135.86 27.89 136 35.01 ;
      RECT 135.8 27.89 136.06 28.21 ;
      RECT 133.04 26.87 133.3 27.19 ;
      RECT 133.04 26.96 133.7 27.1 ;
      RECT 133.56 21.18 133.7 27.1 ;
      RECT 133.04 20.825 133.3 21.41 ;
      RECT 133.04 21.18 133.7 21.32 ;
      RECT 133.03 20.825 133.31 21.195 ;
      RECT 133.03 19.605 133.31 19.975 ;
      RECT 133.1 16.67 133.24 19.975 ;
      RECT 133.04 16.67 133.3 16.99 ;
      RECT 133.03 28.755 133.31 29.125 ;
      RECT 132.64 28.66 133.24 28.8 ;
      RECT 132.64 22.2 132.78 28.8 ;
      RECT 133.04 25.51 133.3 25.83 ;
      RECT 132.64 25.6 133.3 25.74 ;
      RECT 133.04 22.11 133.3 22.43 ;
      RECT 132.64 22.2 133.3 22.34 ;
      RECT 133.04 14.29 133.3 14.61 ;
      RECT 133.1 11.23 133.24 14.61 ;
      RECT 133.04 11.23 133.3 11.55 ;
      RECT 133.04 24.83 133.3 25.15 ;
      RECT 133.1 22.79 133.24 25.15 ;
      RECT 133.04 22.79 133.3 23.11 ;
      RECT 130.28 22.11 130.54 22.43 ;
      RECT 130.34 20.07 130.48 22.43 ;
      RECT 130.34 21.18 130.94 21.32 ;
      RECT 130.8 14.38 130.94 21.32 ;
      RECT 130.28 20.07 130.54 20.39 ;
      RECT 130.28 14.29 130.54 14.61 ;
      RECT 130.28 14.38 130.94 14.52 ;
      RECT 130.28 23.81 130.54 24.13 ;
      RECT 130.34 23.22 130.48 24.13 ;
      RECT 129.88 23.22 130.48 23.36 ;
      RECT 129.88 19.14 130.02 23.36 ;
      RECT 130.28 19.05 130.54 19.37 ;
      RECT 129.88 19.14 130.54 19.28 ;
      RECT 130.28 27.21 130.54 27.53 ;
      RECT 130.34 24.83 130.48 27.53 ;
      RECT 130.28 26.53 130.54 26.85 ;
      RECT 130.28 24.83 130.54 25.15 ;
      RECT 130.28 29.25 130.54 29.57 ;
      RECT 130.34 28.23 130.48 29.57 ;
      RECT 130.28 28.23 130.54 28.55 ;
      RECT 130.28 34.69 130.54 35.01 ;
      RECT 130.34 33.33 130.48 35.01 ;
      RECT 130.28 33.33 130.54 33.65 ;
      RECT 127.52 20.825 127.78 21.41 ;
      RECT 127.51 20.825 127.79 21.195 ;
      RECT 127.51 28.145 127.79 28.515 ;
      RECT 127.58 25.51 127.72 28.515 ;
      RECT 127.52 27.55 127.78 27.87 ;
      RECT 127.52 25.51 127.78 25.83 ;
      RECT 127.52 24.49 127.78 24.81 ;
      RECT 127.58 22.11 127.72 24.81 ;
      RECT 127.52 22.11 127.78 22.43 ;
      RECT 127.52 34.69 127.78 35.01 ;
      RECT 127.58 29.25 127.72 35.01 ;
      RECT 127.52 29.25 127.78 29.57 ;
      RECT 124.76 15.335 125.02 15.97 ;
      RECT 124.75 15.335 125.03 15.705 ;
      RECT 124.82 11.23 124.96 15.97 ;
      RECT 124.76 11.23 125.02 11.55 ;
      RECT 124.76 35.37 125.02 35.69 ;
      RECT 124.82 16.555 124.96 35.69 ;
      RECT 124.76 22.11 125.02 22.43 ;
      RECT 124.76 20.07 125.02 20.39 ;
      RECT 124.75 16.555 125.03 16.925 ;
      RECT 122 19.05 122.26 19.37 ;
      RECT 122.06 14.115 122.2 19.37 ;
      RECT 122 14.63 122.26 14.95 ;
      RECT 121.99 14.115 122.27 14.485 ;
      RECT 122 26.87 122.26 27.19 ;
      RECT 122.06 23.875 122.2 27.19 ;
      RECT 121.99 23.875 122.27 24.245 ;
      RECT 119.23 19.605 119.51 19.975 ;
      RECT 119.3 17.01 119.44 19.975 ;
      RECT 119.24 18.37 119.5 18.69 ;
      RECT 119.24 17.01 119.5 17.33 ;
      RECT 119.24 21.77 119.5 22.09 ;
      RECT 119.3 20.5 119.44 22.09 ;
      RECT 119.23 20.825 119.51 21.195 ;
      RECT 118.84 20.5 119.44 20.64 ;
      RECT 118.84 13.7 118.98 20.64 ;
      RECT 118.84 13.7 119.44 13.84 ;
      RECT 119.3 11.23 119.44 13.84 ;
      RECT 119.24 11.23 119.5 11.55 ;
      RECT 119.24 15.65 119.5 15.97 ;
      RECT 119.3 14.63 119.44 15.97 ;
      RECT 119.24 14.63 119.5 14.95 ;
      RECT 119.24 26.53 119.5 26.85 ;
      RECT 119.3 22.45 119.44 26.85 ;
      RECT 119.24 25.51 119.5 25.83 ;
      RECT 119.24 22.45 119.5 22.77 ;
      RECT 116.48 22.11 116.74 22.43 ;
      RECT 116.54 20.825 116.68 22.43 ;
      RECT 116.54 21.18 117.14 21.32 ;
      RECT 117 16.76 117.14 21.32 ;
      RECT 116.47 20.825 116.75 21.195 ;
      RECT 116.45 16.7 116.77 16.96 ;
      RECT 116.45 16.76 117.14 16.9 ;
      RECT 116.48 20.07 116.74 20.39 ;
      RECT 116.08 20.16 116.74 20.3 ;
      RECT 116.08 16.42 116.22 20.3 ;
      RECT 116.08 16.42 116.68 16.56 ;
      RECT 116.54 11.23 116.68 16.56 ;
      RECT 116.48 12.93 116.74 13.25 ;
      RECT 116.48 11.23 116.74 11.55 ;
      RECT 116.48 19.05 116.74 19.37 ;
      RECT 116.54 17.35 116.68 19.37 ;
      RECT 116.48 17.35 116.74 17.67 ;
      RECT 116.48 27.55 116.74 27.87 ;
      RECT 116.54 22.79 116.68 27.87 ;
      RECT 116.48 22.79 116.74 23.11 ;
      RECT 113.72 26.53 113.98 26.85 ;
      RECT 113.78 25.17 113.92 26.85 ;
      RECT 113.72 25.17 113.98 25.49 ;
      RECT 113.32 25.26 113.98 25.4 ;
      RECT 113.32 13.7 113.46 25.4 ;
      RECT 113.69 22.14 114.01 22.4 ;
      RECT 113.78 21.86 113.92 22.4 ;
      RECT 113.32 21.86 113.92 22 ;
      RECT 113.72 18.37 113.98 18.69 ;
      RECT 113.32 18.46 113.98 18.6 ;
      RECT 113.78 17.35 113.92 18.69 ;
      RECT 113.72 17.35 113.98 17.67 ;
      RECT 113.72 13.61 113.98 13.93 ;
      RECT 113.32 13.7 113.98 13.84 ;
      RECT 111.345 22.11 111.605 22.43 ;
      RECT 111.405 16.42 111.545 22.43 ;
      RECT 110.96 16.33 111.22 16.65 ;
      RECT 110.96 16.42 111.545 16.56 ;
      RECT 111.02 13.27 111.16 16.65 ;
      RECT 110.96 13.27 111.22 13.59 ;
      RECT 110.96 29.93 111.22 30.25 ;
      RECT 111.02 18.71 111.16 30.25 ;
      RECT 110.96 27.55 111.22 27.87 ;
      RECT 110.95 19.605 111.23 19.975 ;
      RECT 110.96 18.71 111.22 19.03 ;
      RECT 108.2 22.11 108.46 22.43 ;
      RECT 108.26 20.5 108.4 22.43 ;
      RECT 108.19 20.825 108.47 21.195 ;
      RECT 107.8 20.5 108.4 20.64 ;
      RECT 107.8 15.74 107.94 20.64 ;
      RECT 107.8 15.74 108.4 15.88 ;
      RECT 108.26 14.29 108.4 15.88 ;
      RECT 108.2 14.29 108.46 14.61 ;
      RECT 108.2 18.37 108.46 18.69 ;
      RECT 108.26 17.35 108.4 18.69 ;
      RECT 108.2 17.35 108.46 17.67 ;
      RECT 108.2 29.59 108.46 29.91 ;
      RECT 108.26 22.79 108.4 29.91 ;
      RECT 108.2 22.79 108.46 23.11 ;
      RECT 105.44 20.825 105.7 21.41 ;
      RECT 105.43 20.825 105.71 21.195 ;
      RECT 105.44 25.51 105.7 25.83 ;
      RECT 105.5 21.86 105.64 25.83 ;
      RECT 105.43 23.875 105.71 24.245 ;
      RECT 105.04 21.86 105.64 22 ;
      RECT 105.04 13.7 105.18 22 ;
      RECT 105.44 19.73 105.7 20.05 ;
      RECT 105.04 19.82 105.7 19.96 ;
      RECT 105.44 13.61 105.7 13.93 ;
      RECT 105.04 13.7 105.7 13.84 ;
      RECT 105.44 19.05 105.7 19.37 ;
      RECT 105.5 14.29 105.64 19.37 ;
      RECT 105.44 14.29 105.7 14.61 ;
      RECT 102.67 19.605 102.95 19.975 ;
      RECT 102.74 16.67 102.88 19.975 ;
      RECT 102.68 16.67 102.94 16.99 ;
      RECT 102.68 24.15 102.94 24.47 ;
      RECT 102.74 22.11 102.88 24.47 ;
      RECT 102.68 22.11 102.94 22.43 ;
      RECT 102.68 34.69 102.94 35.01 ;
      RECT 102.74 28.23 102.88 35.01 ;
      RECT 102.68 28.23 102.94 28.55 ;
      RECT 99.92 29.25 100.18 29.57 ;
      RECT 99.98 19.82 100.12 29.57 ;
      RECT 99.92 24.83 100.18 25.15 ;
      RECT 99.91 20.825 100.19 21.195 ;
      RECT 99.52 19.82 100.12 19.96 ;
      RECT 99.52 11.66 99.66 19.96 ;
      RECT 99.92 11.57 100.18 11.89 ;
      RECT 99.52 11.66 100.18 11.8 ;
      RECT 99.92 32.415 100.18 32.97 ;
      RECT 99.91 32.415 100.19 32.785 ;
      RECT 99.92 18.71 100.18 19.03 ;
      RECT 99.98 13.61 100.12 19.03 ;
      RECT 99.92 17.35 100.18 17.67 ;
      RECT 99.92 13.61 100.18 13.93 ;
      RECT 97.16 20.825 97.42 21.41 ;
      RECT 97.15 20.825 97.43 21.195 ;
      RECT 97.16 32.99 97.42 33.31 ;
      RECT 97.22 24.485 97.36 33.31 ;
      RECT 97.15 24.485 97.43 24.855 ;
      RECT 97.16 19.73 97.42 20.05 ;
      RECT 97.22 19.14 97.36 20.05 ;
      RECT 96.76 19.14 97.36 19.28 ;
      RECT 96.76 15.74 96.9 19.28 ;
      RECT 97.16 15.65 97.42 15.97 ;
      RECT 96.76 15.74 97.42 15.88 ;
      RECT 97.22 11.23 97.36 15.97 ;
      RECT 97.16 11.23 97.42 11.55 ;
      RECT 97.16 18.37 97.42 18.69 ;
      RECT 97.22 16.67 97.36 18.69 ;
      RECT 97.16 16.67 97.42 16.99 ;
      RECT 97.16 23.81 97.42 24.13 ;
      RECT 97.22 22.11 97.36 24.13 ;
      RECT 97.16 22.11 97.42 22.43 ;
      RECT 97.16 35.03 97.42 35.35 ;
      RECT 97.22 33.67 97.36 35.35 ;
      RECT 97.16 33.67 97.42 33.99 ;
      RECT 94.39 36.075 94.67 36.445 ;
      RECT 94.46 16.67 94.6 36.445 ;
      RECT 94.4 22.45 94.66 22.77 ;
      RECT 94.39 19.605 94.67 19.975 ;
      RECT 94.4 16.67 94.66 16.99 ;
      RECT 91.63 36.075 91.91 36.445 ;
      RECT 91.63 36.19 92.3 36.33 ;
      RECT 92.16 35.46 92.3 36.33 ;
      RECT 91.64 35.37 91.9 35.69 ;
      RECT 91.64 35.46 92.3 35.6 ;
      RECT 91.63 16.555 91.91 16.925 ;
      RECT 91.7 11.23 91.84 16.925 ;
      RECT 91.64 11.23 91.9 11.55 ;
      RECT 91.64 25.51 91.9 25.83 ;
      RECT 91.7 20.07 91.84 25.83 ;
      RECT 91.63 24.485 91.91 24.855 ;
      RECT 91.64 21.43 91.9 21.75 ;
      RECT 91.64 20.07 91.9 20.39 ;
      RECT 88.88 31.97 89.14 32.29 ;
      RECT 88.94 23.9 89.08 32.29 ;
      RECT 88.88 26.53 89.14 26.85 ;
      RECT 88.88 24.83 89.14 25.15 ;
      RECT 88.94 23.9 89.54 24.04 ;
      RECT 89.4 19.14 89.54 24.04 ;
      RECT 88.88 19.05 89.14 19.37 ;
      RECT 88.88 19.14 89.54 19.28 ;
      RECT 88.87 20.825 89.15 21.195 ;
      RECT 88.94 19.73 89.08 21.195 ;
      RECT 88.88 19.73 89.14 20.05 ;
      RECT 88.88 22.45 89.14 22.77 ;
      RECT 88.48 22.54 89.14 22.68 ;
      RECT 88.48 15.74 88.62 22.68 ;
      RECT 88.88 15.65 89.14 15.97 ;
      RECT 88.48 15.74 89.14 15.88 ;
      RECT 86.09 32 86.41 32.26 ;
      RECT 86.18 22.54 86.32 32.26 ;
      RECT 86.12 25.17 86.38 25.49 ;
      RECT 86.11 24.485 86.39 24.855 ;
      RECT 85.72 22.54 86.32 22.68 ;
      RECT 85.72 19.14 85.86 22.68 ;
      RECT 86.12 19.05 86.38 19.37 ;
      RECT 85.72 19.14 86.38 19.28 ;
      RECT 86.12 32.99 86.38 33.31 ;
      RECT 86.18 32.415 86.32 33.31 ;
      RECT 86.11 32.415 86.39 32.785 ;
      RECT 86.12 18.37 86.38 18.69 ;
      RECT 86.18 17.35 86.32 18.69 ;
      RECT 86.12 17.35 86.38 17.67 ;
      RECT 83.36 24.49 83.62 24.81 ;
      RECT 83.36 24.58 84.02 24.72 ;
      RECT 83.88 22.54 84.02 24.72 ;
      RECT 83.36 22.45 83.62 22.77 ;
      RECT 83.36 22.54 84.02 22.68 ;
      RECT 83.36 13.95 83.62 14.27 ;
      RECT 83.42 11.23 83.56 14.27 ;
      RECT 83.36 11.23 83.62 11.55 ;
      RECT 83.36 19.73 83.62 20.05 ;
      RECT 83.42 17.01 83.56 20.05 ;
      RECT 83.36 17.01 83.62 17.33 ;
      RECT 83.36 26.53 83.62 26.85 ;
      RECT 83.42 25.26 83.56 26.85 ;
      RECT 82.96 25.26 83.56 25.4 ;
      RECT 82.96 21.86 83.1 25.4 ;
      RECT 83.36 21.77 83.62 22.09 ;
      RECT 82.96 21.86 83.62 22 ;
      RECT 80.6 33.67 80.86 33.99 ;
      RECT 80.66 29.34 80.8 33.99 ;
      RECT 80.66 29.34 81.26 29.48 ;
      RECT 81.12 23.9 81.26 29.48 ;
      RECT 80.57 24.18 80.89 24.44 ;
      RECT 80.66 23.9 80.8 24.44 ;
      RECT 80.66 23.9 81.26 24.04 ;
      RECT 80.57 24.86 80.89 25.12 ;
      RECT 80.66 24.58 80.8 25.12 ;
      RECT 80.2 24.58 80.8 24.72 ;
      RECT 80.2 15.74 80.34 24.72 ;
      RECT 80.6 21.77 80.86 22.09 ;
      RECT 80.2 21.86 80.86 22 ;
      RECT 80.6 19.73 80.86 20.05 ;
      RECT 80.2 19.82 80.86 19.96 ;
      RECT 80.2 15.74 80.8 15.88 ;
      RECT 80.66 11.57 80.8 15.88 ;
      RECT 80.6 11.57 80.86 11.89 ;
      RECT 80.6 18.71 80.86 19.03 ;
      RECT 80.66 16.67 80.8 19.03 ;
      RECT 80.6 16.67 80.86 16.99 ;
      RECT 80.6 27.55 80.86 27.87 ;
      RECT 80.66 25.51 80.8 27.87 ;
      RECT 80.6 25.51 80.86 25.83 ;
      RECT 77.84 18.37 78.1 18.69 ;
      RECT 77.9 15.335 78.04 18.69 ;
      RECT 77.83 15.335 78.11 15.705 ;
      RECT 77.84 33.33 78.1 33.65 ;
      RECT 77.9 25.51 78.04 33.65 ;
      RECT 77.84 25.51 78.1 25.83 ;
      RECT 75.465 24.485 75.725 25.15 ;
      RECT 75.455 24.485 75.735 24.855 ;
      RECT 75.08 16.555 75.34 16.99 ;
      RECT 75.07 16.555 75.35 16.925 ;
      RECT 75.08 32.65 75.34 32.97 ;
      RECT 75.14 18.71 75.28 32.97 ;
      RECT 75.08 27.21 75.34 27.53 ;
      RECT 75.08 18.71 75.34 19.03 ;
      RECT 72.32 19.05 72.58 19.37 ;
      RECT 72.38 14.115 72.52 19.37 ;
      RECT 72.31 16.555 72.59 16.925 ;
      RECT 72.31 14.115 72.59 14.485 ;
      RECT 72.32 19.605 72.58 20.05 ;
      RECT 72.31 19.605 72.59 19.975 ;
      RECT 72.32 23.81 72.58 24.13 ;
      RECT 72.38 21.09 72.52 24.13 ;
      RECT 72.32 21.09 72.58 21.41 ;
      RECT 72.32 26.53 72.58 26.85 ;
      RECT 72.38 24.49 72.52 26.85 ;
      RECT 72.32 24.49 72.58 24.81 ;
      RECT 69.56 15.65 69.82 15.97 ;
      RECT 69.62 11.23 69.76 15.97 ;
      RECT 69.56 11.23 69.82 11.55 ;
      RECT 69.56 27.55 69.82 27.87 ;
      RECT 69.62 16.67 69.76 27.87 ;
      RECT 69.56 18.71 69.82 19.03 ;
      RECT 69.56 16.67 69.82 16.99 ;
      RECT 69.56 38.43 69.82 38.75 ;
      RECT 69.62 29.25 69.76 38.75 ;
      RECT 69.56 33.67 69.82 33.99 ;
      RECT 69.56 29.25 69.82 29.57 ;
      RECT 66.8 21.77 67.06 22.09 ;
      RECT 66.86 19.82 67 22.09 ;
      RECT 66.4 19.82 67 19.96 ;
      RECT 66.4 13.7 66.54 19.96 ;
      RECT 66.8 19.05 67.06 19.37 ;
      RECT 66.4 19.14 67.06 19.28 ;
      RECT 66.8 13.505 67.06 13.93 ;
      RECT 66.79 13.505 67.07 13.875 ;
      RECT 66.4 13.7 67.07 13.84 ;
      RECT 66.8 17.01 67.06 17.33 ;
      RECT 66.86 14.63 67 17.33 ;
      RECT 66.8 14.63 67.06 14.95 ;
      RECT 66.8 29.25 67.06 29.57 ;
      RECT 66.4 29.34 67.06 29.48 ;
      RECT 66.4 22.54 66.54 29.48 ;
      RECT 66.8 22.45 67.06 22.77 ;
      RECT 66.4 22.54 67.06 22.68 ;
      RECT 66.8 25.17 67.06 25.49 ;
      RECT 66.86 24.49 67 25.49 ;
      RECT 66.8 24.49 67.06 24.81 ;
      RECT 64.04 22.11 64.3 22.43 ;
      RECT 64.1 14.29 64.24 22.43 ;
      RECT 64.04 21.09 64.3 21.41 ;
      RECT 64.04 18.71 64.3 19.03 ;
      RECT 64.04 14.29 64.3 14.61 ;
      RECT 64.04 28.23 64.3 28.55 ;
      RECT 64.1 22.79 64.24 28.55 ;
      RECT 64.04 22.79 64.3 23.11 ;
      RECT 61.28 19.05 61.54 19.37 ;
      RECT 61.28 19.14 61.94 19.28 ;
      RECT 61.8 16.42 61.94 19.28 ;
      RECT 61.27 16.555 61.55 16.925 ;
      RECT 61.34 16.42 61.94 16.56 ;
      RECT 61.27 15.335 61.55 15.705 ;
      RECT 61.34 13.27 61.48 15.705 ;
      RECT 61.28 13.27 61.54 13.59 ;
      RECT 61.28 26.53 61.54 26.85 ;
      RECT 61.34 19.82 61.48 26.85 ;
      RECT 61.28 23.81 61.54 24.13 ;
      RECT 60.88 19.82 61.48 19.96 ;
      RECT 60.88 17.44 61.02 19.96 ;
      RECT 61.28 17.35 61.54 17.67 ;
      RECT 60.88 17.44 61.54 17.58 ;
      RECT 58.52 21.77 58.78 22.09 ;
      RECT 58.58 20.5 58.72 22.09 ;
      RECT 58.58 20.5 59.18 20.64 ;
      RECT 59.04 14.38 59.18 20.64 ;
      RECT 58.52 14.29 58.78 14.61 ;
      RECT 58.52 14.38 59.18 14.52 ;
      RECT 58.51 19.605 58.79 19.975 ;
      RECT 58.58 19.05 58.72 19.975 ;
      RECT 58.52 19.05 58.78 19.37 ;
      RECT 58.52 13.27 58.78 13.59 ;
      RECT 58.58 11.91 58.72 13.59 ;
      RECT 58.52 11.91 58.78 12.23 ;
      RECT 58.52 18.37 58.78 18.69 ;
      RECT 58.58 17.35 58.72 18.69 ;
      RECT 58.52 17.35 58.78 17.67 ;
      RECT 58.52 26.53 58.78 26.85 ;
      RECT 58.58 22.45 58.72 26.85 ;
      RECT 58.52 22.45 58.78 22.77 ;
      RECT 55.75 24.485 56.03 24.855 ;
      RECT 55.82 19.73 55.96 24.855 ;
      RECT 55.76 21.77 56.02 22.09 ;
      RECT 55.76 19.73 56.02 20.05 ;
      RECT 55.76 13.61 56.02 13.93 ;
      RECT 55.82 11.91 55.96 13.93 ;
      RECT 55.76 11.91 56.02 12.23 ;
      RECT 55.76 18.37 56.02 18.69 ;
      RECT 55.82 14.29 55.96 18.69 ;
      RECT 55.76 14.29 56.02 14.61 ;
      RECT 53 13.505 53.26 13.93 ;
      RECT 52.99 13.505 53.27 13.875 ;
      RECT 53.06 9.19 53.2 13.93 ;
      RECT 53 9.19 53.26 9.51 ;
      RECT 53 24.485 53.26 25.15 ;
      RECT 52.99 24.485 53.27 24.855 ;
      RECT 53 27.89 53.26 28.21 ;
      RECT 53.06 25.51 53.2 28.21 ;
      RECT 53 25.51 53.26 25.83 ;
      RECT 50.23 14.115 50.51 14.485 ;
      RECT 50.24 13.95 50.5 14.485 ;
      RECT 50.24 17.01 50.5 17.33 ;
      RECT 50.3 14.63 50.44 17.33 ;
      RECT 50.24 14.63 50.5 14.95 ;
      RECT 50.24 26.53 50.5 26.85 ;
      RECT 50.3 25.17 50.44 26.85 ;
      RECT 50.24 25.17 50.5 25.49 ;
      RECT 47.48 15.65 47.74 15.97 ;
      RECT 47.48 15.74 48.14 15.88 ;
      RECT 48 11.66 48.14 15.88 ;
      RECT 47.48 12.93 47.74 13.25 ;
      RECT 47.48 13.02 48.14 13.16 ;
      RECT 47.54 11.66 48.14 11.8 ;
      RECT 47.54 11.26 47.68 11.8 ;
      RECT 47.45 11.26 47.77 11.52 ;
      RECT 47.47 19.605 47.75 19.975 ;
      RECT 47.54 16.67 47.68 19.975 ;
      RECT 47.48 19.05 47.74 19.37 ;
      RECT 47.48 16.67 47.74 16.99 ;
      RECT 47.48 14.29 47.74 14.61 ;
      RECT 47.08 14.38 47.74 14.52 ;
      RECT 47.08 10.98 47.22 14.52 ;
      RECT 47.08 10.98 47.68 11.12 ;
      RECT 47.54 10.21 47.68 11.12 ;
      RECT 47.48 10.21 47.74 10.53 ;
      RECT 47.48 26.53 47.74 26.85 ;
      RECT 47.54 21.77 47.68 26.85 ;
      RECT 47.48 21.77 47.74 22.09 ;
      RECT 47.48 34.69 47.74 35.01 ;
      RECT 47.54 27.89 47.68 35.01 ;
      RECT 47.48 27.89 47.74 28.21 ;
      RECT 44.71 13.98 44.99 14.485 ;
      RECT 44.69 13.98 45.01 14.24 ;
      RECT 44.72 32.31 44.98 32.63 ;
      RECT 44.78 22.79 44.92 32.63 ;
      RECT 44.72 26.87 44.98 27.19 ;
      RECT 44.71 24.485 44.99 24.855 ;
      RECT 44.72 22.79 44.98 23.11 ;
      RECT 44.72 12.93 44.98 13.25 ;
      RECT 44.78 11.57 44.92 13.25 ;
      RECT 44.72 11.57 44.98 11.89 ;
      RECT 44.72 18.37 44.98 18.69 ;
      RECT 44.78 14.63 44.92 18.69 ;
      RECT 44.72 14.63 44.98 14.95 ;
      RECT 41.96 34.69 42.22 35.01 ;
      RECT 42.02 23.875 42.16 35.01 ;
      RECT 41.96 29.59 42.22 29.91 ;
      RECT 41.95 23.875 42.23 24.245 ;
      RECT 41.96 15.65 42.22 15.97 ;
      RECT 42.02 11.23 42.16 15.97 ;
      RECT 41.96 13.27 42.22 13.59 ;
      RECT 41.96 11.23 42.22 11.55 ;
      RECT 41.96 18.37 42.22 18.69 ;
      RECT 42.02 17.35 42.16 18.69 ;
      RECT 41.96 17.35 42.22 17.67 ;
      RECT 39.2 32.99 39.46 33.31 ;
      RECT 39.26 28.66 39.4 33.31 ;
      RECT 39.2 29.93 39.46 30.25 ;
      RECT 38.8 28.66 39.4 28.8 ;
      RECT 38.8 24.58 38.94 28.8 ;
      RECT 39.2 24.49 39.46 24.81 ;
      RECT 38.8 24.58 39.46 24.72 ;
      RECT 39.26 22.54 39.4 24.81 ;
      RECT 39.26 22.54 39.86 22.68 ;
      RECT 39.72 9.19 39.86 22.68 ;
      RECT 39.2 12.93 39.46 13.25 ;
      RECT 39.2 13.02 39.86 13.16 ;
      RECT 39.66 9.19 39.92 9.51 ;
      RECT 39.2 27.89 39.46 28.21 ;
      RECT 39.26 25.51 39.4 28.21 ;
      RECT 39.2 25.51 39.46 25.83 ;
      RECT 36.44 13.95 36.7 14.27 ;
      RECT 36.44 14.04 37.1 14.18 ;
      RECT 36.96 10.98 37.1 14.18 ;
      RECT 36.44 10.89 36.7 11.21 ;
      RECT 36.44 10.98 37.1 11.12 ;
      RECT 36.44 31.97 36.7 32.29 ;
      RECT 36.5 30.02 36.64 32.29 ;
      RECT 36.44 30.95 36.7 31.27 ;
      RECT 36.5 30.02 37.1 30.16 ;
      RECT 36.96 29.34 37.1 30.16 ;
      RECT 36.5 29.34 37.1 29.48 ;
      RECT 36.5 24.83 36.64 29.48 ;
      RECT 36.44 26.53 36.7 26.85 ;
      RECT 36.44 24.83 36.7 25.15 ;
      RECT 36.44 23.875 36.7 24.47 ;
      RECT 36.43 23.875 36.71 24.245 ;
      RECT 36.5 22.79 36.64 24.47 ;
      RECT 36.44 22.79 36.7 23.11 ;
      RECT 36.44 18.71 36.7 19.03 ;
      RECT 36.5 17.78 36.64 19.03 ;
      RECT 36.04 17.78 36.64 17.92 ;
      RECT 36.04 13.02 36.18 17.92 ;
      RECT 36.04 13.02 36.64 13.16 ;
      RECT 36.5 11.91 36.64 13.16 ;
      RECT 36.44 11.91 36.7 12.23 ;
      RECT 36.44 16.67 36.7 16.99 ;
      RECT 36.5 14.63 36.64 16.99 ;
      RECT 36.44 14.63 36.7 14.95 ;
      RECT 36.44 35.03 36.7 35.35 ;
      RECT 36.5 33.67 36.64 35.35 ;
      RECT 36.44 33.67 36.7 33.99 ;
      RECT 33.68 35.37 33.94 35.69 ;
      RECT 33.74 16.67 33.88 35.69 ;
      RECT 33.68 27.55 33.94 27.87 ;
      RECT 33.67 19.605 33.95 19.975 ;
      RECT 33.68 19.05 33.94 19.37 ;
      RECT 33.68 16.67 33.94 16.99 ;
      RECT 33.68 13.95 33.94 14.27 ;
      RECT 33.74 10.55 33.88 14.27 ;
      RECT 33.68 10.55 33.94 10.87 ;
      RECT 30.92 32.65 31.18 32.97 ;
      RECT 30.98 22.54 31.12 32.97 ;
      RECT 30.92 29.93 31.18 30.25 ;
      RECT 30.92 24.49 31.18 24.81 ;
      RECT 30.98 22.54 31.58 22.68 ;
      RECT 31.44 10.3 31.58 22.68 ;
      RECT 30.92 13.61 31.18 13.93 ;
      RECT 30.92 13.7 31.58 13.84 ;
      RECT 30.92 10.21 31.18 10.53 ;
      RECT 30.92 10.3 31.58 10.44 ;
      RECT 28.16 17.35 28.42 17.67 ;
      RECT 28.22 11.91 28.36 17.67 ;
      RECT 28.16 12.93 28.42 13.25 ;
      RECT 28.16 11.91 28.42 12.23 ;
      RECT 28.16 33.33 28.42 33.65 ;
      RECT 28.22 19.05 28.36 33.65 ;
      RECT 28.16 26.53 28.42 26.85 ;
      RECT 28.16 19.05 28.42 19.37 ;
      RECT 25.4 29.25 25.66 29.57 ;
      RECT 25.46 27.89 25.6 29.57 ;
      RECT 25.4 27.89 25.66 28.21 ;
      RECT 19.88 29.59 20.14 29.91 ;
      RECT 19.94 22.11 20.08 29.91 ;
      RECT 19.88 28.23 20.14 28.55 ;
      RECT 19.88 22.11 20.14 22.43 ;
      RECT 189.04 9.86 189.54 60.18 ;
      RECT 187.2 9.84 187.7 60.18 ;
      RECT 186.28 9.86 186.78 60.18 ;
      RECT 184.44 9.84 184.94 60.18 ;
      RECT 183.52 9.86 184.02 60.18 ;
      RECT 181.68 9.84 182.18 60.18 ;
      RECT 180.76 9.86 181.26 60.18 ;
      RECT 178.92 9.84 179.42 60.18 ;
      RECT 178 9.86 178.5 60.18 ;
      RECT 176.16 9.84 176.66 60.18 ;
      RECT 175.24 9.86 175.74 60.18 ;
      RECT 173.4 9.84 173.9 60.18 ;
      RECT 172.48 9.86 172.98 60.18 ;
      RECT 170.64 9.84 171.14 60.18 ;
      RECT 169.72 9.86 170.22 60.18 ;
      RECT 167.88 9.84 168.38 60.18 ;
      RECT 166.96 9.86 167.46 60.18 ;
      RECT 165.12 9.84 165.62 60.18 ;
      RECT 164.2 9.86 164.7 60.18 ;
      RECT 162.36 9.84 162.86 60.18 ;
      RECT 161.44 9.86 161.94 60.18 ;
      RECT 159.6 9.84 160.1 60.18 ;
      RECT 158.68 9.86 159.18 60.18 ;
      RECT 156.84 9.84 157.34 60.18 ;
      RECT 155.92 9.86 156.42 60.18 ;
      RECT 154.08 9.84 154.58 60.18 ;
      RECT 153.16 9.86 153.66 60.18 ;
      RECT 151.32 9.84 151.82 60.18 ;
      RECT 150.4 9.86 150.9 60.18 ;
      RECT 148.56 9.84 149.06 60.18 ;
      RECT 147.64 9.86 148.14 60.18 ;
      RECT 145.8 9.84 146.3 60.18 ;
      RECT 144.88 9.86 145.38 60.18 ;
      RECT 143.04 9.84 143.54 60.18 ;
      RECT 142.12 9.86 142.62 60.18 ;
      RECT 141.31 24.485 141.59 24.855 ;
      RECT 140.28 9.84 140.78 60.18 ;
      RECT 139.36 9.86 139.86 60.18 ;
      RECT 137.52 9.84 138.02 60.18 ;
      RECT 136.6 9.86 137.1 60.18 ;
      RECT 134.76 9.84 135.26 60.18 ;
      RECT 133.84 9.86 134.34 60.18 ;
      RECT 132 9.84 132.5 60.18 ;
      RECT 131.08 9.86 131.58 60.18 ;
      RECT 129.24 9.84 129.74 60.18 ;
      RECT 128.32 9.86 128.82 60.18 ;
      RECT 126.48 9.84 126.98 60.18 ;
      RECT 125.56 9.86 126.06 60.18 ;
      RECT 123.72 9.84 124.22 60.18 ;
      RECT 122.8 9.86 123.3 60.18 ;
      RECT 120.96 9.84 121.46 60.18 ;
      RECT 120.04 9.86 120.54 60.18 ;
      RECT 118.2 9.84 118.7 60.18 ;
      RECT 117.28 9.86 117.78 60.18 ;
      RECT 115.44 9.84 115.94 60.18 ;
      RECT 114.52 9.86 115.02 60.18 ;
      RECT 112.68 9.84 113.18 60.18 ;
      RECT 111.76 9.86 112.26 60.18 ;
      RECT 109.92 9.84 110.42 60.18 ;
      RECT 109 9.86 109.5 60.18 ;
      RECT 107.16 9.84 107.66 60.18 ;
      RECT 106.24 9.86 106.74 60.18 ;
      RECT 104.4 9.84 104.9 60.18 ;
      RECT 103.48 9.86 103.98 60.18 ;
      RECT 101.64 9.84 102.14 60.18 ;
      RECT 100.72 9.86 101.22 60.18 ;
      RECT 98.88 9.84 99.38 60.18 ;
      RECT 97.96 9.86 98.46 60.18 ;
      RECT 96.12 9.84 96.62 60.18 ;
      RECT 95.2 9.86 95.7 60.18 ;
      RECT 93.36 9.84 93.86 60.18 ;
      RECT 92.44 9.86 92.94 60.18 ;
      RECT 90.6 9.84 91.1 60.18 ;
      RECT 89.68 9.86 90.18 60.18 ;
      RECT 87.84 9.84 88.34 60.18 ;
      RECT 86.92 9.86 87.42 60.18 ;
      RECT 85.08 9.84 85.58 60.18 ;
      RECT 84.16 9.86 84.66 60.18 ;
      RECT 82.32 9.84 82.82 60.18 ;
      RECT 81.4 9.86 81.9 60.18 ;
      RECT 79.56 9.84 80.06 60.18 ;
      RECT 78.64 9.86 79.14 60.18 ;
      RECT 77.83 24.485 78.11 24.855 ;
      RECT 76.8 9.84 77.3 60.18 ;
      RECT 75.88 9.86 76.38 60.18 ;
      RECT 74.04 9.84 74.54 60.18 ;
      RECT 73.12 9.86 73.62 60.18 ;
      RECT 71.28 9.84 71.78 60.18 ;
      RECT 70.36 9.86 70.86 60.18 ;
      RECT 68.52 9.84 69.02 60.18 ;
      RECT 67.6 9.86 68.1 60.18 ;
      RECT 65.76 9.84 66.26 60.18 ;
      RECT 64.84 9.86 65.34 60.18 ;
      RECT 63 9.84 63.5 60.18 ;
      RECT 62.08 9.86 62.58 60.18 ;
      RECT 60.24 9.84 60.74 60.18 ;
      RECT 59.32 9.86 59.82 60.18 ;
      RECT 57.48 9.84 57.98 60.18 ;
      RECT 56.56 9.86 57.06 60.18 ;
      RECT 54.72 9.84 55.22 60.18 ;
      RECT 53.8 9.86 54.3 60.18 ;
      RECT 51.96 9.84 52.46 60.18 ;
      RECT 51.04 9.86 51.54 60.18 ;
      RECT 49.2 9.84 49.7 60.18 ;
      RECT 48.28 9.86 48.78 60.18 ;
      RECT 46.44 9.84 46.94 60.18 ;
      RECT 45.52 9.86 46.02 60.18 ;
      RECT 43.68 9.84 44.18 60.18 ;
      RECT 42.76 9.86 43.26 60.18 ;
      RECT 40.92 9.84 41.42 60.18 ;
      RECT 40 9.86 40.5 60.18 ;
      RECT 38.16 9.84 38.66 60.18 ;
      RECT 37.24 9.86 37.74 60.18 ;
      RECT 35.4 9.84 35.9 60.18 ;
      RECT 34.48 9.86 34.98 60.18 ;
      RECT 32.64 9.84 33.14 60.18 ;
      RECT 31.72 9.86 32.22 60.18 ;
      RECT 29.88 9.84 30.38 60.18 ;
      RECT 28.96 9.86 29.46 60.18 ;
      RECT 27.12 9.84 27.62 60.18 ;
      RECT 26.2 9.86 26.7 60.18 ;
      RECT 24.36 9.84 24.86 60.18 ;
      RECT 23.44 9.86 23.94 60.18 ;
      RECT 21.6 9.84 22.1 60.18 ;
      RECT 20.68 9.86 21.18 60.18 ;
      RECT 18.84 9.84 19.34 60.18 ;
      RECT 17.92 9.86 18.42 60.18 ;
      RECT 16.08 9.84 16.58 60.18 ;
      RECT 15.16 9.86 15.66 60.18 ;
    LAYER via2 ;
      RECT 189.19 17.58 189.39 17.78 ;
      RECT 189.19 21.66 189.39 21.86 ;
      RECT 189.19 25.74 189.39 25.94 ;
      RECT 189.19 29.82 189.39 30.02 ;
      RECT 189.19 33.9 189.39 34.1 ;
      RECT 189.19 37.98 189.39 38.18 ;
      RECT 189.19 42.06 189.39 42.26 ;
      RECT 189.19 46.14 189.39 46.34 ;
      RECT 189.19 50.22 189.39 50.42 ;
      RECT 189.19 54.3 189.39 54.5 ;
      RECT 189.19 58.38 189.39 58.58 ;
      RECT 187.35 18.94 187.55 19.14 ;
      RECT 187.35 23.02 187.55 23.22 ;
      RECT 187.35 27.1 187.55 27.3 ;
      RECT 187.35 31.18 187.55 31.38 ;
      RECT 187.35 35.26 187.55 35.46 ;
      RECT 187.35 39.34 187.55 39.54 ;
      RECT 187.35 43.42 187.55 43.62 ;
      RECT 187.35 47.5 187.55 47.7 ;
      RECT 187.35 51.58 187.55 51.78 ;
      RECT 187.35 55.66 187.55 55.86 ;
      RECT 187.35 59.74 187.55 59.94 ;
      RECT 186.43 17.58 186.63 17.78 ;
      RECT 186.43 21.66 186.63 21.86 ;
      RECT 186.43 25.74 186.63 25.94 ;
      RECT 186.43 29.82 186.63 30.02 ;
      RECT 186.43 33.9 186.63 34.1 ;
      RECT 186.43 37.98 186.63 38.18 ;
      RECT 186.43 42.06 186.63 42.26 ;
      RECT 186.43 46.14 186.63 46.34 ;
      RECT 186.43 50.22 186.63 50.42 ;
      RECT 186.43 54.3 186.63 54.5 ;
      RECT 186.43 58.38 186.63 58.58 ;
      RECT 184.59 18.94 184.79 19.14 ;
      RECT 184.59 23.02 184.79 23.22 ;
      RECT 184.59 27.1 184.79 27.3 ;
      RECT 184.59 31.18 184.79 31.38 ;
      RECT 184.59 35.26 184.79 35.46 ;
      RECT 184.59 39.34 184.79 39.54 ;
      RECT 184.59 43.42 184.79 43.62 ;
      RECT 184.59 47.5 184.79 47.7 ;
      RECT 184.59 51.58 184.79 51.78 ;
      RECT 184.59 55.66 184.79 55.86 ;
      RECT 184.59 59.74 184.79 59.94 ;
      RECT 183.67 17.58 183.87 17.78 ;
      RECT 183.67 21.66 183.87 21.86 ;
      RECT 183.67 25.74 183.87 25.94 ;
      RECT 183.67 29.82 183.87 30.02 ;
      RECT 183.67 33.9 183.87 34.1 ;
      RECT 183.67 37.98 183.87 38.18 ;
      RECT 183.67 42.06 183.87 42.26 ;
      RECT 183.67 46.14 183.87 46.34 ;
      RECT 183.67 50.22 183.87 50.42 ;
      RECT 183.67 54.3 183.87 54.5 ;
      RECT 183.67 58.38 183.87 58.58 ;
      RECT 181.83 18.94 182.03 19.14 ;
      RECT 181.83 23.02 182.03 23.22 ;
      RECT 181.83 27.1 182.03 27.3 ;
      RECT 181.83 31.18 182.03 31.38 ;
      RECT 181.83 35.26 182.03 35.46 ;
      RECT 181.83 39.34 182.03 39.54 ;
      RECT 181.83 43.42 182.03 43.62 ;
      RECT 181.83 47.5 182.03 47.7 ;
      RECT 181.83 51.58 182.03 51.78 ;
      RECT 181.83 55.66 182.03 55.86 ;
      RECT 181.83 59.74 182.03 59.94 ;
      RECT 180.91 17.58 181.11 17.78 ;
      RECT 180.91 21.66 181.11 21.86 ;
      RECT 180.91 25.74 181.11 25.94 ;
      RECT 180.91 29.82 181.11 30.02 ;
      RECT 180.91 33.9 181.11 34.1 ;
      RECT 180.91 37.98 181.11 38.18 ;
      RECT 180.91 42.06 181.11 42.26 ;
      RECT 180.91 46.14 181.11 46.34 ;
      RECT 180.91 50.22 181.11 50.42 ;
      RECT 180.91 54.3 181.11 54.5 ;
      RECT 180.91 58.38 181.11 58.58 ;
      RECT 179.07 18.94 179.27 19.14 ;
      RECT 179.07 23.02 179.27 23.22 ;
      RECT 179.07 27.1 179.27 27.3 ;
      RECT 179.07 31.18 179.27 31.38 ;
      RECT 179.07 35.26 179.27 35.46 ;
      RECT 179.07 39.34 179.27 39.54 ;
      RECT 179.07 43.42 179.27 43.62 ;
      RECT 179.07 47.5 179.27 47.7 ;
      RECT 179.07 51.58 179.27 51.78 ;
      RECT 179.07 55.66 179.27 55.86 ;
      RECT 179.07 59.74 179.27 59.94 ;
      RECT 178.15 17.58 178.35 17.78 ;
      RECT 178.15 21.66 178.35 21.86 ;
      RECT 178.15 25.74 178.35 25.94 ;
      RECT 178.15 29.82 178.35 30.02 ;
      RECT 178.15 33.9 178.35 34.1 ;
      RECT 178.15 37.98 178.35 38.18 ;
      RECT 178.15 42.06 178.35 42.26 ;
      RECT 178.15 46.14 178.35 46.34 ;
      RECT 178.15 50.22 178.35 50.42 ;
      RECT 178.15 54.3 178.35 54.5 ;
      RECT 178.15 58.38 178.35 58.58 ;
      RECT 177.23 15.42 177.43 15.62 ;
      RECT 176.31 18.94 176.51 19.14 ;
      RECT 176.31 23.02 176.51 23.22 ;
      RECT 176.31 27.1 176.51 27.3 ;
      RECT 176.31 31.18 176.51 31.38 ;
      RECT 176.31 35.26 176.51 35.46 ;
      RECT 176.31 39.34 176.51 39.54 ;
      RECT 176.31 43.42 176.51 43.62 ;
      RECT 176.31 47.5 176.51 47.7 ;
      RECT 176.31 51.58 176.51 51.78 ;
      RECT 176.31 55.66 176.51 55.86 ;
      RECT 176.31 59.74 176.51 59.94 ;
      RECT 175.39 17.58 175.59 17.78 ;
      RECT 175.39 21.66 175.59 21.86 ;
      RECT 175.39 25.74 175.59 25.94 ;
      RECT 175.39 29.82 175.59 30.02 ;
      RECT 175.39 33.9 175.59 34.1 ;
      RECT 175.39 37.98 175.59 38.18 ;
      RECT 175.39 42.06 175.59 42.26 ;
      RECT 175.39 46.14 175.59 46.34 ;
      RECT 175.39 50.22 175.59 50.42 ;
      RECT 175.39 54.3 175.59 54.5 ;
      RECT 175.39 58.38 175.59 58.58 ;
      RECT 173.55 18.94 173.75 19.14 ;
      RECT 173.55 23.02 173.75 23.22 ;
      RECT 173.55 27.1 173.75 27.3 ;
      RECT 173.55 31.18 173.75 31.38 ;
      RECT 173.55 35.26 173.75 35.46 ;
      RECT 173.55 39.34 173.75 39.54 ;
      RECT 173.55 43.42 173.75 43.62 ;
      RECT 173.55 47.5 173.75 47.7 ;
      RECT 173.55 51.58 173.75 51.78 ;
      RECT 173.55 55.66 173.75 55.86 ;
      RECT 173.55 59.74 173.75 59.94 ;
      RECT 172.63 17.58 172.83 17.78 ;
      RECT 172.63 21.66 172.83 21.86 ;
      RECT 172.63 25.74 172.83 25.94 ;
      RECT 172.63 29.82 172.83 30.02 ;
      RECT 172.63 33.9 172.83 34.1 ;
      RECT 172.63 37.98 172.83 38.18 ;
      RECT 172.63 42.06 172.83 42.26 ;
      RECT 172.63 46.14 172.83 46.34 ;
      RECT 172.63 50.22 172.83 50.42 ;
      RECT 172.63 54.3 172.83 54.5 ;
      RECT 172.63 58.38 172.83 58.58 ;
      RECT 170.79 18.94 170.99 19.14 ;
      RECT 170.79 23.02 170.99 23.22 ;
      RECT 170.79 27.1 170.99 27.3 ;
      RECT 170.79 31.18 170.99 31.38 ;
      RECT 170.79 35.26 170.99 35.46 ;
      RECT 170.79 39.34 170.99 39.54 ;
      RECT 170.79 43.42 170.99 43.62 ;
      RECT 170.79 47.5 170.99 47.7 ;
      RECT 170.79 51.58 170.99 51.78 ;
      RECT 170.79 55.66 170.99 55.86 ;
      RECT 170.79 59.74 170.99 59.94 ;
      RECT 169.87 17.58 170.07 17.78 ;
      RECT 169.87 21.66 170.07 21.86 ;
      RECT 169.87 25.74 170.07 25.94 ;
      RECT 169.87 29.82 170.07 30.02 ;
      RECT 169.87 33.9 170.07 34.1 ;
      RECT 169.87 37.98 170.07 38.18 ;
      RECT 169.87 42.06 170.07 42.26 ;
      RECT 169.87 46.14 170.07 46.34 ;
      RECT 169.87 50.22 170.07 50.42 ;
      RECT 169.87 54.3 170.07 54.5 ;
      RECT 169.87 58.38 170.07 58.58 ;
      RECT 168.95 9.32 169.15 9.52 ;
      RECT 168.03 18.94 168.23 19.14 ;
      RECT 168.03 23.02 168.23 23.22 ;
      RECT 168.03 27.1 168.23 27.3 ;
      RECT 168.03 31.18 168.23 31.38 ;
      RECT 168.03 35.26 168.23 35.46 ;
      RECT 168.03 39.34 168.23 39.54 ;
      RECT 168.03 43.42 168.23 43.62 ;
      RECT 168.03 47.5 168.23 47.7 ;
      RECT 168.03 51.58 168.23 51.78 ;
      RECT 168.03 55.66 168.23 55.86 ;
      RECT 168.03 59.74 168.23 59.94 ;
      RECT 167.11 17.58 167.31 17.78 ;
      RECT 167.11 21.66 167.31 21.86 ;
      RECT 167.11 25.74 167.31 25.94 ;
      RECT 167.11 29.82 167.31 30.02 ;
      RECT 167.11 33.9 167.31 34.1 ;
      RECT 167.11 37.98 167.31 38.18 ;
      RECT 167.11 42.06 167.31 42.26 ;
      RECT 167.11 46.14 167.31 46.34 ;
      RECT 167.11 50.22 167.31 50.42 ;
      RECT 167.11 54.3 167.31 54.5 ;
      RECT 167.11 58.38 167.31 58.58 ;
      RECT 165.27 18.94 165.47 19.14 ;
      RECT 165.27 23.02 165.47 23.22 ;
      RECT 165.27 27.1 165.47 27.3 ;
      RECT 165.27 31.18 165.47 31.38 ;
      RECT 165.27 35.26 165.47 35.46 ;
      RECT 165.27 39.34 165.47 39.54 ;
      RECT 165.27 43.42 165.47 43.62 ;
      RECT 165.27 47.5 165.47 47.7 ;
      RECT 165.27 51.58 165.47 51.78 ;
      RECT 165.27 55.66 165.47 55.86 ;
      RECT 165.27 59.74 165.47 59.94 ;
      RECT 164.35 17.58 164.55 17.78 ;
      RECT 164.35 21.66 164.55 21.86 ;
      RECT 164.35 25.74 164.55 25.94 ;
      RECT 164.35 29.82 164.55 30.02 ;
      RECT 164.35 33.9 164.55 34.1 ;
      RECT 164.35 37.98 164.55 38.18 ;
      RECT 164.35 42.06 164.55 42.26 ;
      RECT 164.35 46.14 164.55 46.34 ;
      RECT 164.35 50.22 164.55 50.42 ;
      RECT 164.35 54.3 164.55 54.5 ;
      RECT 164.35 58.38 164.55 58.58 ;
      RECT 162.51 18.94 162.71 19.14 ;
      RECT 162.51 23.02 162.71 23.22 ;
      RECT 162.51 27.1 162.71 27.3 ;
      RECT 162.51 31.18 162.71 31.38 ;
      RECT 162.51 35.26 162.71 35.46 ;
      RECT 162.51 39.34 162.71 39.54 ;
      RECT 162.51 43.42 162.71 43.62 ;
      RECT 162.51 47.5 162.71 47.7 ;
      RECT 162.51 51.58 162.71 51.78 ;
      RECT 162.51 55.66 162.71 55.86 ;
      RECT 162.51 59.74 162.71 59.94 ;
      RECT 161.59 17.58 161.79 17.78 ;
      RECT 161.59 21.66 161.79 21.86 ;
      RECT 161.59 25.74 161.79 25.94 ;
      RECT 161.59 29.82 161.79 30.02 ;
      RECT 161.59 33.9 161.79 34.1 ;
      RECT 161.59 37.98 161.79 38.18 ;
      RECT 161.59 42.06 161.79 42.26 ;
      RECT 161.59 46.14 161.79 46.34 ;
      RECT 161.59 50.22 161.79 50.42 ;
      RECT 161.59 54.3 161.79 54.5 ;
      RECT 161.59 58.38 161.79 58.58 ;
      RECT 160.67 16.64 160.87 16.84 ;
      RECT 160.67 19.69 160.87 19.89 ;
      RECT 159.75 18.94 159.95 19.14 ;
      RECT 159.75 23.02 159.95 23.22 ;
      RECT 159.75 27.1 159.95 27.3 ;
      RECT 159.75 31.18 159.95 31.38 ;
      RECT 159.75 35.26 159.95 35.46 ;
      RECT 159.75 39.34 159.95 39.54 ;
      RECT 159.75 43.42 159.95 43.62 ;
      RECT 159.75 47.5 159.95 47.7 ;
      RECT 159.75 51.58 159.95 51.78 ;
      RECT 159.75 55.66 159.95 55.86 ;
      RECT 159.75 59.74 159.95 59.94 ;
      RECT 158.83 17.58 159.03 17.78 ;
      RECT 158.83 21.66 159.03 21.86 ;
      RECT 158.83 25.74 159.03 25.94 ;
      RECT 158.83 29.82 159.03 30.02 ;
      RECT 158.83 33.9 159.03 34.1 ;
      RECT 158.83 37.98 159.03 38.18 ;
      RECT 158.83 42.06 159.03 42.26 ;
      RECT 158.83 46.14 159.03 46.34 ;
      RECT 158.83 50.22 159.03 50.42 ;
      RECT 158.83 54.3 159.03 54.5 ;
      RECT 158.83 58.38 159.03 58.58 ;
      RECT 157.91 15.42 158.11 15.62 ;
      RECT 156.99 18.94 157.19 19.14 ;
      RECT 156.99 23.02 157.19 23.22 ;
      RECT 156.99 27.1 157.19 27.3 ;
      RECT 156.99 31.18 157.19 31.38 ;
      RECT 156.99 35.26 157.19 35.46 ;
      RECT 156.99 39.34 157.19 39.54 ;
      RECT 156.99 43.42 157.19 43.62 ;
      RECT 156.99 47.5 157.19 47.7 ;
      RECT 156.99 51.58 157.19 51.78 ;
      RECT 156.99 55.66 157.19 55.86 ;
      RECT 156.99 59.74 157.19 59.94 ;
      RECT 156.07 17.58 156.27 17.78 ;
      RECT 156.07 21.66 156.27 21.86 ;
      RECT 156.07 25.74 156.27 25.94 ;
      RECT 156.07 29.82 156.27 30.02 ;
      RECT 156.07 33.9 156.27 34.1 ;
      RECT 156.07 37.98 156.27 38.18 ;
      RECT 156.07 42.06 156.27 42.26 ;
      RECT 156.07 46.14 156.27 46.34 ;
      RECT 156.07 50.22 156.27 50.42 ;
      RECT 156.07 54.3 156.27 54.5 ;
      RECT 156.07 58.38 156.27 58.58 ;
      RECT 154.23 18.94 154.43 19.14 ;
      RECT 154.23 23.02 154.43 23.22 ;
      RECT 154.23 27.1 154.43 27.3 ;
      RECT 154.23 31.18 154.43 31.38 ;
      RECT 154.23 35.26 154.43 35.46 ;
      RECT 154.23 39.34 154.43 39.54 ;
      RECT 154.23 43.42 154.43 43.62 ;
      RECT 154.23 47.5 154.43 47.7 ;
      RECT 154.23 51.58 154.43 51.78 ;
      RECT 154.23 55.66 154.43 55.86 ;
      RECT 154.23 59.74 154.43 59.94 ;
      RECT 153.31 17.58 153.51 17.78 ;
      RECT 153.31 21.66 153.51 21.86 ;
      RECT 153.31 25.74 153.51 25.94 ;
      RECT 153.31 29.82 153.51 30.02 ;
      RECT 153.31 33.9 153.51 34.1 ;
      RECT 153.31 37.98 153.51 38.18 ;
      RECT 153.31 42.06 153.51 42.26 ;
      RECT 153.31 46.14 153.51 46.34 ;
      RECT 153.31 50.22 153.51 50.42 ;
      RECT 153.31 54.3 153.51 54.5 ;
      RECT 153.31 58.38 153.51 58.58 ;
      RECT 151.47 18.94 151.67 19.14 ;
      RECT 151.47 23.02 151.67 23.22 ;
      RECT 151.47 27.1 151.67 27.3 ;
      RECT 151.47 31.18 151.67 31.38 ;
      RECT 151.47 35.26 151.67 35.46 ;
      RECT 151.47 39.34 151.67 39.54 ;
      RECT 151.47 43.42 151.67 43.62 ;
      RECT 151.47 47.5 151.67 47.7 ;
      RECT 151.47 51.58 151.67 51.78 ;
      RECT 151.47 55.66 151.67 55.86 ;
      RECT 151.47 59.74 151.67 59.94 ;
      RECT 150.55 17.58 150.75 17.78 ;
      RECT 150.55 21.66 150.75 21.86 ;
      RECT 150.55 25.74 150.75 25.94 ;
      RECT 150.55 29.82 150.75 30.02 ;
      RECT 150.55 33.9 150.75 34.1 ;
      RECT 150.55 37.98 150.75 38.18 ;
      RECT 150.55 42.06 150.75 42.26 ;
      RECT 150.55 46.14 150.75 46.34 ;
      RECT 150.55 50.22 150.75 50.42 ;
      RECT 150.55 54.3 150.75 54.5 ;
      RECT 150.55 58.38 150.75 58.58 ;
      RECT 150.09 9.32 150.29 9.52 ;
      RECT 149.63 24.57 149.83 24.77 ;
      RECT 148.71 18.94 148.91 19.14 ;
      RECT 148.71 23.02 148.91 23.22 ;
      RECT 148.71 27.1 148.91 27.3 ;
      RECT 148.71 31.18 148.91 31.38 ;
      RECT 148.71 35.26 148.91 35.46 ;
      RECT 148.71 39.34 148.91 39.54 ;
      RECT 148.71 43.42 148.91 43.62 ;
      RECT 148.71 47.5 148.91 47.7 ;
      RECT 148.71 51.58 148.91 51.78 ;
      RECT 148.71 55.66 148.91 55.86 ;
      RECT 148.71 59.74 148.91 59.94 ;
      RECT 147.79 17.58 147.99 17.78 ;
      RECT 147.79 21.66 147.99 21.86 ;
      RECT 147.79 25.74 147.99 25.94 ;
      RECT 147.79 29.82 147.99 30.02 ;
      RECT 147.79 33.9 147.99 34.1 ;
      RECT 147.79 37.98 147.99 38.18 ;
      RECT 147.79 42.06 147.99 42.26 ;
      RECT 147.79 46.14 147.99 46.34 ;
      RECT 147.79 50.22 147.99 50.42 ;
      RECT 147.79 54.3 147.99 54.5 ;
      RECT 147.79 58.38 147.99 58.58 ;
      RECT 145.95 18.94 146.15 19.14 ;
      RECT 145.95 23.02 146.15 23.22 ;
      RECT 145.95 27.1 146.15 27.3 ;
      RECT 145.95 31.18 146.15 31.38 ;
      RECT 145.95 35.26 146.15 35.46 ;
      RECT 145.95 39.34 146.15 39.54 ;
      RECT 145.95 43.42 146.15 43.62 ;
      RECT 145.95 47.5 146.15 47.7 ;
      RECT 145.95 51.58 146.15 51.78 ;
      RECT 145.95 55.66 146.15 55.86 ;
      RECT 145.95 59.74 146.15 59.94 ;
      RECT 145.03 17.58 145.23 17.78 ;
      RECT 145.03 21.66 145.23 21.86 ;
      RECT 145.03 25.74 145.23 25.94 ;
      RECT 145.03 29.82 145.23 30.02 ;
      RECT 145.03 33.9 145.23 34.1 ;
      RECT 145.03 37.98 145.23 38.18 ;
      RECT 145.03 42.06 145.23 42.26 ;
      RECT 145.03 46.14 145.23 46.34 ;
      RECT 145.03 50.22 145.23 50.42 ;
      RECT 145.03 54.3 145.23 54.5 ;
      RECT 145.03 58.38 145.23 58.58 ;
      RECT 143.19 18.94 143.39 19.14 ;
      RECT 143.19 23.02 143.39 23.22 ;
      RECT 143.19 27.1 143.39 27.3 ;
      RECT 143.19 31.18 143.39 31.38 ;
      RECT 143.19 35.26 143.39 35.46 ;
      RECT 143.19 39.34 143.39 39.54 ;
      RECT 143.19 43.42 143.39 43.62 ;
      RECT 143.19 47.5 143.39 47.7 ;
      RECT 143.19 51.58 143.39 51.78 ;
      RECT 143.19 55.66 143.39 55.86 ;
      RECT 143.19 59.74 143.39 59.94 ;
      RECT 142.27 17.58 142.47 17.78 ;
      RECT 142.27 21.66 142.47 21.86 ;
      RECT 142.27 25.74 142.47 25.94 ;
      RECT 142.27 29.82 142.47 30.02 ;
      RECT 142.27 33.9 142.47 34.1 ;
      RECT 142.27 37.98 142.47 38.18 ;
      RECT 142.27 42.06 142.47 42.26 ;
      RECT 142.27 46.14 142.47 46.34 ;
      RECT 142.27 50.22 142.47 50.42 ;
      RECT 142.27 54.3 142.47 54.5 ;
      RECT 142.27 58.38 142.47 58.58 ;
      RECT 141.35 20.91 141.55 21.11 ;
      RECT 141.35 24.57 141.55 24.77 ;
      RECT 140.43 18.94 140.63 19.14 ;
      RECT 140.43 23.02 140.63 23.22 ;
      RECT 140.43 27.1 140.63 27.3 ;
      RECT 140.43 31.18 140.63 31.38 ;
      RECT 140.43 35.26 140.63 35.46 ;
      RECT 140.43 39.34 140.63 39.54 ;
      RECT 140.43 43.42 140.63 43.62 ;
      RECT 140.43 47.5 140.63 47.7 ;
      RECT 140.43 51.58 140.63 51.78 ;
      RECT 140.43 55.66 140.63 55.86 ;
      RECT 140.43 59.74 140.63 59.94 ;
      RECT 139.51 17.58 139.71 17.78 ;
      RECT 139.51 21.66 139.71 21.86 ;
      RECT 139.51 25.74 139.71 25.94 ;
      RECT 139.51 29.82 139.71 30.02 ;
      RECT 139.51 33.9 139.71 34.1 ;
      RECT 139.51 37.98 139.71 38.18 ;
      RECT 139.51 42.06 139.71 42.26 ;
      RECT 139.51 46.14 139.71 46.34 ;
      RECT 139.51 50.22 139.71 50.42 ;
      RECT 139.51 54.3 139.71 54.5 ;
      RECT 139.51 58.38 139.71 58.58 ;
      RECT 138.59 16.64 138.79 16.84 ;
      RECT 137.67 18.94 137.87 19.14 ;
      RECT 137.67 23.02 137.87 23.22 ;
      RECT 137.67 27.1 137.87 27.3 ;
      RECT 137.67 31.18 137.87 31.38 ;
      RECT 137.67 35.26 137.87 35.46 ;
      RECT 137.67 39.34 137.87 39.54 ;
      RECT 137.67 43.42 137.87 43.62 ;
      RECT 137.67 47.5 137.87 47.7 ;
      RECT 137.67 51.58 137.87 51.78 ;
      RECT 137.67 55.66 137.87 55.86 ;
      RECT 137.67 59.74 137.87 59.94 ;
      RECT 136.75 17.58 136.95 17.78 ;
      RECT 136.75 21.66 136.95 21.86 ;
      RECT 136.75 25.74 136.95 25.94 ;
      RECT 136.75 29.82 136.95 30.02 ;
      RECT 136.75 33.9 136.95 34.1 ;
      RECT 136.75 37.98 136.95 38.18 ;
      RECT 136.75 42.06 136.95 42.26 ;
      RECT 136.75 46.14 136.95 46.34 ;
      RECT 136.75 50.22 136.95 50.42 ;
      RECT 136.75 54.3 136.95 54.5 ;
      RECT 136.75 58.38 136.95 58.58 ;
      RECT 135.83 23.96 136.03 24.16 ;
      RECT 134.91 18.94 135.11 19.14 ;
      RECT 134.91 23.02 135.11 23.22 ;
      RECT 134.91 27.1 135.11 27.3 ;
      RECT 134.91 31.18 135.11 31.38 ;
      RECT 134.91 35.26 135.11 35.46 ;
      RECT 134.91 39.34 135.11 39.54 ;
      RECT 134.91 43.42 135.11 43.62 ;
      RECT 134.91 47.5 135.11 47.7 ;
      RECT 134.91 51.58 135.11 51.78 ;
      RECT 134.91 55.66 135.11 55.86 ;
      RECT 134.91 59.74 135.11 59.94 ;
      RECT 133.99 17.58 134.19 17.78 ;
      RECT 133.99 21.66 134.19 21.86 ;
      RECT 133.99 25.74 134.19 25.94 ;
      RECT 133.99 29.82 134.19 30.02 ;
      RECT 133.99 33.9 134.19 34.1 ;
      RECT 133.99 37.98 134.19 38.18 ;
      RECT 133.99 42.06 134.19 42.26 ;
      RECT 133.99 46.14 134.19 46.34 ;
      RECT 133.99 50.22 134.19 50.42 ;
      RECT 133.99 54.3 134.19 54.5 ;
      RECT 133.99 58.38 134.19 58.58 ;
      RECT 133.07 19.69 133.27 19.89 ;
      RECT 133.07 20.91 133.27 21.11 ;
      RECT 133.07 28.84 133.27 29.04 ;
      RECT 132.15 18.94 132.35 19.14 ;
      RECT 132.15 23.02 132.35 23.22 ;
      RECT 132.15 27.1 132.35 27.3 ;
      RECT 132.15 31.18 132.35 31.38 ;
      RECT 132.15 35.26 132.35 35.46 ;
      RECT 132.15 39.34 132.35 39.54 ;
      RECT 132.15 43.42 132.35 43.62 ;
      RECT 132.15 47.5 132.35 47.7 ;
      RECT 132.15 51.58 132.35 51.78 ;
      RECT 132.15 55.66 132.35 55.86 ;
      RECT 132.15 59.74 132.35 59.94 ;
      RECT 131.23 17.58 131.43 17.78 ;
      RECT 131.23 21.66 131.43 21.86 ;
      RECT 131.23 25.74 131.43 25.94 ;
      RECT 131.23 29.82 131.43 30.02 ;
      RECT 131.23 33.9 131.43 34.1 ;
      RECT 131.23 37.98 131.43 38.18 ;
      RECT 131.23 42.06 131.43 42.26 ;
      RECT 131.23 46.14 131.43 46.34 ;
      RECT 131.23 50.22 131.43 50.42 ;
      RECT 131.23 54.3 131.43 54.5 ;
      RECT 131.23 58.38 131.43 58.58 ;
      RECT 129.39 18.94 129.59 19.14 ;
      RECT 129.39 23.02 129.59 23.22 ;
      RECT 129.39 27.1 129.59 27.3 ;
      RECT 129.39 31.18 129.59 31.38 ;
      RECT 129.39 35.26 129.59 35.46 ;
      RECT 129.39 39.34 129.59 39.54 ;
      RECT 129.39 43.42 129.59 43.62 ;
      RECT 129.39 47.5 129.59 47.7 ;
      RECT 129.39 51.58 129.59 51.78 ;
      RECT 129.39 55.66 129.59 55.86 ;
      RECT 129.39 59.74 129.59 59.94 ;
      RECT 128.47 17.58 128.67 17.78 ;
      RECT 128.47 21.66 128.67 21.86 ;
      RECT 128.47 25.74 128.67 25.94 ;
      RECT 128.47 29.82 128.67 30.02 ;
      RECT 128.47 33.9 128.67 34.1 ;
      RECT 128.47 37.98 128.67 38.18 ;
      RECT 128.47 42.06 128.67 42.26 ;
      RECT 128.47 46.14 128.67 46.34 ;
      RECT 128.47 50.22 128.67 50.42 ;
      RECT 128.47 54.3 128.67 54.5 ;
      RECT 128.47 58.38 128.67 58.58 ;
      RECT 127.55 20.91 127.75 21.11 ;
      RECT 127.55 28.23 127.75 28.43 ;
      RECT 126.63 18.94 126.83 19.14 ;
      RECT 126.63 23.02 126.83 23.22 ;
      RECT 126.63 27.1 126.83 27.3 ;
      RECT 126.63 31.18 126.83 31.38 ;
      RECT 126.63 35.26 126.83 35.46 ;
      RECT 126.63 39.34 126.83 39.54 ;
      RECT 126.63 43.42 126.83 43.62 ;
      RECT 126.63 47.5 126.83 47.7 ;
      RECT 126.63 51.58 126.83 51.78 ;
      RECT 126.63 55.66 126.83 55.86 ;
      RECT 126.63 59.74 126.83 59.94 ;
      RECT 125.71 17.58 125.91 17.78 ;
      RECT 125.71 21.66 125.91 21.86 ;
      RECT 125.71 25.74 125.91 25.94 ;
      RECT 125.71 29.82 125.91 30.02 ;
      RECT 125.71 33.9 125.91 34.1 ;
      RECT 125.71 37.98 125.91 38.18 ;
      RECT 125.71 42.06 125.91 42.26 ;
      RECT 125.71 46.14 125.91 46.34 ;
      RECT 125.71 50.22 125.91 50.42 ;
      RECT 125.71 54.3 125.91 54.5 ;
      RECT 125.71 58.38 125.91 58.58 ;
      RECT 124.79 15.42 124.99 15.62 ;
      RECT 124.79 16.64 124.99 16.84 ;
      RECT 123.87 18.94 124.07 19.14 ;
      RECT 123.87 23.02 124.07 23.22 ;
      RECT 123.87 27.1 124.07 27.3 ;
      RECT 123.87 31.18 124.07 31.38 ;
      RECT 123.87 35.26 124.07 35.46 ;
      RECT 123.87 39.34 124.07 39.54 ;
      RECT 123.87 43.42 124.07 43.62 ;
      RECT 123.87 47.5 124.07 47.7 ;
      RECT 123.87 51.58 124.07 51.78 ;
      RECT 123.87 55.66 124.07 55.86 ;
      RECT 123.87 59.74 124.07 59.94 ;
      RECT 122.95 17.58 123.15 17.78 ;
      RECT 122.95 21.66 123.15 21.86 ;
      RECT 122.95 25.74 123.15 25.94 ;
      RECT 122.95 29.82 123.15 30.02 ;
      RECT 122.95 33.9 123.15 34.1 ;
      RECT 122.95 37.98 123.15 38.18 ;
      RECT 122.95 42.06 123.15 42.26 ;
      RECT 122.95 46.14 123.15 46.34 ;
      RECT 122.95 50.22 123.15 50.42 ;
      RECT 122.95 54.3 123.15 54.5 ;
      RECT 122.95 58.38 123.15 58.58 ;
      RECT 122.03 14.2 122.23 14.4 ;
      RECT 122.03 23.96 122.23 24.16 ;
      RECT 121.11 18.94 121.31 19.14 ;
      RECT 121.11 23.02 121.31 23.22 ;
      RECT 121.11 27.1 121.31 27.3 ;
      RECT 121.11 31.18 121.31 31.38 ;
      RECT 121.11 35.26 121.31 35.46 ;
      RECT 121.11 39.34 121.31 39.54 ;
      RECT 121.11 43.42 121.31 43.62 ;
      RECT 121.11 47.5 121.31 47.7 ;
      RECT 121.11 51.58 121.31 51.78 ;
      RECT 121.11 55.66 121.31 55.86 ;
      RECT 121.11 59.74 121.31 59.94 ;
      RECT 120.19 17.58 120.39 17.78 ;
      RECT 120.19 21.66 120.39 21.86 ;
      RECT 120.19 25.74 120.39 25.94 ;
      RECT 120.19 29.82 120.39 30.02 ;
      RECT 120.19 33.9 120.39 34.1 ;
      RECT 120.19 37.98 120.39 38.18 ;
      RECT 120.19 42.06 120.39 42.26 ;
      RECT 120.19 46.14 120.39 46.34 ;
      RECT 120.19 50.22 120.39 50.42 ;
      RECT 120.19 54.3 120.39 54.5 ;
      RECT 120.19 58.38 120.39 58.58 ;
      RECT 119.27 19.69 119.47 19.89 ;
      RECT 119.27 20.91 119.47 21.11 ;
      RECT 118.35 18.94 118.55 19.14 ;
      RECT 118.35 23.02 118.55 23.22 ;
      RECT 118.35 27.1 118.55 27.3 ;
      RECT 118.35 31.18 118.55 31.38 ;
      RECT 118.35 35.26 118.55 35.46 ;
      RECT 118.35 39.34 118.55 39.54 ;
      RECT 118.35 43.42 118.55 43.62 ;
      RECT 118.35 47.5 118.55 47.7 ;
      RECT 118.35 51.58 118.55 51.78 ;
      RECT 118.35 55.66 118.55 55.86 ;
      RECT 118.35 59.74 118.55 59.94 ;
      RECT 117.43 17.58 117.63 17.78 ;
      RECT 117.43 21.66 117.63 21.86 ;
      RECT 117.43 25.74 117.63 25.94 ;
      RECT 117.43 29.82 117.63 30.02 ;
      RECT 117.43 33.9 117.63 34.1 ;
      RECT 117.43 37.98 117.63 38.18 ;
      RECT 117.43 42.06 117.63 42.26 ;
      RECT 117.43 46.14 117.63 46.34 ;
      RECT 117.43 50.22 117.63 50.42 ;
      RECT 117.43 54.3 117.63 54.5 ;
      RECT 117.43 58.38 117.63 58.58 ;
      RECT 116.51 20.91 116.71 21.11 ;
      RECT 115.59 18.94 115.79 19.14 ;
      RECT 115.59 23.02 115.79 23.22 ;
      RECT 115.59 27.1 115.79 27.3 ;
      RECT 115.59 31.18 115.79 31.38 ;
      RECT 115.59 35.26 115.79 35.46 ;
      RECT 115.59 39.34 115.79 39.54 ;
      RECT 115.59 43.42 115.79 43.62 ;
      RECT 115.59 47.5 115.79 47.7 ;
      RECT 115.59 51.58 115.79 51.78 ;
      RECT 115.59 55.66 115.79 55.86 ;
      RECT 115.59 59.74 115.79 59.94 ;
      RECT 114.67 17.58 114.87 17.78 ;
      RECT 114.67 21.66 114.87 21.86 ;
      RECT 114.67 25.74 114.87 25.94 ;
      RECT 114.67 29.82 114.87 30.02 ;
      RECT 114.67 33.9 114.87 34.1 ;
      RECT 114.67 37.98 114.87 38.18 ;
      RECT 114.67 42.06 114.87 42.26 ;
      RECT 114.67 46.14 114.87 46.34 ;
      RECT 114.67 50.22 114.87 50.42 ;
      RECT 114.67 54.3 114.87 54.5 ;
      RECT 114.67 58.38 114.87 58.58 ;
      RECT 112.83 18.94 113.03 19.14 ;
      RECT 112.83 23.02 113.03 23.22 ;
      RECT 112.83 27.1 113.03 27.3 ;
      RECT 112.83 31.18 113.03 31.38 ;
      RECT 112.83 35.26 113.03 35.46 ;
      RECT 112.83 39.34 113.03 39.54 ;
      RECT 112.83 43.42 113.03 43.62 ;
      RECT 112.83 47.5 113.03 47.7 ;
      RECT 112.83 51.58 113.03 51.78 ;
      RECT 112.83 55.66 113.03 55.86 ;
      RECT 112.83 59.74 113.03 59.94 ;
      RECT 111.91 17.58 112.11 17.78 ;
      RECT 111.91 21.66 112.11 21.86 ;
      RECT 111.91 25.74 112.11 25.94 ;
      RECT 111.91 29.82 112.11 30.02 ;
      RECT 111.91 33.9 112.11 34.1 ;
      RECT 111.91 37.98 112.11 38.18 ;
      RECT 111.91 42.06 112.11 42.26 ;
      RECT 111.91 46.14 112.11 46.34 ;
      RECT 111.91 50.22 112.11 50.42 ;
      RECT 111.91 54.3 112.11 54.5 ;
      RECT 111.91 58.38 112.11 58.58 ;
      RECT 110.99 19.69 111.19 19.89 ;
      RECT 110.07 18.94 110.27 19.14 ;
      RECT 110.07 23.02 110.27 23.22 ;
      RECT 110.07 27.1 110.27 27.3 ;
      RECT 110.07 31.18 110.27 31.38 ;
      RECT 110.07 35.26 110.27 35.46 ;
      RECT 110.07 39.34 110.27 39.54 ;
      RECT 110.07 43.42 110.27 43.62 ;
      RECT 110.07 47.5 110.27 47.7 ;
      RECT 110.07 51.58 110.27 51.78 ;
      RECT 110.07 55.66 110.27 55.86 ;
      RECT 110.07 59.74 110.27 59.94 ;
      RECT 109.15 17.58 109.35 17.78 ;
      RECT 109.15 21.66 109.35 21.86 ;
      RECT 109.15 25.74 109.35 25.94 ;
      RECT 109.15 29.82 109.35 30.02 ;
      RECT 109.15 33.9 109.35 34.1 ;
      RECT 109.15 37.98 109.35 38.18 ;
      RECT 109.15 42.06 109.35 42.26 ;
      RECT 109.15 46.14 109.35 46.34 ;
      RECT 109.15 50.22 109.35 50.42 ;
      RECT 109.15 54.3 109.35 54.5 ;
      RECT 109.15 58.38 109.35 58.58 ;
      RECT 108.23 20.91 108.43 21.11 ;
      RECT 107.31 18.94 107.51 19.14 ;
      RECT 107.31 23.02 107.51 23.22 ;
      RECT 107.31 27.1 107.51 27.3 ;
      RECT 107.31 31.18 107.51 31.38 ;
      RECT 107.31 35.26 107.51 35.46 ;
      RECT 107.31 39.34 107.51 39.54 ;
      RECT 107.31 43.42 107.51 43.62 ;
      RECT 107.31 47.5 107.51 47.7 ;
      RECT 107.31 51.58 107.51 51.78 ;
      RECT 107.31 55.66 107.51 55.86 ;
      RECT 107.31 59.74 107.51 59.94 ;
      RECT 106.39 17.58 106.59 17.78 ;
      RECT 106.39 21.66 106.59 21.86 ;
      RECT 106.39 25.74 106.59 25.94 ;
      RECT 106.39 29.82 106.59 30.02 ;
      RECT 106.39 33.9 106.59 34.1 ;
      RECT 106.39 37.98 106.59 38.18 ;
      RECT 106.39 42.06 106.59 42.26 ;
      RECT 106.39 46.14 106.59 46.34 ;
      RECT 106.39 50.22 106.59 50.42 ;
      RECT 106.39 54.3 106.59 54.5 ;
      RECT 106.39 58.38 106.59 58.58 ;
      RECT 105.47 20.91 105.67 21.11 ;
      RECT 105.47 23.96 105.67 24.16 ;
      RECT 104.55 18.94 104.75 19.14 ;
      RECT 104.55 23.02 104.75 23.22 ;
      RECT 104.55 27.1 104.75 27.3 ;
      RECT 104.55 31.18 104.75 31.38 ;
      RECT 104.55 35.26 104.75 35.46 ;
      RECT 104.55 39.34 104.75 39.54 ;
      RECT 104.55 43.42 104.75 43.62 ;
      RECT 104.55 47.5 104.75 47.7 ;
      RECT 104.55 51.58 104.75 51.78 ;
      RECT 104.55 55.66 104.75 55.86 ;
      RECT 104.55 59.74 104.75 59.94 ;
      RECT 103.63 17.58 103.83 17.78 ;
      RECT 103.63 21.66 103.83 21.86 ;
      RECT 103.63 25.74 103.83 25.94 ;
      RECT 103.63 29.82 103.83 30.02 ;
      RECT 103.63 33.9 103.83 34.1 ;
      RECT 103.63 37.98 103.83 38.18 ;
      RECT 103.63 42.06 103.83 42.26 ;
      RECT 103.63 46.14 103.83 46.34 ;
      RECT 103.63 50.22 103.83 50.42 ;
      RECT 103.63 54.3 103.83 54.5 ;
      RECT 103.63 58.38 103.83 58.58 ;
      RECT 102.71 19.69 102.91 19.89 ;
      RECT 101.79 18.94 101.99 19.14 ;
      RECT 101.79 23.02 101.99 23.22 ;
      RECT 101.79 27.1 101.99 27.3 ;
      RECT 101.79 31.18 101.99 31.38 ;
      RECT 101.79 35.26 101.99 35.46 ;
      RECT 101.79 39.34 101.99 39.54 ;
      RECT 101.79 43.42 101.99 43.62 ;
      RECT 101.79 47.5 101.99 47.7 ;
      RECT 101.79 51.58 101.99 51.78 ;
      RECT 101.79 55.66 101.99 55.86 ;
      RECT 101.79 59.74 101.99 59.94 ;
      RECT 100.87 17.58 101.07 17.78 ;
      RECT 100.87 21.66 101.07 21.86 ;
      RECT 100.87 25.74 101.07 25.94 ;
      RECT 100.87 29.82 101.07 30.02 ;
      RECT 100.87 33.9 101.07 34.1 ;
      RECT 100.87 37.98 101.07 38.18 ;
      RECT 100.87 42.06 101.07 42.26 ;
      RECT 100.87 46.14 101.07 46.34 ;
      RECT 100.87 50.22 101.07 50.42 ;
      RECT 100.87 54.3 101.07 54.5 ;
      RECT 100.87 58.38 101.07 58.58 ;
      RECT 99.95 20.91 100.15 21.11 ;
      RECT 99.95 32.5 100.15 32.7 ;
      RECT 99.03 18.94 99.23 19.14 ;
      RECT 99.03 23.02 99.23 23.22 ;
      RECT 99.03 27.1 99.23 27.3 ;
      RECT 99.03 31.18 99.23 31.38 ;
      RECT 99.03 35.26 99.23 35.46 ;
      RECT 99.03 39.34 99.23 39.54 ;
      RECT 99.03 43.42 99.23 43.62 ;
      RECT 99.03 47.5 99.23 47.7 ;
      RECT 99.03 51.58 99.23 51.78 ;
      RECT 99.03 55.66 99.23 55.86 ;
      RECT 99.03 59.74 99.23 59.94 ;
      RECT 98.11 17.58 98.31 17.78 ;
      RECT 98.11 21.66 98.31 21.86 ;
      RECT 98.11 25.74 98.31 25.94 ;
      RECT 98.11 29.82 98.31 30.02 ;
      RECT 98.11 33.9 98.31 34.1 ;
      RECT 98.11 37.98 98.31 38.18 ;
      RECT 98.11 42.06 98.31 42.26 ;
      RECT 98.11 46.14 98.31 46.34 ;
      RECT 98.11 50.22 98.31 50.42 ;
      RECT 98.11 54.3 98.31 54.5 ;
      RECT 98.11 58.38 98.31 58.58 ;
      RECT 97.19 20.91 97.39 21.11 ;
      RECT 97.19 24.57 97.39 24.77 ;
      RECT 96.27 18.94 96.47 19.14 ;
      RECT 96.27 23.02 96.47 23.22 ;
      RECT 96.27 27.1 96.47 27.3 ;
      RECT 96.27 31.18 96.47 31.38 ;
      RECT 96.27 35.26 96.47 35.46 ;
      RECT 96.27 39.34 96.47 39.54 ;
      RECT 96.27 43.42 96.47 43.62 ;
      RECT 96.27 47.5 96.47 47.7 ;
      RECT 96.27 51.58 96.47 51.78 ;
      RECT 96.27 55.66 96.47 55.86 ;
      RECT 96.27 59.74 96.47 59.94 ;
      RECT 95.35 17.58 95.55 17.78 ;
      RECT 95.35 21.66 95.55 21.86 ;
      RECT 95.35 25.74 95.55 25.94 ;
      RECT 95.35 29.82 95.55 30.02 ;
      RECT 95.35 33.9 95.55 34.1 ;
      RECT 95.35 37.98 95.55 38.18 ;
      RECT 95.35 42.06 95.55 42.26 ;
      RECT 95.35 46.14 95.55 46.34 ;
      RECT 95.35 50.22 95.55 50.42 ;
      RECT 95.35 54.3 95.55 54.5 ;
      RECT 95.35 58.38 95.55 58.58 ;
      RECT 94.43 19.69 94.63 19.89 ;
      RECT 94.43 36.16 94.63 36.36 ;
      RECT 93.51 18.94 93.71 19.14 ;
      RECT 93.51 23.02 93.71 23.22 ;
      RECT 93.51 27.1 93.71 27.3 ;
      RECT 93.51 31.18 93.71 31.38 ;
      RECT 93.51 35.26 93.71 35.46 ;
      RECT 93.51 39.34 93.71 39.54 ;
      RECT 93.51 43.42 93.71 43.62 ;
      RECT 93.51 47.5 93.71 47.7 ;
      RECT 93.51 51.58 93.71 51.78 ;
      RECT 93.51 55.66 93.71 55.86 ;
      RECT 93.51 59.74 93.71 59.94 ;
      RECT 92.59 17.58 92.79 17.78 ;
      RECT 92.59 21.66 92.79 21.86 ;
      RECT 92.59 25.74 92.79 25.94 ;
      RECT 92.59 29.82 92.79 30.02 ;
      RECT 92.59 33.9 92.79 34.1 ;
      RECT 92.59 37.98 92.79 38.18 ;
      RECT 92.59 42.06 92.79 42.26 ;
      RECT 92.59 46.14 92.79 46.34 ;
      RECT 92.59 50.22 92.79 50.42 ;
      RECT 92.59 54.3 92.79 54.5 ;
      RECT 92.59 58.38 92.79 58.58 ;
      RECT 91.67 16.64 91.87 16.84 ;
      RECT 91.67 24.57 91.87 24.77 ;
      RECT 91.67 36.16 91.87 36.36 ;
      RECT 90.75 18.94 90.95 19.14 ;
      RECT 90.75 23.02 90.95 23.22 ;
      RECT 90.75 27.1 90.95 27.3 ;
      RECT 90.75 31.18 90.95 31.38 ;
      RECT 90.75 35.26 90.95 35.46 ;
      RECT 90.75 39.34 90.95 39.54 ;
      RECT 90.75 43.42 90.95 43.62 ;
      RECT 90.75 47.5 90.95 47.7 ;
      RECT 90.75 51.58 90.95 51.78 ;
      RECT 90.75 55.66 90.95 55.86 ;
      RECT 90.75 59.74 90.95 59.94 ;
      RECT 89.83 17.58 90.03 17.78 ;
      RECT 89.83 21.66 90.03 21.86 ;
      RECT 89.83 25.74 90.03 25.94 ;
      RECT 89.83 29.82 90.03 30.02 ;
      RECT 89.83 33.9 90.03 34.1 ;
      RECT 89.83 37.98 90.03 38.18 ;
      RECT 89.83 42.06 90.03 42.26 ;
      RECT 89.83 46.14 90.03 46.34 ;
      RECT 89.83 50.22 90.03 50.42 ;
      RECT 89.83 54.3 90.03 54.5 ;
      RECT 89.83 58.38 90.03 58.58 ;
      RECT 88.91 20.91 89.11 21.11 ;
      RECT 87.99 18.94 88.19 19.14 ;
      RECT 87.99 23.02 88.19 23.22 ;
      RECT 87.99 27.1 88.19 27.3 ;
      RECT 87.99 31.18 88.19 31.38 ;
      RECT 87.99 35.26 88.19 35.46 ;
      RECT 87.99 39.34 88.19 39.54 ;
      RECT 87.99 43.42 88.19 43.62 ;
      RECT 87.99 47.5 88.19 47.7 ;
      RECT 87.99 51.58 88.19 51.78 ;
      RECT 87.99 55.66 88.19 55.86 ;
      RECT 87.99 59.74 88.19 59.94 ;
      RECT 87.07 17.58 87.27 17.78 ;
      RECT 87.07 21.66 87.27 21.86 ;
      RECT 87.07 25.74 87.27 25.94 ;
      RECT 87.07 29.82 87.27 30.02 ;
      RECT 87.07 33.9 87.27 34.1 ;
      RECT 87.07 37.98 87.27 38.18 ;
      RECT 87.07 42.06 87.27 42.26 ;
      RECT 87.07 46.14 87.27 46.34 ;
      RECT 87.07 50.22 87.27 50.42 ;
      RECT 87.07 54.3 87.27 54.5 ;
      RECT 87.07 58.38 87.27 58.58 ;
      RECT 86.15 24.57 86.35 24.77 ;
      RECT 86.15 32.5 86.35 32.7 ;
      RECT 85.23 18.94 85.43 19.14 ;
      RECT 85.23 23.02 85.43 23.22 ;
      RECT 85.23 27.1 85.43 27.3 ;
      RECT 85.23 31.18 85.43 31.38 ;
      RECT 85.23 35.26 85.43 35.46 ;
      RECT 85.23 39.34 85.43 39.54 ;
      RECT 85.23 43.42 85.43 43.62 ;
      RECT 85.23 47.5 85.43 47.7 ;
      RECT 85.23 51.58 85.43 51.78 ;
      RECT 85.23 55.66 85.43 55.86 ;
      RECT 85.23 59.74 85.43 59.94 ;
      RECT 84.31 17.58 84.51 17.78 ;
      RECT 84.31 21.66 84.51 21.86 ;
      RECT 84.31 25.74 84.51 25.94 ;
      RECT 84.31 29.82 84.51 30.02 ;
      RECT 84.31 33.9 84.51 34.1 ;
      RECT 84.31 37.98 84.51 38.18 ;
      RECT 84.31 42.06 84.51 42.26 ;
      RECT 84.31 46.14 84.51 46.34 ;
      RECT 84.31 50.22 84.51 50.42 ;
      RECT 84.31 54.3 84.51 54.5 ;
      RECT 84.31 58.38 84.51 58.58 ;
      RECT 82.47 18.94 82.67 19.14 ;
      RECT 82.47 23.02 82.67 23.22 ;
      RECT 82.47 27.1 82.67 27.3 ;
      RECT 82.47 31.18 82.67 31.38 ;
      RECT 82.47 35.26 82.67 35.46 ;
      RECT 82.47 39.34 82.67 39.54 ;
      RECT 82.47 43.42 82.67 43.62 ;
      RECT 82.47 47.5 82.67 47.7 ;
      RECT 82.47 51.58 82.67 51.78 ;
      RECT 82.47 55.66 82.67 55.86 ;
      RECT 82.47 59.74 82.67 59.94 ;
      RECT 81.55 17.58 81.75 17.78 ;
      RECT 81.55 21.66 81.75 21.86 ;
      RECT 81.55 25.74 81.75 25.94 ;
      RECT 81.55 29.82 81.75 30.02 ;
      RECT 81.55 33.9 81.75 34.1 ;
      RECT 81.55 37.98 81.75 38.18 ;
      RECT 81.55 42.06 81.75 42.26 ;
      RECT 81.55 46.14 81.75 46.34 ;
      RECT 81.55 50.22 81.75 50.42 ;
      RECT 81.55 54.3 81.75 54.5 ;
      RECT 81.55 58.38 81.75 58.58 ;
      RECT 79.71 18.94 79.91 19.14 ;
      RECT 79.71 23.02 79.91 23.22 ;
      RECT 79.71 27.1 79.91 27.3 ;
      RECT 79.71 31.18 79.91 31.38 ;
      RECT 79.71 35.26 79.91 35.46 ;
      RECT 79.71 39.34 79.91 39.54 ;
      RECT 79.71 43.42 79.91 43.62 ;
      RECT 79.71 47.5 79.91 47.7 ;
      RECT 79.71 51.58 79.91 51.78 ;
      RECT 79.71 55.66 79.91 55.86 ;
      RECT 79.71 59.74 79.91 59.94 ;
      RECT 78.79 17.58 78.99 17.78 ;
      RECT 78.79 21.66 78.99 21.86 ;
      RECT 78.79 25.74 78.99 25.94 ;
      RECT 78.79 29.82 78.99 30.02 ;
      RECT 78.79 33.9 78.99 34.1 ;
      RECT 78.79 37.98 78.99 38.18 ;
      RECT 78.79 42.06 78.99 42.26 ;
      RECT 78.79 46.14 78.99 46.34 ;
      RECT 78.79 50.22 78.99 50.42 ;
      RECT 78.79 54.3 78.99 54.5 ;
      RECT 78.79 58.38 78.99 58.58 ;
      RECT 77.87 15.42 78.07 15.62 ;
      RECT 77.87 24.57 78.07 24.77 ;
      RECT 76.95 18.94 77.15 19.14 ;
      RECT 76.95 23.02 77.15 23.22 ;
      RECT 76.95 27.1 77.15 27.3 ;
      RECT 76.95 31.18 77.15 31.38 ;
      RECT 76.95 35.26 77.15 35.46 ;
      RECT 76.95 39.34 77.15 39.54 ;
      RECT 76.95 43.42 77.15 43.62 ;
      RECT 76.95 47.5 77.15 47.7 ;
      RECT 76.95 51.58 77.15 51.78 ;
      RECT 76.95 55.66 77.15 55.86 ;
      RECT 76.95 59.74 77.15 59.94 ;
      RECT 76.03 17.58 76.23 17.78 ;
      RECT 76.03 21.66 76.23 21.86 ;
      RECT 76.03 25.74 76.23 25.94 ;
      RECT 76.03 29.82 76.23 30.02 ;
      RECT 76.03 33.9 76.23 34.1 ;
      RECT 76.03 37.98 76.23 38.18 ;
      RECT 76.03 42.06 76.23 42.26 ;
      RECT 76.03 46.14 76.23 46.34 ;
      RECT 76.03 50.22 76.23 50.42 ;
      RECT 76.03 54.3 76.23 54.5 ;
      RECT 76.03 58.38 76.23 58.58 ;
      RECT 75.495 24.57 75.695 24.77 ;
      RECT 75.11 16.64 75.31 16.84 ;
      RECT 74.19 18.94 74.39 19.14 ;
      RECT 74.19 23.02 74.39 23.22 ;
      RECT 74.19 27.1 74.39 27.3 ;
      RECT 74.19 31.18 74.39 31.38 ;
      RECT 74.19 35.26 74.39 35.46 ;
      RECT 74.19 39.34 74.39 39.54 ;
      RECT 74.19 43.42 74.39 43.62 ;
      RECT 74.19 47.5 74.39 47.7 ;
      RECT 74.19 51.58 74.39 51.78 ;
      RECT 74.19 55.66 74.39 55.86 ;
      RECT 74.19 59.74 74.39 59.94 ;
      RECT 73.27 17.58 73.47 17.78 ;
      RECT 73.27 21.66 73.47 21.86 ;
      RECT 73.27 25.74 73.47 25.94 ;
      RECT 73.27 29.82 73.47 30.02 ;
      RECT 73.27 33.9 73.47 34.1 ;
      RECT 73.27 37.98 73.47 38.18 ;
      RECT 73.27 42.06 73.47 42.26 ;
      RECT 73.27 46.14 73.47 46.34 ;
      RECT 73.27 50.22 73.47 50.42 ;
      RECT 73.27 54.3 73.47 54.5 ;
      RECT 73.27 58.38 73.47 58.58 ;
      RECT 72.35 14.2 72.55 14.4 ;
      RECT 72.35 16.64 72.55 16.84 ;
      RECT 72.35 19.69 72.55 19.89 ;
      RECT 71.43 18.94 71.63 19.14 ;
      RECT 71.43 23.02 71.63 23.22 ;
      RECT 71.43 27.1 71.63 27.3 ;
      RECT 71.43 31.18 71.63 31.38 ;
      RECT 71.43 35.26 71.63 35.46 ;
      RECT 71.43 39.34 71.63 39.54 ;
      RECT 71.43 43.42 71.63 43.62 ;
      RECT 71.43 47.5 71.63 47.7 ;
      RECT 71.43 51.58 71.63 51.78 ;
      RECT 71.43 55.66 71.63 55.86 ;
      RECT 71.43 59.74 71.63 59.94 ;
      RECT 70.51 17.58 70.71 17.78 ;
      RECT 70.51 21.66 70.71 21.86 ;
      RECT 70.51 25.74 70.71 25.94 ;
      RECT 70.51 29.82 70.71 30.02 ;
      RECT 70.51 33.9 70.71 34.1 ;
      RECT 70.51 37.98 70.71 38.18 ;
      RECT 70.51 42.06 70.71 42.26 ;
      RECT 70.51 46.14 70.71 46.34 ;
      RECT 70.51 50.22 70.71 50.42 ;
      RECT 70.51 54.3 70.71 54.5 ;
      RECT 70.51 58.38 70.71 58.58 ;
      RECT 68.67 18.94 68.87 19.14 ;
      RECT 68.67 23.02 68.87 23.22 ;
      RECT 68.67 27.1 68.87 27.3 ;
      RECT 68.67 31.18 68.87 31.38 ;
      RECT 68.67 35.26 68.87 35.46 ;
      RECT 68.67 39.34 68.87 39.54 ;
      RECT 68.67 43.42 68.87 43.62 ;
      RECT 68.67 47.5 68.87 47.7 ;
      RECT 68.67 51.58 68.87 51.78 ;
      RECT 68.67 55.66 68.87 55.86 ;
      RECT 68.67 59.74 68.87 59.94 ;
      RECT 67.75 17.58 67.95 17.78 ;
      RECT 67.75 21.66 67.95 21.86 ;
      RECT 67.75 25.74 67.95 25.94 ;
      RECT 67.75 29.82 67.95 30.02 ;
      RECT 67.75 33.9 67.95 34.1 ;
      RECT 67.75 37.98 67.95 38.18 ;
      RECT 67.75 42.06 67.95 42.26 ;
      RECT 67.75 46.14 67.95 46.34 ;
      RECT 67.75 50.22 67.95 50.42 ;
      RECT 67.75 54.3 67.95 54.5 ;
      RECT 67.75 58.38 67.95 58.58 ;
      RECT 66.83 13.59 67.03 13.79 ;
      RECT 65.91 18.94 66.11 19.14 ;
      RECT 65.91 23.02 66.11 23.22 ;
      RECT 65.91 27.1 66.11 27.3 ;
      RECT 65.91 31.18 66.11 31.38 ;
      RECT 65.91 35.26 66.11 35.46 ;
      RECT 65.91 39.34 66.11 39.54 ;
      RECT 65.91 43.42 66.11 43.62 ;
      RECT 65.91 47.5 66.11 47.7 ;
      RECT 65.91 51.58 66.11 51.78 ;
      RECT 65.91 55.66 66.11 55.86 ;
      RECT 65.91 59.74 66.11 59.94 ;
      RECT 64.99 17.58 65.19 17.78 ;
      RECT 64.99 21.66 65.19 21.86 ;
      RECT 64.99 25.74 65.19 25.94 ;
      RECT 64.99 29.82 65.19 30.02 ;
      RECT 64.99 33.9 65.19 34.1 ;
      RECT 64.99 37.98 65.19 38.18 ;
      RECT 64.99 42.06 65.19 42.26 ;
      RECT 64.99 46.14 65.19 46.34 ;
      RECT 64.99 50.22 65.19 50.42 ;
      RECT 64.99 54.3 65.19 54.5 ;
      RECT 64.99 58.38 65.19 58.58 ;
      RECT 63.15 18.94 63.35 19.14 ;
      RECT 63.15 23.02 63.35 23.22 ;
      RECT 63.15 27.1 63.35 27.3 ;
      RECT 63.15 31.18 63.35 31.38 ;
      RECT 63.15 35.26 63.35 35.46 ;
      RECT 63.15 39.34 63.35 39.54 ;
      RECT 63.15 43.42 63.35 43.62 ;
      RECT 63.15 47.5 63.35 47.7 ;
      RECT 63.15 51.58 63.35 51.78 ;
      RECT 63.15 55.66 63.35 55.86 ;
      RECT 63.15 59.74 63.35 59.94 ;
      RECT 62.23 17.58 62.43 17.78 ;
      RECT 62.23 21.66 62.43 21.86 ;
      RECT 62.23 25.74 62.43 25.94 ;
      RECT 62.23 29.82 62.43 30.02 ;
      RECT 62.23 33.9 62.43 34.1 ;
      RECT 62.23 37.98 62.43 38.18 ;
      RECT 62.23 42.06 62.43 42.26 ;
      RECT 62.23 46.14 62.43 46.34 ;
      RECT 62.23 50.22 62.43 50.42 ;
      RECT 62.23 54.3 62.43 54.5 ;
      RECT 62.23 58.38 62.43 58.58 ;
      RECT 61.31 15.42 61.51 15.62 ;
      RECT 61.31 16.64 61.51 16.84 ;
      RECT 60.39 18.94 60.59 19.14 ;
      RECT 60.39 23.02 60.59 23.22 ;
      RECT 60.39 27.1 60.59 27.3 ;
      RECT 60.39 31.18 60.59 31.38 ;
      RECT 60.39 35.26 60.59 35.46 ;
      RECT 60.39 39.34 60.59 39.54 ;
      RECT 60.39 43.42 60.59 43.62 ;
      RECT 60.39 47.5 60.59 47.7 ;
      RECT 60.39 51.58 60.59 51.78 ;
      RECT 60.39 55.66 60.59 55.86 ;
      RECT 60.39 59.74 60.59 59.94 ;
      RECT 59.47 17.58 59.67 17.78 ;
      RECT 59.47 21.66 59.67 21.86 ;
      RECT 59.47 25.74 59.67 25.94 ;
      RECT 59.47 29.82 59.67 30.02 ;
      RECT 59.47 33.9 59.67 34.1 ;
      RECT 59.47 37.98 59.67 38.18 ;
      RECT 59.47 42.06 59.67 42.26 ;
      RECT 59.47 46.14 59.67 46.34 ;
      RECT 59.47 50.22 59.67 50.42 ;
      RECT 59.47 54.3 59.67 54.5 ;
      RECT 59.47 58.38 59.67 58.58 ;
      RECT 58.55 19.69 58.75 19.89 ;
      RECT 57.63 18.94 57.83 19.14 ;
      RECT 57.63 23.02 57.83 23.22 ;
      RECT 57.63 27.1 57.83 27.3 ;
      RECT 57.63 31.18 57.83 31.38 ;
      RECT 57.63 35.26 57.83 35.46 ;
      RECT 57.63 39.34 57.83 39.54 ;
      RECT 57.63 43.42 57.83 43.62 ;
      RECT 57.63 47.5 57.83 47.7 ;
      RECT 57.63 51.58 57.83 51.78 ;
      RECT 57.63 55.66 57.83 55.86 ;
      RECT 57.63 59.74 57.83 59.94 ;
      RECT 56.71 17.58 56.91 17.78 ;
      RECT 56.71 21.66 56.91 21.86 ;
      RECT 56.71 25.74 56.91 25.94 ;
      RECT 56.71 29.82 56.91 30.02 ;
      RECT 56.71 33.9 56.91 34.1 ;
      RECT 56.71 37.98 56.91 38.18 ;
      RECT 56.71 42.06 56.91 42.26 ;
      RECT 56.71 46.14 56.91 46.34 ;
      RECT 56.71 50.22 56.91 50.42 ;
      RECT 56.71 54.3 56.91 54.5 ;
      RECT 56.71 58.38 56.91 58.58 ;
      RECT 55.79 24.57 55.99 24.77 ;
      RECT 54.87 18.94 55.07 19.14 ;
      RECT 54.87 23.02 55.07 23.22 ;
      RECT 54.87 27.1 55.07 27.3 ;
      RECT 54.87 31.18 55.07 31.38 ;
      RECT 54.87 35.26 55.07 35.46 ;
      RECT 54.87 39.34 55.07 39.54 ;
      RECT 54.87 43.42 55.07 43.62 ;
      RECT 54.87 47.5 55.07 47.7 ;
      RECT 54.87 51.58 55.07 51.78 ;
      RECT 54.87 55.66 55.07 55.86 ;
      RECT 54.87 59.74 55.07 59.94 ;
      RECT 53.95 17.58 54.15 17.78 ;
      RECT 53.95 21.66 54.15 21.86 ;
      RECT 53.95 25.74 54.15 25.94 ;
      RECT 53.95 29.82 54.15 30.02 ;
      RECT 53.95 33.9 54.15 34.1 ;
      RECT 53.95 37.98 54.15 38.18 ;
      RECT 53.95 42.06 54.15 42.26 ;
      RECT 53.95 46.14 54.15 46.34 ;
      RECT 53.95 50.22 54.15 50.42 ;
      RECT 53.95 54.3 54.15 54.5 ;
      RECT 53.95 58.38 54.15 58.58 ;
      RECT 53.03 13.59 53.23 13.79 ;
      RECT 53.03 24.57 53.23 24.77 ;
      RECT 52.11 18.94 52.31 19.14 ;
      RECT 52.11 23.02 52.31 23.22 ;
      RECT 52.11 27.1 52.31 27.3 ;
      RECT 52.11 31.18 52.31 31.38 ;
      RECT 52.11 35.26 52.31 35.46 ;
      RECT 52.11 39.34 52.31 39.54 ;
      RECT 52.11 43.42 52.31 43.62 ;
      RECT 52.11 47.5 52.31 47.7 ;
      RECT 52.11 51.58 52.31 51.78 ;
      RECT 52.11 55.66 52.31 55.86 ;
      RECT 52.11 59.74 52.31 59.94 ;
      RECT 51.19 17.58 51.39 17.78 ;
      RECT 51.19 21.66 51.39 21.86 ;
      RECT 51.19 25.74 51.39 25.94 ;
      RECT 51.19 29.82 51.39 30.02 ;
      RECT 51.19 33.9 51.39 34.1 ;
      RECT 51.19 37.98 51.39 38.18 ;
      RECT 51.19 42.06 51.39 42.26 ;
      RECT 51.19 46.14 51.39 46.34 ;
      RECT 51.19 50.22 51.39 50.42 ;
      RECT 51.19 54.3 51.39 54.5 ;
      RECT 51.19 58.38 51.39 58.58 ;
      RECT 50.27 14.2 50.47 14.4 ;
      RECT 49.35 18.94 49.55 19.14 ;
      RECT 49.35 23.02 49.55 23.22 ;
      RECT 49.35 27.1 49.55 27.3 ;
      RECT 49.35 31.18 49.55 31.38 ;
      RECT 49.35 35.26 49.55 35.46 ;
      RECT 49.35 39.34 49.55 39.54 ;
      RECT 49.35 43.42 49.55 43.62 ;
      RECT 49.35 47.5 49.55 47.7 ;
      RECT 49.35 51.58 49.55 51.78 ;
      RECT 49.35 55.66 49.55 55.86 ;
      RECT 49.35 59.74 49.55 59.94 ;
      RECT 48.43 17.58 48.63 17.78 ;
      RECT 48.43 21.66 48.63 21.86 ;
      RECT 48.43 25.74 48.63 25.94 ;
      RECT 48.43 29.82 48.63 30.02 ;
      RECT 48.43 33.9 48.63 34.1 ;
      RECT 48.43 37.98 48.63 38.18 ;
      RECT 48.43 42.06 48.63 42.26 ;
      RECT 48.43 46.14 48.63 46.34 ;
      RECT 48.43 50.22 48.63 50.42 ;
      RECT 48.43 54.3 48.63 54.5 ;
      RECT 48.43 58.38 48.63 58.58 ;
      RECT 47.51 19.69 47.71 19.89 ;
      RECT 46.59 18.94 46.79 19.14 ;
      RECT 46.59 23.02 46.79 23.22 ;
      RECT 46.59 27.1 46.79 27.3 ;
      RECT 46.59 31.18 46.79 31.38 ;
      RECT 46.59 35.26 46.79 35.46 ;
      RECT 46.59 39.34 46.79 39.54 ;
      RECT 46.59 43.42 46.79 43.62 ;
      RECT 46.59 47.5 46.79 47.7 ;
      RECT 46.59 51.58 46.79 51.78 ;
      RECT 46.59 55.66 46.79 55.86 ;
      RECT 46.59 59.74 46.79 59.94 ;
      RECT 45.67 17.58 45.87 17.78 ;
      RECT 45.67 21.66 45.87 21.86 ;
      RECT 45.67 25.74 45.87 25.94 ;
      RECT 45.67 29.82 45.87 30.02 ;
      RECT 45.67 33.9 45.87 34.1 ;
      RECT 45.67 37.98 45.87 38.18 ;
      RECT 45.67 42.06 45.87 42.26 ;
      RECT 45.67 46.14 45.87 46.34 ;
      RECT 45.67 50.22 45.87 50.42 ;
      RECT 45.67 54.3 45.87 54.5 ;
      RECT 45.67 58.38 45.87 58.58 ;
      RECT 44.75 14.2 44.95 14.4 ;
      RECT 44.75 24.57 44.95 24.77 ;
      RECT 43.83 18.94 44.03 19.14 ;
      RECT 43.83 23.02 44.03 23.22 ;
      RECT 43.83 27.1 44.03 27.3 ;
      RECT 43.83 31.18 44.03 31.38 ;
      RECT 43.83 35.26 44.03 35.46 ;
      RECT 43.83 39.34 44.03 39.54 ;
      RECT 43.83 43.42 44.03 43.62 ;
      RECT 43.83 47.5 44.03 47.7 ;
      RECT 43.83 51.58 44.03 51.78 ;
      RECT 43.83 55.66 44.03 55.86 ;
      RECT 43.83 59.74 44.03 59.94 ;
      RECT 42.91 17.58 43.11 17.78 ;
      RECT 42.91 21.66 43.11 21.86 ;
      RECT 42.91 25.74 43.11 25.94 ;
      RECT 42.91 29.82 43.11 30.02 ;
      RECT 42.91 33.9 43.11 34.1 ;
      RECT 42.91 37.98 43.11 38.18 ;
      RECT 42.91 42.06 43.11 42.26 ;
      RECT 42.91 46.14 43.11 46.34 ;
      RECT 42.91 50.22 43.11 50.42 ;
      RECT 42.91 54.3 43.11 54.5 ;
      RECT 42.91 58.38 43.11 58.58 ;
      RECT 41.99 23.96 42.19 24.16 ;
      RECT 41.07 18.94 41.27 19.14 ;
      RECT 41.07 23.02 41.27 23.22 ;
      RECT 41.07 27.1 41.27 27.3 ;
      RECT 41.07 31.18 41.27 31.38 ;
      RECT 41.07 35.26 41.27 35.46 ;
      RECT 41.07 39.34 41.27 39.54 ;
      RECT 41.07 43.42 41.27 43.62 ;
      RECT 41.07 47.5 41.27 47.7 ;
      RECT 41.07 51.58 41.27 51.78 ;
      RECT 41.07 55.66 41.27 55.86 ;
      RECT 41.07 59.74 41.27 59.94 ;
      RECT 40.15 17.58 40.35 17.78 ;
      RECT 40.15 21.66 40.35 21.86 ;
      RECT 40.15 25.74 40.35 25.94 ;
      RECT 40.15 29.82 40.35 30.02 ;
      RECT 40.15 33.9 40.35 34.1 ;
      RECT 40.15 37.98 40.35 38.18 ;
      RECT 40.15 42.06 40.35 42.26 ;
      RECT 40.15 46.14 40.35 46.34 ;
      RECT 40.15 50.22 40.35 50.42 ;
      RECT 40.15 54.3 40.35 54.5 ;
      RECT 40.15 58.38 40.35 58.58 ;
      RECT 38.31 18.94 38.51 19.14 ;
      RECT 38.31 23.02 38.51 23.22 ;
      RECT 38.31 27.1 38.51 27.3 ;
      RECT 38.31 31.18 38.51 31.38 ;
      RECT 38.31 35.26 38.51 35.46 ;
      RECT 38.31 39.34 38.51 39.54 ;
      RECT 38.31 43.42 38.51 43.62 ;
      RECT 38.31 47.5 38.51 47.7 ;
      RECT 38.31 51.58 38.51 51.78 ;
      RECT 38.31 55.66 38.51 55.86 ;
      RECT 38.31 59.74 38.51 59.94 ;
      RECT 37.39 17.58 37.59 17.78 ;
      RECT 37.39 21.66 37.59 21.86 ;
      RECT 37.39 25.74 37.59 25.94 ;
      RECT 37.39 29.82 37.59 30.02 ;
      RECT 37.39 33.9 37.59 34.1 ;
      RECT 37.39 37.98 37.59 38.18 ;
      RECT 37.39 42.06 37.59 42.26 ;
      RECT 37.39 46.14 37.59 46.34 ;
      RECT 37.39 50.22 37.59 50.42 ;
      RECT 37.39 54.3 37.59 54.5 ;
      RECT 37.39 58.38 37.59 58.58 ;
      RECT 36.47 23.96 36.67 24.16 ;
      RECT 35.55 18.94 35.75 19.14 ;
      RECT 35.55 23.02 35.75 23.22 ;
      RECT 35.55 27.1 35.75 27.3 ;
      RECT 35.55 31.18 35.75 31.38 ;
      RECT 35.55 35.26 35.75 35.46 ;
      RECT 35.55 39.34 35.75 39.54 ;
      RECT 35.55 43.42 35.75 43.62 ;
      RECT 35.55 47.5 35.75 47.7 ;
      RECT 35.55 51.58 35.75 51.78 ;
      RECT 35.55 55.66 35.75 55.86 ;
      RECT 35.55 59.74 35.75 59.94 ;
      RECT 34.63 17.58 34.83 17.78 ;
      RECT 34.63 21.66 34.83 21.86 ;
      RECT 34.63 25.74 34.83 25.94 ;
      RECT 34.63 29.82 34.83 30.02 ;
      RECT 34.63 33.9 34.83 34.1 ;
      RECT 34.63 37.98 34.83 38.18 ;
      RECT 34.63 42.06 34.83 42.26 ;
      RECT 34.63 46.14 34.83 46.34 ;
      RECT 34.63 50.22 34.83 50.42 ;
      RECT 34.63 54.3 34.83 54.5 ;
      RECT 34.63 58.38 34.83 58.58 ;
      RECT 33.71 19.69 33.91 19.89 ;
      RECT 32.79 18.94 32.99 19.14 ;
      RECT 32.79 23.02 32.99 23.22 ;
      RECT 32.79 27.1 32.99 27.3 ;
      RECT 32.79 31.18 32.99 31.38 ;
      RECT 32.79 35.26 32.99 35.46 ;
      RECT 32.79 39.34 32.99 39.54 ;
      RECT 32.79 43.42 32.99 43.62 ;
      RECT 32.79 47.5 32.99 47.7 ;
      RECT 32.79 51.58 32.99 51.78 ;
      RECT 32.79 55.66 32.99 55.86 ;
      RECT 32.79 59.74 32.99 59.94 ;
      RECT 31.87 17.58 32.07 17.78 ;
      RECT 31.87 21.66 32.07 21.86 ;
      RECT 31.87 25.74 32.07 25.94 ;
      RECT 31.87 29.82 32.07 30.02 ;
      RECT 31.87 33.9 32.07 34.1 ;
      RECT 31.87 37.98 32.07 38.18 ;
      RECT 31.87 42.06 32.07 42.26 ;
      RECT 31.87 46.14 32.07 46.34 ;
      RECT 31.87 50.22 32.07 50.42 ;
      RECT 31.87 54.3 32.07 54.5 ;
      RECT 31.87 58.38 32.07 58.58 ;
      RECT 30.03 18.94 30.23 19.14 ;
      RECT 30.03 23.02 30.23 23.22 ;
      RECT 30.03 27.1 30.23 27.3 ;
      RECT 30.03 31.18 30.23 31.38 ;
      RECT 30.03 35.26 30.23 35.46 ;
      RECT 30.03 39.34 30.23 39.54 ;
      RECT 30.03 43.42 30.23 43.62 ;
      RECT 30.03 47.5 30.23 47.7 ;
      RECT 30.03 51.58 30.23 51.78 ;
      RECT 30.03 55.66 30.23 55.86 ;
      RECT 30.03 59.74 30.23 59.94 ;
      RECT 29.11 17.58 29.31 17.78 ;
      RECT 29.11 21.66 29.31 21.86 ;
      RECT 29.11 25.74 29.31 25.94 ;
      RECT 29.11 29.82 29.31 30.02 ;
      RECT 29.11 33.9 29.31 34.1 ;
      RECT 29.11 37.98 29.31 38.18 ;
      RECT 29.11 42.06 29.31 42.26 ;
      RECT 29.11 46.14 29.31 46.34 ;
      RECT 29.11 50.22 29.31 50.42 ;
      RECT 29.11 54.3 29.31 54.5 ;
      RECT 29.11 58.38 29.31 58.58 ;
      RECT 27.27 18.94 27.47 19.14 ;
      RECT 27.27 23.02 27.47 23.22 ;
      RECT 27.27 27.1 27.47 27.3 ;
      RECT 27.27 31.18 27.47 31.38 ;
      RECT 27.27 35.26 27.47 35.46 ;
      RECT 27.27 39.34 27.47 39.54 ;
      RECT 27.27 43.42 27.47 43.62 ;
      RECT 27.27 47.5 27.47 47.7 ;
      RECT 27.27 51.58 27.47 51.78 ;
      RECT 27.27 55.66 27.47 55.86 ;
      RECT 27.27 59.74 27.47 59.94 ;
      RECT 26.35 17.58 26.55 17.78 ;
      RECT 26.35 21.66 26.55 21.86 ;
      RECT 26.35 25.74 26.55 25.94 ;
      RECT 26.35 29.82 26.55 30.02 ;
      RECT 26.35 33.9 26.55 34.1 ;
      RECT 26.35 37.98 26.55 38.18 ;
      RECT 26.35 42.06 26.55 42.26 ;
      RECT 26.35 46.14 26.55 46.34 ;
      RECT 26.35 50.22 26.55 50.42 ;
      RECT 26.35 54.3 26.55 54.5 ;
      RECT 26.35 58.38 26.55 58.58 ;
      RECT 24.51 18.94 24.71 19.14 ;
      RECT 24.51 23.02 24.71 23.22 ;
      RECT 24.51 27.1 24.71 27.3 ;
      RECT 24.51 31.18 24.71 31.38 ;
      RECT 24.51 35.26 24.71 35.46 ;
      RECT 24.51 39.34 24.71 39.54 ;
      RECT 24.51 43.42 24.71 43.62 ;
      RECT 24.51 47.5 24.71 47.7 ;
      RECT 24.51 51.58 24.71 51.78 ;
      RECT 24.51 55.66 24.71 55.86 ;
      RECT 24.51 59.74 24.71 59.94 ;
      RECT 23.59 17.58 23.79 17.78 ;
      RECT 23.59 21.66 23.79 21.86 ;
      RECT 23.59 25.74 23.79 25.94 ;
      RECT 23.59 29.82 23.79 30.02 ;
      RECT 23.59 33.9 23.79 34.1 ;
      RECT 23.59 37.98 23.79 38.18 ;
      RECT 23.59 42.06 23.79 42.26 ;
      RECT 23.59 46.14 23.79 46.34 ;
      RECT 23.59 50.22 23.79 50.42 ;
      RECT 23.59 54.3 23.79 54.5 ;
      RECT 23.59 58.38 23.79 58.58 ;
      RECT 21.75 18.94 21.95 19.14 ;
      RECT 21.75 23.02 21.95 23.22 ;
      RECT 21.75 27.1 21.95 27.3 ;
      RECT 21.75 31.18 21.95 31.38 ;
      RECT 21.75 35.26 21.95 35.46 ;
      RECT 21.75 39.34 21.95 39.54 ;
      RECT 21.75 43.42 21.95 43.62 ;
      RECT 21.75 47.5 21.95 47.7 ;
      RECT 21.75 51.58 21.95 51.78 ;
      RECT 21.75 55.66 21.95 55.86 ;
      RECT 21.75 59.74 21.95 59.94 ;
      RECT 20.83 17.58 21.03 17.78 ;
      RECT 20.83 21.66 21.03 21.86 ;
      RECT 20.83 25.74 21.03 25.94 ;
      RECT 20.83 29.82 21.03 30.02 ;
      RECT 20.83 33.9 21.03 34.1 ;
      RECT 20.83 37.98 21.03 38.18 ;
      RECT 20.83 42.06 21.03 42.26 ;
      RECT 20.83 46.14 21.03 46.34 ;
      RECT 20.83 50.22 21.03 50.42 ;
      RECT 20.83 54.3 21.03 54.5 ;
      RECT 20.83 58.38 21.03 58.58 ;
      RECT 18.99 18.94 19.19 19.14 ;
      RECT 18.99 23.02 19.19 23.22 ;
      RECT 18.99 27.1 19.19 27.3 ;
      RECT 18.99 31.18 19.19 31.38 ;
      RECT 18.99 35.26 19.19 35.46 ;
      RECT 18.99 39.34 19.19 39.54 ;
      RECT 18.99 43.42 19.19 43.62 ;
      RECT 18.99 47.5 19.19 47.7 ;
      RECT 18.99 51.58 19.19 51.78 ;
      RECT 18.99 55.66 19.19 55.86 ;
      RECT 18.99 59.74 19.19 59.94 ;
      RECT 18.07 17.58 18.27 17.78 ;
      RECT 18.07 21.66 18.27 21.86 ;
      RECT 18.07 25.74 18.27 25.94 ;
      RECT 18.07 29.82 18.27 30.02 ;
      RECT 18.07 33.9 18.27 34.1 ;
      RECT 18.07 37.98 18.27 38.18 ;
      RECT 18.07 42.06 18.27 42.26 ;
      RECT 18.07 46.14 18.27 46.34 ;
      RECT 18.07 50.22 18.27 50.42 ;
      RECT 18.07 54.3 18.27 54.5 ;
      RECT 18.07 58.38 18.27 58.58 ;
      RECT 16.23 18.94 16.43 19.14 ;
      RECT 16.23 23.02 16.43 23.22 ;
      RECT 16.23 27.1 16.43 27.3 ;
      RECT 16.23 31.18 16.43 31.38 ;
      RECT 16.23 35.26 16.43 35.46 ;
      RECT 16.23 39.34 16.43 39.54 ;
      RECT 16.23 43.42 16.43 43.62 ;
      RECT 16.23 47.5 16.43 47.7 ;
      RECT 16.23 51.58 16.43 51.78 ;
      RECT 16.23 55.66 16.43 55.86 ;
      RECT 16.23 59.74 16.43 59.94 ;
      RECT 15.31 17.58 15.51 17.78 ;
      RECT 15.31 21.66 15.51 21.86 ;
      RECT 15.31 25.74 15.51 25.94 ;
      RECT 15.31 29.82 15.51 30.02 ;
      RECT 15.31 33.9 15.51 34.1 ;
      RECT 15.31 37.98 15.51 38.18 ;
      RECT 15.31 42.06 15.51 42.26 ;
      RECT 15.31 46.14 15.51 46.34 ;
      RECT 15.31 50.22 15.51 50.42 ;
      RECT 15.31 54.3 15.51 54.5 ;
      RECT 15.31 58.38 15.51 58.58 ;
    LAYER met3 ;
      RECT 177.165 15.355 177.495 15.685 ;
      RECT 157.845 15.355 158.175 15.685 ;
      RECT 157.845 15.37 177.495 15.67 ;
      RECT 168.885 9.255 169.215 9.585 ;
      RECT 150.025 9.255 150.355 9.585 ;
      RECT 150.025 9.27 169.215 9.57 ;
      RECT 160.605 16.575 160.935 16.905 ;
      RECT 138.525 16.575 138.855 16.905 ;
      RECT 124.725 16.575 125.055 16.905 ;
      RECT 124.725 16.59 160.935 16.89 ;
      RECT 146.09 20.85 146.47 21.17 ;
      RECT 146.09 20.86 149.42 21.16 ;
      RECT 149.12 19.64 149.42 21.16 ;
      RECT 160.605 19.625 160.935 19.955 ;
      RECT 149.12 19.64 160.935 19.94 ;
      RECT 149.565 24.505 149.895 24.835 ;
      RECT 141.285 24.505 141.615 24.835 ;
      RECT 146.09 24.51 146.47 24.83 ;
      RECT 139.88 24.51 140.26 24.83 ;
      RECT 139.88 24.52 149.895 24.82 ;
      RECT 141.285 20.845 141.615 21.175 ;
      RECT 133.005 20.845 133.335 21.175 ;
      RECT 133.005 20.86 141.615 21.16 ;
      RECT 133.005 28.775 133.335 29.105 ;
      RECT 139.88 28.78 140.26 29.1 ;
      RECT 133.005 28.79 140.26 29.09 ;
      RECT 135.765 23.895 136.095 24.225 ;
      RECT 135.05 23.9 135.43 24.22 ;
      RECT 135.05 23.91 136.095 24.21 ;
      RECT 124.725 15.355 125.055 15.685 ;
      RECT 135.05 15.36 135.43 15.68 ;
      RECT 133.48 15.37 135.43 15.67 ;
      RECT 124.725 15.37 126.42 15.67 ;
      RECT 126.12 14.76 126.42 15.67 ;
      RECT 133.48 14.76 133.78 15.67 ;
      RECT 126.12 14.76 133.78 15.06 ;
      RECT 133.005 19.625 133.335 19.955 ;
      RECT 119.205 19.625 119.535 19.955 ;
      RECT 110.925 19.625 111.255 19.955 ;
      RECT 102.645 19.625 102.975 19.955 ;
      RECT 94.365 19.625 94.695 19.955 ;
      RECT 94.365 19.64 133.335 19.94 ;
      RECT 127.485 20.845 127.815 21.175 ;
      RECT 119.205 20.845 119.535 21.175 ;
      RECT 119.205 20.86 127.815 21.16 ;
      RECT 127.485 28.165 127.815 28.495 ;
      RECT 118.49 28.17 118.87 28.49 ;
      RECT 118.49 28.18 127.815 28.48 ;
      RECT 121.965 14.135 122.295 14.465 ;
      RECT 72.285 14.135 72.615 14.465 ;
      RECT 72.285 14.15 122.295 14.45 ;
      RECT 106.8 24.215 120.9 24.515 ;
      RECT 120.6 23.91 120.9 24.515 ;
      RECT 121.965 23.895 122.295 24.225 ;
      RECT 105.405 23.895 105.735 24.225 ;
      RECT 106.8 23.91 107.1 24.515 ;
      RECT 120.6 23.91 122.295 24.21 ;
      RECT 105.405 23.91 107.1 24.21 ;
      RECT 116.445 20.845 116.775 21.175 ;
      RECT 108.165 20.845 108.495 21.175 ;
      RECT 118.49 20.85 118.87 21.17 ;
      RECT 108.165 20.86 118.87 21.16 ;
      RECT 105.405 20.845 105.735 21.175 ;
      RECT 99.885 20.845 100.215 21.175 ;
      RECT 99.885 20.86 105.735 21.16 ;
      RECT 99.885 32.435 100.215 32.765 ;
      RECT 86.085 32.435 86.415 32.765 ;
      RECT 86.085 32.45 100.215 32.75 ;
      RECT 97.125 20.845 97.455 21.175 ;
      RECT 88.845 20.845 89.175 21.175 ;
      RECT 95.72 20.85 96.1 21.17 ;
      RECT 88.845 20.86 97.455 21.16 ;
      RECT 97.125 24.505 97.455 24.835 ;
      RECT 91.605 24.505 91.935 24.835 ;
      RECT 91.605 24.52 97.455 24.82 ;
      RECT 91.605 16.575 91.935 16.905 ;
      RECT 95.72 16.58 96.1 16.9 ;
      RECT 91.605 16.59 96.1 16.89 ;
      RECT 94.365 36.095 94.695 36.425 ;
      RECT 91.605 36.095 91.935 36.425 ;
      RECT 91.605 36.11 94.695 36.41 ;
      RECT 86.085 24.505 86.415 24.835 ;
      RECT 77.805 24.505 78.135 24.835 ;
      RECT 75.43 24.505 75.76 24.835 ;
      RECT 55.725 24.505 56.055 24.835 ;
      RECT 55.725 24.52 86.415 24.82 ;
      RECT 77.805 15.355 78.135 15.685 ;
      RECT 61.245 15.355 61.575 15.685 ;
      RECT 61.245 15.37 78.135 15.67 ;
      RECT 75.045 16.575 75.375 16.905 ;
      RECT 74.33 16.58 74.71 16.9 ;
      RECT 74.33 16.59 75.375 16.89 ;
      RECT 72.285 19.625 72.615 19.955 ;
      RECT 74.33 19.63 74.71 19.95 ;
      RECT 72.285 19.64 74.71 19.94 ;
      RECT 72.285 16.575 72.615 16.905 ;
      RECT 61.245 16.575 61.575 16.905 ;
      RECT 61.245 16.59 72.615 16.89 ;
      RECT 66.765 13.525 67.095 13.855 ;
      RECT 52.965 13.525 53.295 13.855 ;
      RECT 52.965 13.54 67.095 13.84 ;
      RECT 58.485 19.625 58.815 19.955 ;
      RECT 47.445 19.625 47.775 19.955 ;
      RECT 33.645 19.625 33.975 19.955 ;
      RECT 33.645 19.64 58.815 19.94 ;
      RECT 52.965 24.505 53.295 24.835 ;
      RECT 44.685 24.505 45.015 24.835 ;
      RECT 44.685 24.52 53.295 24.82 ;
      RECT 50.205 14.135 50.535 14.465 ;
      RECT 44.685 14.135 45.015 14.465 ;
      RECT 44.685 14.15 50.535 14.45 ;
      RECT 41.925 23.895 42.255 24.225 ;
      RECT 36.405 23.895 36.735 24.225 ;
      RECT 36.405 23.91 42.255 24.21 ;
      RECT 10.12 17.45 189.98 17.91 ;
      RECT 10.12 18.81 189.98 19.27 ;
      RECT 10.12 21.53 189.98 21.99 ;
      RECT 10.12 22.89 189.98 23.35 ;
      RECT 10.12 25.61 189.98 26.07 ;
      RECT 10.12 26.97 189.98 27.43 ;
      RECT 10.12 29.69 189.98 30.15 ;
      RECT 10.12 31.05 189.98 31.51 ;
      RECT 10.12 33.77 189.98 34.23 ;
      RECT 10.12 35.13 189.98 35.59 ;
      RECT 10.12 37.85 189.98 38.31 ;
      RECT 10.12 39.21 189.98 39.67 ;
      RECT 10.12 41.93 189.98 42.39 ;
      RECT 10.12 43.29 189.98 43.75 ;
      RECT 10.12 46.01 189.98 46.47 ;
      RECT 10.12 47.37 189.98 47.83 ;
      RECT 10.12 50.09 189.98 50.55 ;
      RECT 10.12 51.45 189.98 51.91 ;
      RECT 10.12 54.17 189.98 54.63 ;
      RECT 10.12 55.53 189.98 55.99 ;
      RECT 10.12 58.25 189.98 58.71 ;
      RECT 10.12 59.61 189.98 60.07 ;
    LAYER via3 ;
      RECT 188.24 18.94 188.44 19.14 ;
      RECT 188.24 23.02 188.44 23.22 ;
      RECT 188.24 27.1 188.44 27.3 ;
      RECT 188.24 31.18 188.44 31.38 ;
      RECT 188.24 35.26 188.44 35.46 ;
      RECT 188.24 39.34 188.44 39.54 ;
      RECT 188.24 43.42 188.44 43.62 ;
      RECT 188.24 47.5 188.44 47.7 ;
      RECT 188.24 51.58 188.44 51.78 ;
      RECT 188.24 55.66 188.44 55.86 ;
      RECT 188.24 59.74 188.44 59.94 ;
      RECT 187.84 18.94 188.04 19.14 ;
      RECT 187.84 23.02 188.04 23.22 ;
      RECT 187.84 27.1 188.04 27.3 ;
      RECT 187.84 31.18 188.04 31.38 ;
      RECT 187.84 35.26 188.04 35.46 ;
      RECT 187.84 39.34 188.04 39.54 ;
      RECT 187.84 43.42 188.04 43.62 ;
      RECT 187.84 47.5 188.04 47.7 ;
      RECT 187.84 51.58 188.04 51.78 ;
      RECT 187.84 55.66 188.04 55.86 ;
      RECT 187.84 59.74 188.04 59.94 ;
      RECT 186.4 17.58 186.6 17.78 ;
      RECT 186.4 21.66 186.6 21.86 ;
      RECT 186.4 25.74 186.6 25.94 ;
      RECT 186.4 29.82 186.6 30.02 ;
      RECT 186.4 33.9 186.6 34.1 ;
      RECT 186.4 37.98 186.6 38.18 ;
      RECT 186.4 42.06 186.6 42.26 ;
      RECT 186.4 46.14 186.6 46.34 ;
      RECT 186.4 50.22 186.6 50.42 ;
      RECT 186.4 54.3 186.6 54.5 ;
      RECT 186.4 58.38 186.6 58.58 ;
      RECT 186 17.58 186.2 17.78 ;
      RECT 186 21.66 186.2 21.86 ;
      RECT 186 25.74 186.2 25.94 ;
      RECT 186 29.82 186.2 30.02 ;
      RECT 186 33.9 186.2 34.1 ;
      RECT 186 37.98 186.2 38.18 ;
      RECT 186 42.06 186.2 42.26 ;
      RECT 186 46.14 186.2 46.34 ;
      RECT 186 50.22 186.2 50.42 ;
      RECT 186 54.3 186.2 54.5 ;
      RECT 186 58.38 186.2 58.58 ;
      RECT 182.72 18.94 182.92 19.14 ;
      RECT 182.72 23.02 182.92 23.22 ;
      RECT 182.72 27.1 182.92 27.3 ;
      RECT 182.72 31.18 182.92 31.38 ;
      RECT 182.72 35.26 182.92 35.46 ;
      RECT 182.72 39.34 182.92 39.54 ;
      RECT 182.72 43.42 182.92 43.62 ;
      RECT 182.72 47.5 182.92 47.7 ;
      RECT 182.72 51.58 182.92 51.78 ;
      RECT 182.72 55.66 182.92 55.86 ;
      RECT 182.72 59.74 182.92 59.94 ;
      RECT 182.32 18.94 182.52 19.14 ;
      RECT 182.32 23.02 182.52 23.22 ;
      RECT 182.32 27.1 182.52 27.3 ;
      RECT 182.32 31.18 182.52 31.38 ;
      RECT 182.32 35.26 182.52 35.46 ;
      RECT 182.32 39.34 182.52 39.54 ;
      RECT 182.32 43.42 182.52 43.62 ;
      RECT 182.32 47.5 182.52 47.7 ;
      RECT 182.32 51.58 182.52 51.78 ;
      RECT 182.32 55.66 182.52 55.86 ;
      RECT 182.32 59.74 182.52 59.94 ;
      RECT 180.88 17.58 181.08 17.78 ;
      RECT 180.88 21.66 181.08 21.86 ;
      RECT 180.88 25.74 181.08 25.94 ;
      RECT 180.88 29.82 181.08 30.02 ;
      RECT 180.88 33.9 181.08 34.1 ;
      RECT 180.88 37.98 181.08 38.18 ;
      RECT 180.88 42.06 181.08 42.26 ;
      RECT 180.88 46.14 181.08 46.34 ;
      RECT 180.88 50.22 181.08 50.42 ;
      RECT 180.88 54.3 181.08 54.5 ;
      RECT 180.88 58.38 181.08 58.58 ;
      RECT 180.48 17.58 180.68 17.78 ;
      RECT 180.48 21.66 180.68 21.86 ;
      RECT 180.48 25.74 180.68 25.94 ;
      RECT 180.48 29.82 180.68 30.02 ;
      RECT 180.48 33.9 180.68 34.1 ;
      RECT 180.48 37.98 180.68 38.18 ;
      RECT 180.48 42.06 180.68 42.26 ;
      RECT 180.48 46.14 180.68 46.34 ;
      RECT 180.48 50.22 180.68 50.42 ;
      RECT 180.48 54.3 180.68 54.5 ;
      RECT 180.48 58.38 180.68 58.58 ;
      RECT 177.2 18.94 177.4 19.14 ;
      RECT 177.2 23.02 177.4 23.22 ;
      RECT 177.2 27.1 177.4 27.3 ;
      RECT 177.2 31.18 177.4 31.38 ;
      RECT 177.2 35.26 177.4 35.46 ;
      RECT 177.2 39.34 177.4 39.54 ;
      RECT 177.2 43.42 177.4 43.62 ;
      RECT 177.2 47.5 177.4 47.7 ;
      RECT 177.2 51.58 177.4 51.78 ;
      RECT 177.2 55.66 177.4 55.86 ;
      RECT 177.2 59.74 177.4 59.94 ;
      RECT 176.8 18.94 177 19.14 ;
      RECT 176.8 23.02 177 23.22 ;
      RECT 176.8 27.1 177 27.3 ;
      RECT 176.8 31.18 177 31.38 ;
      RECT 176.8 35.26 177 35.46 ;
      RECT 176.8 39.34 177 39.54 ;
      RECT 176.8 43.42 177 43.62 ;
      RECT 176.8 47.5 177 47.7 ;
      RECT 176.8 51.58 177 51.78 ;
      RECT 176.8 55.66 177 55.86 ;
      RECT 176.8 59.74 177 59.94 ;
      RECT 175.36 17.58 175.56 17.78 ;
      RECT 175.36 21.66 175.56 21.86 ;
      RECT 175.36 25.74 175.56 25.94 ;
      RECT 175.36 29.82 175.56 30.02 ;
      RECT 175.36 33.9 175.56 34.1 ;
      RECT 175.36 37.98 175.56 38.18 ;
      RECT 175.36 42.06 175.56 42.26 ;
      RECT 175.36 46.14 175.56 46.34 ;
      RECT 175.36 50.22 175.56 50.42 ;
      RECT 175.36 54.3 175.56 54.5 ;
      RECT 175.36 58.38 175.56 58.58 ;
      RECT 174.96 17.58 175.16 17.78 ;
      RECT 174.96 21.66 175.16 21.86 ;
      RECT 174.96 25.74 175.16 25.94 ;
      RECT 174.96 29.82 175.16 30.02 ;
      RECT 174.96 33.9 175.16 34.1 ;
      RECT 174.96 37.98 175.16 38.18 ;
      RECT 174.96 42.06 175.16 42.26 ;
      RECT 174.96 46.14 175.16 46.34 ;
      RECT 174.96 50.22 175.16 50.42 ;
      RECT 174.96 54.3 175.16 54.5 ;
      RECT 174.96 58.38 175.16 58.58 ;
      RECT 171.68 18.94 171.88 19.14 ;
      RECT 171.68 23.02 171.88 23.22 ;
      RECT 171.68 27.1 171.88 27.3 ;
      RECT 171.68 31.18 171.88 31.38 ;
      RECT 171.68 35.26 171.88 35.46 ;
      RECT 171.68 39.34 171.88 39.54 ;
      RECT 171.68 43.42 171.88 43.62 ;
      RECT 171.68 47.5 171.88 47.7 ;
      RECT 171.68 51.58 171.88 51.78 ;
      RECT 171.68 55.66 171.88 55.86 ;
      RECT 171.68 59.74 171.88 59.94 ;
      RECT 171.28 18.94 171.48 19.14 ;
      RECT 171.28 23.02 171.48 23.22 ;
      RECT 171.28 27.1 171.48 27.3 ;
      RECT 171.28 31.18 171.48 31.38 ;
      RECT 171.28 35.26 171.48 35.46 ;
      RECT 171.28 39.34 171.48 39.54 ;
      RECT 171.28 43.42 171.48 43.62 ;
      RECT 171.28 47.5 171.48 47.7 ;
      RECT 171.28 51.58 171.48 51.78 ;
      RECT 171.28 55.66 171.48 55.86 ;
      RECT 171.28 59.74 171.48 59.94 ;
      RECT 169.84 17.58 170.04 17.78 ;
      RECT 169.84 21.66 170.04 21.86 ;
      RECT 169.84 25.74 170.04 25.94 ;
      RECT 169.84 29.82 170.04 30.02 ;
      RECT 169.84 33.9 170.04 34.1 ;
      RECT 169.84 37.98 170.04 38.18 ;
      RECT 169.84 42.06 170.04 42.26 ;
      RECT 169.84 46.14 170.04 46.34 ;
      RECT 169.84 50.22 170.04 50.42 ;
      RECT 169.84 54.3 170.04 54.5 ;
      RECT 169.84 58.38 170.04 58.58 ;
      RECT 169.44 17.58 169.64 17.78 ;
      RECT 169.44 21.66 169.64 21.86 ;
      RECT 169.44 25.74 169.64 25.94 ;
      RECT 169.44 29.82 169.64 30.02 ;
      RECT 169.44 33.9 169.64 34.1 ;
      RECT 169.44 37.98 169.64 38.18 ;
      RECT 169.44 42.06 169.64 42.26 ;
      RECT 169.44 46.14 169.64 46.34 ;
      RECT 169.44 50.22 169.64 50.42 ;
      RECT 169.44 54.3 169.64 54.5 ;
      RECT 169.44 58.38 169.64 58.58 ;
      RECT 166.16 18.94 166.36 19.14 ;
      RECT 166.16 23.02 166.36 23.22 ;
      RECT 166.16 27.1 166.36 27.3 ;
      RECT 166.16 31.18 166.36 31.38 ;
      RECT 166.16 35.26 166.36 35.46 ;
      RECT 166.16 39.34 166.36 39.54 ;
      RECT 166.16 43.42 166.36 43.62 ;
      RECT 166.16 47.5 166.36 47.7 ;
      RECT 166.16 51.58 166.36 51.78 ;
      RECT 166.16 55.66 166.36 55.86 ;
      RECT 166.16 59.74 166.36 59.94 ;
      RECT 165.76 18.94 165.96 19.14 ;
      RECT 165.76 23.02 165.96 23.22 ;
      RECT 165.76 27.1 165.96 27.3 ;
      RECT 165.76 31.18 165.96 31.38 ;
      RECT 165.76 35.26 165.96 35.46 ;
      RECT 165.76 39.34 165.96 39.54 ;
      RECT 165.76 43.42 165.96 43.62 ;
      RECT 165.76 47.5 165.96 47.7 ;
      RECT 165.76 51.58 165.96 51.78 ;
      RECT 165.76 55.66 165.96 55.86 ;
      RECT 165.76 59.74 165.96 59.94 ;
      RECT 164.32 17.58 164.52 17.78 ;
      RECT 164.32 21.66 164.52 21.86 ;
      RECT 164.32 25.74 164.52 25.94 ;
      RECT 164.32 29.82 164.52 30.02 ;
      RECT 164.32 33.9 164.52 34.1 ;
      RECT 164.32 37.98 164.52 38.18 ;
      RECT 164.32 42.06 164.52 42.26 ;
      RECT 164.32 46.14 164.52 46.34 ;
      RECT 164.32 50.22 164.52 50.42 ;
      RECT 164.32 54.3 164.52 54.5 ;
      RECT 164.32 58.38 164.52 58.58 ;
      RECT 163.92 17.58 164.12 17.78 ;
      RECT 163.92 21.66 164.12 21.86 ;
      RECT 163.92 25.74 164.12 25.94 ;
      RECT 163.92 29.82 164.12 30.02 ;
      RECT 163.92 33.9 164.12 34.1 ;
      RECT 163.92 37.98 164.12 38.18 ;
      RECT 163.92 42.06 164.12 42.26 ;
      RECT 163.92 46.14 164.12 46.34 ;
      RECT 163.92 50.22 164.12 50.42 ;
      RECT 163.92 54.3 164.12 54.5 ;
      RECT 163.92 58.38 164.12 58.58 ;
      RECT 160.64 18.94 160.84 19.14 ;
      RECT 160.64 23.02 160.84 23.22 ;
      RECT 160.64 27.1 160.84 27.3 ;
      RECT 160.64 31.18 160.84 31.38 ;
      RECT 160.64 35.26 160.84 35.46 ;
      RECT 160.64 39.34 160.84 39.54 ;
      RECT 160.64 43.42 160.84 43.62 ;
      RECT 160.64 47.5 160.84 47.7 ;
      RECT 160.64 51.58 160.84 51.78 ;
      RECT 160.64 55.66 160.84 55.86 ;
      RECT 160.64 59.74 160.84 59.94 ;
      RECT 160.24 18.94 160.44 19.14 ;
      RECT 160.24 23.02 160.44 23.22 ;
      RECT 160.24 27.1 160.44 27.3 ;
      RECT 160.24 31.18 160.44 31.38 ;
      RECT 160.24 35.26 160.44 35.46 ;
      RECT 160.24 39.34 160.44 39.54 ;
      RECT 160.24 43.42 160.44 43.62 ;
      RECT 160.24 47.5 160.44 47.7 ;
      RECT 160.24 51.58 160.44 51.78 ;
      RECT 160.24 55.66 160.44 55.86 ;
      RECT 160.24 59.74 160.44 59.94 ;
      RECT 158.8 17.58 159 17.78 ;
      RECT 158.8 21.66 159 21.86 ;
      RECT 158.8 25.74 159 25.94 ;
      RECT 158.8 29.82 159 30.02 ;
      RECT 158.8 33.9 159 34.1 ;
      RECT 158.8 37.98 159 38.18 ;
      RECT 158.8 42.06 159 42.26 ;
      RECT 158.8 46.14 159 46.34 ;
      RECT 158.8 50.22 159 50.42 ;
      RECT 158.8 54.3 159 54.5 ;
      RECT 158.8 58.38 159 58.58 ;
      RECT 158.4 17.58 158.6 17.78 ;
      RECT 158.4 21.66 158.6 21.86 ;
      RECT 158.4 25.74 158.6 25.94 ;
      RECT 158.4 29.82 158.6 30.02 ;
      RECT 158.4 33.9 158.6 34.1 ;
      RECT 158.4 37.98 158.6 38.18 ;
      RECT 158.4 42.06 158.6 42.26 ;
      RECT 158.4 46.14 158.6 46.34 ;
      RECT 158.4 50.22 158.6 50.42 ;
      RECT 158.4 54.3 158.6 54.5 ;
      RECT 158.4 58.38 158.6 58.58 ;
      RECT 155.12 18.94 155.32 19.14 ;
      RECT 155.12 23.02 155.32 23.22 ;
      RECT 155.12 27.1 155.32 27.3 ;
      RECT 155.12 31.18 155.32 31.38 ;
      RECT 155.12 35.26 155.32 35.46 ;
      RECT 155.12 39.34 155.32 39.54 ;
      RECT 155.12 43.42 155.32 43.62 ;
      RECT 155.12 47.5 155.32 47.7 ;
      RECT 155.12 51.58 155.32 51.78 ;
      RECT 155.12 55.66 155.32 55.86 ;
      RECT 155.12 59.74 155.32 59.94 ;
      RECT 154.72 18.94 154.92 19.14 ;
      RECT 154.72 23.02 154.92 23.22 ;
      RECT 154.72 27.1 154.92 27.3 ;
      RECT 154.72 31.18 154.92 31.38 ;
      RECT 154.72 35.26 154.92 35.46 ;
      RECT 154.72 39.34 154.92 39.54 ;
      RECT 154.72 43.42 154.92 43.62 ;
      RECT 154.72 47.5 154.92 47.7 ;
      RECT 154.72 51.58 154.92 51.78 ;
      RECT 154.72 55.66 154.92 55.86 ;
      RECT 154.72 59.74 154.92 59.94 ;
      RECT 153.28 17.58 153.48 17.78 ;
      RECT 153.28 21.66 153.48 21.86 ;
      RECT 153.28 25.74 153.48 25.94 ;
      RECT 153.28 29.82 153.48 30.02 ;
      RECT 153.28 33.9 153.48 34.1 ;
      RECT 153.28 37.98 153.48 38.18 ;
      RECT 153.28 42.06 153.48 42.26 ;
      RECT 153.28 46.14 153.48 46.34 ;
      RECT 153.28 50.22 153.48 50.42 ;
      RECT 153.28 54.3 153.48 54.5 ;
      RECT 153.28 58.38 153.48 58.58 ;
      RECT 152.88 17.58 153.08 17.78 ;
      RECT 152.88 21.66 153.08 21.86 ;
      RECT 152.88 25.74 153.08 25.94 ;
      RECT 152.88 29.82 153.08 30.02 ;
      RECT 152.88 33.9 153.08 34.1 ;
      RECT 152.88 37.98 153.08 38.18 ;
      RECT 152.88 42.06 153.08 42.26 ;
      RECT 152.88 46.14 153.08 46.34 ;
      RECT 152.88 50.22 153.08 50.42 ;
      RECT 152.88 54.3 153.08 54.5 ;
      RECT 152.88 58.38 153.08 58.58 ;
      RECT 149.6 18.94 149.8 19.14 ;
      RECT 149.6 23.02 149.8 23.22 ;
      RECT 149.6 27.1 149.8 27.3 ;
      RECT 149.6 31.18 149.8 31.38 ;
      RECT 149.6 35.26 149.8 35.46 ;
      RECT 149.6 39.34 149.8 39.54 ;
      RECT 149.6 43.42 149.8 43.62 ;
      RECT 149.6 47.5 149.8 47.7 ;
      RECT 149.6 51.58 149.8 51.78 ;
      RECT 149.6 55.66 149.8 55.86 ;
      RECT 149.6 59.74 149.8 59.94 ;
      RECT 149.2 18.94 149.4 19.14 ;
      RECT 149.2 23.02 149.4 23.22 ;
      RECT 149.2 27.1 149.4 27.3 ;
      RECT 149.2 31.18 149.4 31.38 ;
      RECT 149.2 35.26 149.4 35.46 ;
      RECT 149.2 39.34 149.4 39.54 ;
      RECT 149.2 43.42 149.4 43.62 ;
      RECT 149.2 47.5 149.4 47.7 ;
      RECT 149.2 51.58 149.4 51.78 ;
      RECT 149.2 55.66 149.4 55.86 ;
      RECT 149.2 59.74 149.4 59.94 ;
      RECT 147.76 17.58 147.96 17.78 ;
      RECT 147.76 21.66 147.96 21.86 ;
      RECT 147.76 25.74 147.96 25.94 ;
      RECT 147.76 29.82 147.96 30.02 ;
      RECT 147.76 33.9 147.96 34.1 ;
      RECT 147.76 37.98 147.96 38.18 ;
      RECT 147.76 42.06 147.96 42.26 ;
      RECT 147.76 46.14 147.96 46.34 ;
      RECT 147.76 50.22 147.96 50.42 ;
      RECT 147.76 54.3 147.96 54.5 ;
      RECT 147.76 58.38 147.96 58.58 ;
      RECT 147.36 17.58 147.56 17.78 ;
      RECT 147.36 21.66 147.56 21.86 ;
      RECT 147.36 25.74 147.56 25.94 ;
      RECT 147.36 29.82 147.56 30.02 ;
      RECT 147.36 33.9 147.56 34.1 ;
      RECT 147.36 37.98 147.56 38.18 ;
      RECT 147.36 42.06 147.56 42.26 ;
      RECT 147.36 46.14 147.56 46.34 ;
      RECT 147.36 50.22 147.56 50.42 ;
      RECT 147.36 54.3 147.56 54.5 ;
      RECT 147.36 58.38 147.56 58.58 ;
      RECT 146.18 20.91 146.38 21.11 ;
      RECT 146.18 24.57 146.38 24.77 ;
      RECT 144.08 18.94 144.28 19.14 ;
      RECT 144.08 23.02 144.28 23.22 ;
      RECT 144.08 27.1 144.28 27.3 ;
      RECT 144.08 31.18 144.28 31.38 ;
      RECT 144.08 35.26 144.28 35.46 ;
      RECT 144.08 39.34 144.28 39.54 ;
      RECT 144.08 43.42 144.28 43.62 ;
      RECT 144.08 47.5 144.28 47.7 ;
      RECT 144.08 51.58 144.28 51.78 ;
      RECT 144.08 55.66 144.28 55.86 ;
      RECT 144.08 59.74 144.28 59.94 ;
      RECT 143.68 18.94 143.88 19.14 ;
      RECT 143.68 23.02 143.88 23.22 ;
      RECT 143.68 27.1 143.88 27.3 ;
      RECT 143.68 31.18 143.88 31.38 ;
      RECT 143.68 35.26 143.88 35.46 ;
      RECT 143.68 39.34 143.88 39.54 ;
      RECT 143.68 43.42 143.88 43.62 ;
      RECT 143.68 47.5 143.88 47.7 ;
      RECT 143.68 51.58 143.88 51.78 ;
      RECT 143.68 55.66 143.88 55.86 ;
      RECT 143.68 59.74 143.88 59.94 ;
      RECT 142.24 17.58 142.44 17.78 ;
      RECT 142.24 21.66 142.44 21.86 ;
      RECT 142.24 25.74 142.44 25.94 ;
      RECT 142.24 29.82 142.44 30.02 ;
      RECT 142.24 33.9 142.44 34.1 ;
      RECT 142.24 37.98 142.44 38.18 ;
      RECT 142.24 42.06 142.44 42.26 ;
      RECT 142.24 46.14 142.44 46.34 ;
      RECT 142.24 50.22 142.44 50.42 ;
      RECT 142.24 54.3 142.44 54.5 ;
      RECT 142.24 58.38 142.44 58.58 ;
      RECT 141.84 17.58 142.04 17.78 ;
      RECT 141.84 21.66 142.04 21.86 ;
      RECT 141.84 25.74 142.04 25.94 ;
      RECT 141.84 29.82 142.04 30.02 ;
      RECT 141.84 33.9 142.04 34.1 ;
      RECT 141.84 37.98 142.04 38.18 ;
      RECT 141.84 42.06 142.04 42.26 ;
      RECT 141.84 46.14 142.04 46.34 ;
      RECT 141.84 50.22 142.04 50.42 ;
      RECT 141.84 54.3 142.04 54.5 ;
      RECT 141.84 58.38 142.04 58.58 ;
      RECT 139.97 24.57 140.17 24.77 ;
      RECT 139.97 28.84 140.17 29.04 ;
      RECT 138.56 18.94 138.76 19.14 ;
      RECT 138.56 23.02 138.76 23.22 ;
      RECT 138.56 27.1 138.76 27.3 ;
      RECT 138.56 31.18 138.76 31.38 ;
      RECT 138.56 35.26 138.76 35.46 ;
      RECT 138.56 39.34 138.76 39.54 ;
      RECT 138.56 43.42 138.76 43.62 ;
      RECT 138.56 47.5 138.76 47.7 ;
      RECT 138.56 51.58 138.76 51.78 ;
      RECT 138.56 55.66 138.76 55.86 ;
      RECT 138.56 59.74 138.76 59.94 ;
      RECT 138.16 18.94 138.36 19.14 ;
      RECT 138.16 23.02 138.36 23.22 ;
      RECT 138.16 27.1 138.36 27.3 ;
      RECT 138.16 31.18 138.36 31.38 ;
      RECT 138.16 35.26 138.36 35.46 ;
      RECT 138.16 39.34 138.36 39.54 ;
      RECT 138.16 43.42 138.36 43.62 ;
      RECT 138.16 47.5 138.36 47.7 ;
      RECT 138.16 51.58 138.36 51.78 ;
      RECT 138.16 55.66 138.36 55.86 ;
      RECT 138.16 59.74 138.36 59.94 ;
      RECT 136.72 17.58 136.92 17.78 ;
      RECT 136.72 21.66 136.92 21.86 ;
      RECT 136.72 25.74 136.92 25.94 ;
      RECT 136.72 29.82 136.92 30.02 ;
      RECT 136.72 33.9 136.92 34.1 ;
      RECT 136.72 37.98 136.92 38.18 ;
      RECT 136.72 42.06 136.92 42.26 ;
      RECT 136.72 46.14 136.92 46.34 ;
      RECT 136.72 50.22 136.92 50.42 ;
      RECT 136.72 54.3 136.92 54.5 ;
      RECT 136.72 58.38 136.92 58.58 ;
      RECT 136.32 17.58 136.52 17.78 ;
      RECT 136.32 21.66 136.52 21.86 ;
      RECT 136.32 25.74 136.52 25.94 ;
      RECT 136.32 29.82 136.52 30.02 ;
      RECT 136.32 33.9 136.52 34.1 ;
      RECT 136.32 37.98 136.52 38.18 ;
      RECT 136.32 42.06 136.52 42.26 ;
      RECT 136.32 46.14 136.52 46.34 ;
      RECT 136.32 50.22 136.52 50.42 ;
      RECT 136.32 54.3 136.52 54.5 ;
      RECT 136.32 58.38 136.52 58.58 ;
      RECT 135.14 15.42 135.34 15.62 ;
      RECT 135.14 23.96 135.34 24.16 ;
      RECT 133.04 18.94 133.24 19.14 ;
      RECT 133.04 23.02 133.24 23.22 ;
      RECT 133.04 27.1 133.24 27.3 ;
      RECT 133.04 31.18 133.24 31.38 ;
      RECT 133.04 35.26 133.24 35.46 ;
      RECT 133.04 39.34 133.24 39.54 ;
      RECT 133.04 43.42 133.24 43.62 ;
      RECT 133.04 47.5 133.24 47.7 ;
      RECT 133.04 51.58 133.24 51.78 ;
      RECT 133.04 55.66 133.24 55.86 ;
      RECT 133.04 59.74 133.24 59.94 ;
      RECT 132.64 18.94 132.84 19.14 ;
      RECT 132.64 23.02 132.84 23.22 ;
      RECT 132.64 27.1 132.84 27.3 ;
      RECT 132.64 31.18 132.84 31.38 ;
      RECT 132.64 35.26 132.84 35.46 ;
      RECT 132.64 39.34 132.84 39.54 ;
      RECT 132.64 43.42 132.84 43.62 ;
      RECT 132.64 47.5 132.84 47.7 ;
      RECT 132.64 51.58 132.84 51.78 ;
      RECT 132.64 55.66 132.84 55.86 ;
      RECT 132.64 59.74 132.84 59.94 ;
      RECT 131.2 17.58 131.4 17.78 ;
      RECT 131.2 21.66 131.4 21.86 ;
      RECT 131.2 25.74 131.4 25.94 ;
      RECT 131.2 29.82 131.4 30.02 ;
      RECT 131.2 33.9 131.4 34.1 ;
      RECT 131.2 37.98 131.4 38.18 ;
      RECT 131.2 42.06 131.4 42.26 ;
      RECT 131.2 46.14 131.4 46.34 ;
      RECT 131.2 50.22 131.4 50.42 ;
      RECT 131.2 54.3 131.4 54.5 ;
      RECT 131.2 58.38 131.4 58.58 ;
      RECT 130.8 17.58 131 17.78 ;
      RECT 130.8 21.66 131 21.86 ;
      RECT 130.8 25.74 131 25.94 ;
      RECT 130.8 29.82 131 30.02 ;
      RECT 130.8 33.9 131 34.1 ;
      RECT 130.8 37.98 131 38.18 ;
      RECT 130.8 42.06 131 42.26 ;
      RECT 130.8 46.14 131 46.34 ;
      RECT 130.8 50.22 131 50.42 ;
      RECT 130.8 54.3 131 54.5 ;
      RECT 130.8 58.38 131 58.58 ;
      RECT 127.52 18.94 127.72 19.14 ;
      RECT 127.52 23.02 127.72 23.22 ;
      RECT 127.52 27.1 127.72 27.3 ;
      RECT 127.52 31.18 127.72 31.38 ;
      RECT 127.52 35.26 127.72 35.46 ;
      RECT 127.52 39.34 127.72 39.54 ;
      RECT 127.52 43.42 127.72 43.62 ;
      RECT 127.52 47.5 127.72 47.7 ;
      RECT 127.52 51.58 127.72 51.78 ;
      RECT 127.52 55.66 127.72 55.86 ;
      RECT 127.52 59.74 127.72 59.94 ;
      RECT 127.12 18.94 127.32 19.14 ;
      RECT 127.12 23.02 127.32 23.22 ;
      RECT 127.12 27.1 127.32 27.3 ;
      RECT 127.12 31.18 127.32 31.38 ;
      RECT 127.12 35.26 127.32 35.46 ;
      RECT 127.12 39.34 127.32 39.54 ;
      RECT 127.12 43.42 127.32 43.62 ;
      RECT 127.12 47.5 127.32 47.7 ;
      RECT 127.12 51.58 127.32 51.78 ;
      RECT 127.12 55.66 127.32 55.86 ;
      RECT 127.12 59.74 127.32 59.94 ;
      RECT 125.68 17.58 125.88 17.78 ;
      RECT 125.68 21.66 125.88 21.86 ;
      RECT 125.68 25.74 125.88 25.94 ;
      RECT 125.68 29.82 125.88 30.02 ;
      RECT 125.68 33.9 125.88 34.1 ;
      RECT 125.68 37.98 125.88 38.18 ;
      RECT 125.68 42.06 125.88 42.26 ;
      RECT 125.68 46.14 125.88 46.34 ;
      RECT 125.68 50.22 125.88 50.42 ;
      RECT 125.68 54.3 125.88 54.5 ;
      RECT 125.68 58.38 125.88 58.58 ;
      RECT 125.28 17.58 125.48 17.78 ;
      RECT 125.28 21.66 125.48 21.86 ;
      RECT 125.28 25.74 125.48 25.94 ;
      RECT 125.28 29.82 125.48 30.02 ;
      RECT 125.28 33.9 125.48 34.1 ;
      RECT 125.28 37.98 125.48 38.18 ;
      RECT 125.28 42.06 125.48 42.26 ;
      RECT 125.28 46.14 125.48 46.34 ;
      RECT 125.28 50.22 125.48 50.42 ;
      RECT 125.28 54.3 125.48 54.5 ;
      RECT 125.28 58.38 125.48 58.58 ;
      RECT 122 18.94 122.2 19.14 ;
      RECT 122 23.02 122.2 23.22 ;
      RECT 122 27.1 122.2 27.3 ;
      RECT 122 31.18 122.2 31.38 ;
      RECT 122 35.26 122.2 35.46 ;
      RECT 122 39.34 122.2 39.54 ;
      RECT 122 43.42 122.2 43.62 ;
      RECT 122 47.5 122.2 47.7 ;
      RECT 122 51.58 122.2 51.78 ;
      RECT 122 55.66 122.2 55.86 ;
      RECT 122 59.74 122.2 59.94 ;
      RECT 121.6 18.94 121.8 19.14 ;
      RECT 121.6 23.02 121.8 23.22 ;
      RECT 121.6 27.1 121.8 27.3 ;
      RECT 121.6 31.18 121.8 31.38 ;
      RECT 121.6 35.26 121.8 35.46 ;
      RECT 121.6 39.34 121.8 39.54 ;
      RECT 121.6 43.42 121.8 43.62 ;
      RECT 121.6 47.5 121.8 47.7 ;
      RECT 121.6 51.58 121.8 51.78 ;
      RECT 121.6 55.66 121.8 55.86 ;
      RECT 121.6 59.74 121.8 59.94 ;
      RECT 120.16 17.58 120.36 17.78 ;
      RECT 120.16 21.66 120.36 21.86 ;
      RECT 120.16 25.74 120.36 25.94 ;
      RECT 120.16 29.82 120.36 30.02 ;
      RECT 120.16 33.9 120.36 34.1 ;
      RECT 120.16 37.98 120.36 38.18 ;
      RECT 120.16 42.06 120.36 42.26 ;
      RECT 120.16 46.14 120.36 46.34 ;
      RECT 120.16 50.22 120.36 50.42 ;
      RECT 120.16 54.3 120.36 54.5 ;
      RECT 120.16 58.38 120.36 58.58 ;
      RECT 119.76 17.58 119.96 17.78 ;
      RECT 119.76 21.66 119.96 21.86 ;
      RECT 119.76 25.74 119.96 25.94 ;
      RECT 119.76 29.82 119.96 30.02 ;
      RECT 119.76 33.9 119.96 34.1 ;
      RECT 119.76 37.98 119.96 38.18 ;
      RECT 119.76 42.06 119.96 42.26 ;
      RECT 119.76 46.14 119.96 46.34 ;
      RECT 119.76 50.22 119.96 50.42 ;
      RECT 119.76 54.3 119.96 54.5 ;
      RECT 119.76 58.38 119.96 58.58 ;
      RECT 118.58 20.91 118.78 21.11 ;
      RECT 118.58 28.23 118.78 28.43 ;
      RECT 116.48 18.94 116.68 19.14 ;
      RECT 116.48 23.02 116.68 23.22 ;
      RECT 116.48 27.1 116.68 27.3 ;
      RECT 116.48 31.18 116.68 31.38 ;
      RECT 116.48 35.26 116.68 35.46 ;
      RECT 116.48 39.34 116.68 39.54 ;
      RECT 116.48 43.42 116.68 43.62 ;
      RECT 116.48 47.5 116.68 47.7 ;
      RECT 116.48 51.58 116.68 51.78 ;
      RECT 116.48 55.66 116.68 55.86 ;
      RECT 116.48 59.74 116.68 59.94 ;
      RECT 116.08 18.94 116.28 19.14 ;
      RECT 116.08 23.02 116.28 23.22 ;
      RECT 116.08 27.1 116.28 27.3 ;
      RECT 116.08 31.18 116.28 31.38 ;
      RECT 116.08 35.26 116.28 35.46 ;
      RECT 116.08 39.34 116.28 39.54 ;
      RECT 116.08 43.42 116.28 43.62 ;
      RECT 116.08 47.5 116.28 47.7 ;
      RECT 116.08 51.58 116.28 51.78 ;
      RECT 116.08 55.66 116.28 55.86 ;
      RECT 116.08 59.74 116.28 59.94 ;
      RECT 114.64 17.58 114.84 17.78 ;
      RECT 114.64 21.66 114.84 21.86 ;
      RECT 114.64 25.74 114.84 25.94 ;
      RECT 114.64 29.82 114.84 30.02 ;
      RECT 114.64 33.9 114.84 34.1 ;
      RECT 114.64 37.98 114.84 38.18 ;
      RECT 114.64 42.06 114.84 42.26 ;
      RECT 114.64 46.14 114.84 46.34 ;
      RECT 114.64 50.22 114.84 50.42 ;
      RECT 114.64 54.3 114.84 54.5 ;
      RECT 114.64 58.38 114.84 58.58 ;
      RECT 114.24 17.58 114.44 17.78 ;
      RECT 114.24 21.66 114.44 21.86 ;
      RECT 114.24 25.74 114.44 25.94 ;
      RECT 114.24 29.82 114.44 30.02 ;
      RECT 114.24 33.9 114.44 34.1 ;
      RECT 114.24 37.98 114.44 38.18 ;
      RECT 114.24 42.06 114.44 42.26 ;
      RECT 114.24 46.14 114.44 46.34 ;
      RECT 114.24 50.22 114.44 50.42 ;
      RECT 114.24 54.3 114.44 54.5 ;
      RECT 114.24 58.38 114.44 58.58 ;
      RECT 110.96 18.94 111.16 19.14 ;
      RECT 110.96 23.02 111.16 23.22 ;
      RECT 110.96 27.1 111.16 27.3 ;
      RECT 110.96 31.18 111.16 31.38 ;
      RECT 110.96 35.26 111.16 35.46 ;
      RECT 110.96 39.34 111.16 39.54 ;
      RECT 110.96 43.42 111.16 43.62 ;
      RECT 110.96 47.5 111.16 47.7 ;
      RECT 110.96 51.58 111.16 51.78 ;
      RECT 110.96 55.66 111.16 55.86 ;
      RECT 110.96 59.74 111.16 59.94 ;
      RECT 110.56 18.94 110.76 19.14 ;
      RECT 110.56 23.02 110.76 23.22 ;
      RECT 110.56 27.1 110.76 27.3 ;
      RECT 110.56 31.18 110.76 31.38 ;
      RECT 110.56 35.26 110.76 35.46 ;
      RECT 110.56 39.34 110.76 39.54 ;
      RECT 110.56 43.42 110.76 43.62 ;
      RECT 110.56 47.5 110.76 47.7 ;
      RECT 110.56 51.58 110.76 51.78 ;
      RECT 110.56 55.66 110.76 55.86 ;
      RECT 110.56 59.74 110.76 59.94 ;
      RECT 109.12 17.58 109.32 17.78 ;
      RECT 109.12 21.66 109.32 21.86 ;
      RECT 109.12 25.74 109.32 25.94 ;
      RECT 109.12 29.82 109.32 30.02 ;
      RECT 109.12 33.9 109.32 34.1 ;
      RECT 109.12 37.98 109.32 38.18 ;
      RECT 109.12 42.06 109.32 42.26 ;
      RECT 109.12 46.14 109.32 46.34 ;
      RECT 109.12 50.22 109.32 50.42 ;
      RECT 109.12 54.3 109.32 54.5 ;
      RECT 109.12 58.38 109.32 58.58 ;
      RECT 108.72 17.58 108.92 17.78 ;
      RECT 108.72 21.66 108.92 21.86 ;
      RECT 108.72 25.74 108.92 25.94 ;
      RECT 108.72 29.82 108.92 30.02 ;
      RECT 108.72 33.9 108.92 34.1 ;
      RECT 108.72 37.98 108.92 38.18 ;
      RECT 108.72 42.06 108.92 42.26 ;
      RECT 108.72 46.14 108.92 46.34 ;
      RECT 108.72 50.22 108.92 50.42 ;
      RECT 108.72 54.3 108.92 54.5 ;
      RECT 108.72 58.38 108.92 58.58 ;
      RECT 105.44 18.94 105.64 19.14 ;
      RECT 105.44 23.02 105.64 23.22 ;
      RECT 105.44 27.1 105.64 27.3 ;
      RECT 105.44 31.18 105.64 31.38 ;
      RECT 105.44 35.26 105.64 35.46 ;
      RECT 105.44 39.34 105.64 39.54 ;
      RECT 105.44 43.42 105.64 43.62 ;
      RECT 105.44 47.5 105.64 47.7 ;
      RECT 105.44 51.58 105.64 51.78 ;
      RECT 105.44 55.66 105.64 55.86 ;
      RECT 105.44 59.74 105.64 59.94 ;
      RECT 105.04 18.94 105.24 19.14 ;
      RECT 105.04 23.02 105.24 23.22 ;
      RECT 105.04 27.1 105.24 27.3 ;
      RECT 105.04 31.18 105.24 31.38 ;
      RECT 105.04 35.26 105.24 35.46 ;
      RECT 105.04 39.34 105.24 39.54 ;
      RECT 105.04 43.42 105.24 43.62 ;
      RECT 105.04 47.5 105.24 47.7 ;
      RECT 105.04 51.58 105.24 51.78 ;
      RECT 105.04 55.66 105.24 55.86 ;
      RECT 105.04 59.74 105.24 59.94 ;
      RECT 103.6 17.58 103.8 17.78 ;
      RECT 103.6 21.66 103.8 21.86 ;
      RECT 103.6 25.74 103.8 25.94 ;
      RECT 103.6 29.82 103.8 30.02 ;
      RECT 103.6 33.9 103.8 34.1 ;
      RECT 103.6 37.98 103.8 38.18 ;
      RECT 103.6 42.06 103.8 42.26 ;
      RECT 103.6 46.14 103.8 46.34 ;
      RECT 103.6 50.22 103.8 50.42 ;
      RECT 103.6 54.3 103.8 54.5 ;
      RECT 103.6 58.38 103.8 58.58 ;
      RECT 103.2 17.58 103.4 17.78 ;
      RECT 103.2 21.66 103.4 21.86 ;
      RECT 103.2 25.74 103.4 25.94 ;
      RECT 103.2 29.82 103.4 30.02 ;
      RECT 103.2 33.9 103.4 34.1 ;
      RECT 103.2 37.98 103.4 38.18 ;
      RECT 103.2 42.06 103.4 42.26 ;
      RECT 103.2 46.14 103.4 46.34 ;
      RECT 103.2 50.22 103.4 50.42 ;
      RECT 103.2 54.3 103.4 54.5 ;
      RECT 103.2 58.38 103.4 58.58 ;
      RECT 99.92 18.94 100.12 19.14 ;
      RECT 99.92 23.02 100.12 23.22 ;
      RECT 99.92 27.1 100.12 27.3 ;
      RECT 99.92 31.18 100.12 31.38 ;
      RECT 99.92 35.26 100.12 35.46 ;
      RECT 99.92 39.34 100.12 39.54 ;
      RECT 99.92 43.42 100.12 43.62 ;
      RECT 99.92 47.5 100.12 47.7 ;
      RECT 99.92 51.58 100.12 51.78 ;
      RECT 99.92 55.66 100.12 55.86 ;
      RECT 99.92 59.74 100.12 59.94 ;
      RECT 99.52 18.94 99.72 19.14 ;
      RECT 99.52 23.02 99.72 23.22 ;
      RECT 99.52 27.1 99.72 27.3 ;
      RECT 99.52 31.18 99.72 31.38 ;
      RECT 99.52 35.26 99.72 35.46 ;
      RECT 99.52 39.34 99.72 39.54 ;
      RECT 99.52 43.42 99.72 43.62 ;
      RECT 99.52 47.5 99.72 47.7 ;
      RECT 99.52 51.58 99.72 51.78 ;
      RECT 99.52 55.66 99.72 55.86 ;
      RECT 99.52 59.74 99.72 59.94 ;
      RECT 98.08 17.58 98.28 17.78 ;
      RECT 98.08 21.66 98.28 21.86 ;
      RECT 98.08 25.74 98.28 25.94 ;
      RECT 98.08 29.82 98.28 30.02 ;
      RECT 98.08 33.9 98.28 34.1 ;
      RECT 98.08 37.98 98.28 38.18 ;
      RECT 98.08 42.06 98.28 42.26 ;
      RECT 98.08 46.14 98.28 46.34 ;
      RECT 98.08 50.22 98.28 50.42 ;
      RECT 98.08 54.3 98.28 54.5 ;
      RECT 98.08 58.38 98.28 58.58 ;
      RECT 97.68 17.58 97.88 17.78 ;
      RECT 97.68 21.66 97.88 21.86 ;
      RECT 97.68 25.74 97.88 25.94 ;
      RECT 97.68 29.82 97.88 30.02 ;
      RECT 97.68 33.9 97.88 34.1 ;
      RECT 97.68 37.98 97.88 38.18 ;
      RECT 97.68 42.06 97.88 42.26 ;
      RECT 97.68 46.14 97.88 46.34 ;
      RECT 97.68 50.22 97.88 50.42 ;
      RECT 97.68 54.3 97.88 54.5 ;
      RECT 97.68 58.38 97.88 58.58 ;
      RECT 95.81 16.64 96.01 16.84 ;
      RECT 95.81 20.91 96.01 21.11 ;
      RECT 94.4 18.94 94.6 19.14 ;
      RECT 94.4 23.02 94.6 23.22 ;
      RECT 94.4 27.1 94.6 27.3 ;
      RECT 94.4 31.18 94.6 31.38 ;
      RECT 94.4 35.26 94.6 35.46 ;
      RECT 94.4 39.34 94.6 39.54 ;
      RECT 94.4 43.42 94.6 43.62 ;
      RECT 94.4 47.5 94.6 47.7 ;
      RECT 94.4 51.58 94.6 51.78 ;
      RECT 94.4 55.66 94.6 55.86 ;
      RECT 94.4 59.74 94.6 59.94 ;
      RECT 94 18.94 94.2 19.14 ;
      RECT 94 23.02 94.2 23.22 ;
      RECT 94 27.1 94.2 27.3 ;
      RECT 94 31.18 94.2 31.38 ;
      RECT 94 35.26 94.2 35.46 ;
      RECT 94 39.34 94.2 39.54 ;
      RECT 94 43.42 94.2 43.62 ;
      RECT 94 47.5 94.2 47.7 ;
      RECT 94 51.58 94.2 51.78 ;
      RECT 94 55.66 94.2 55.86 ;
      RECT 94 59.74 94.2 59.94 ;
      RECT 92.56 17.58 92.76 17.78 ;
      RECT 92.56 21.66 92.76 21.86 ;
      RECT 92.56 25.74 92.76 25.94 ;
      RECT 92.56 29.82 92.76 30.02 ;
      RECT 92.56 33.9 92.76 34.1 ;
      RECT 92.56 37.98 92.76 38.18 ;
      RECT 92.56 42.06 92.76 42.26 ;
      RECT 92.56 46.14 92.76 46.34 ;
      RECT 92.56 50.22 92.76 50.42 ;
      RECT 92.56 54.3 92.76 54.5 ;
      RECT 92.56 58.38 92.76 58.58 ;
      RECT 92.16 17.58 92.36 17.78 ;
      RECT 92.16 21.66 92.36 21.86 ;
      RECT 92.16 25.74 92.36 25.94 ;
      RECT 92.16 29.82 92.36 30.02 ;
      RECT 92.16 33.9 92.36 34.1 ;
      RECT 92.16 37.98 92.36 38.18 ;
      RECT 92.16 42.06 92.36 42.26 ;
      RECT 92.16 46.14 92.36 46.34 ;
      RECT 92.16 50.22 92.36 50.42 ;
      RECT 92.16 54.3 92.36 54.5 ;
      RECT 92.16 58.38 92.36 58.58 ;
      RECT 88.88 18.94 89.08 19.14 ;
      RECT 88.88 23.02 89.08 23.22 ;
      RECT 88.88 27.1 89.08 27.3 ;
      RECT 88.88 31.18 89.08 31.38 ;
      RECT 88.88 35.26 89.08 35.46 ;
      RECT 88.88 39.34 89.08 39.54 ;
      RECT 88.88 43.42 89.08 43.62 ;
      RECT 88.88 47.5 89.08 47.7 ;
      RECT 88.88 51.58 89.08 51.78 ;
      RECT 88.88 55.66 89.08 55.86 ;
      RECT 88.88 59.74 89.08 59.94 ;
      RECT 88.48 18.94 88.68 19.14 ;
      RECT 88.48 23.02 88.68 23.22 ;
      RECT 88.48 27.1 88.68 27.3 ;
      RECT 88.48 31.18 88.68 31.38 ;
      RECT 88.48 35.26 88.68 35.46 ;
      RECT 88.48 39.34 88.68 39.54 ;
      RECT 88.48 43.42 88.68 43.62 ;
      RECT 88.48 47.5 88.68 47.7 ;
      RECT 88.48 51.58 88.68 51.78 ;
      RECT 88.48 55.66 88.68 55.86 ;
      RECT 88.48 59.74 88.68 59.94 ;
      RECT 87.04 17.58 87.24 17.78 ;
      RECT 87.04 21.66 87.24 21.86 ;
      RECT 87.04 25.74 87.24 25.94 ;
      RECT 87.04 29.82 87.24 30.02 ;
      RECT 87.04 33.9 87.24 34.1 ;
      RECT 87.04 37.98 87.24 38.18 ;
      RECT 87.04 42.06 87.24 42.26 ;
      RECT 87.04 46.14 87.24 46.34 ;
      RECT 87.04 50.22 87.24 50.42 ;
      RECT 87.04 54.3 87.24 54.5 ;
      RECT 87.04 58.38 87.24 58.58 ;
      RECT 86.64 17.58 86.84 17.78 ;
      RECT 86.64 21.66 86.84 21.86 ;
      RECT 86.64 25.74 86.84 25.94 ;
      RECT 86.64 29.82 86.84 30.02 ;
      RECT 86.64 33.9 86.84 34.1 ;
      RECT 86.64 37.98 86.84 38.18 ;
      RECT 86.64 42.06 86.84 42.26 ;
      RECT 86.64 46.14 86.84 46.34 ;
      RECT 86.64 50.22 86.84 50.42 ;
      RECT 86.64 54.3 86.84 54.5 ;
      RECT 86.64 58.38 86.84 58.58 ;
      RECT 83.36 18.94 83.56 19.14 ;
      RECT 83.36 23.02 83.56 23.22 ;
      RECT 83.36 27.1 83.56 27.3 ;
      RECT 83.36 31.18 83.56 31.38 ;
      RECT 83.36 35.26 83.56 35.46 ;
      RECT 83.36 39.34 83.56 39.54 ;
      RECT 83.36 43.42 83.56 43.62 ;
      RECT 83.36 47.5 83.56 47.7 ;
      RECT 83.36 51.58 83.56 51.78 ;
      RECT 83.36 55.66 83.56 55.86 ;
      RECT 83.36 59.74 83.56 59.94 ;
      RECT 82.96 18.94 83.16 19.14 ;
      RECT 82.96 23.02 83.16 23.22 ;
      RECT 82.96 27.1 83.16 27.3 ;
      RECT 82.96 31.18 83.16 31.38 ;
      RECT 82.96 35.26 83.16 35.46 ;
      RECT 82.96 39.34 83.16 39.54 ;
      RECT 82.96 43.42 83.16 43.62 ;
      RECT 82.96 47.5 83.16 47.7 ;
      RECT 82.96 51.58 83.16 51.78 ;
      RECT 82.96 55.66 83.16 55.86 ;
      RECT 82.96 59.74 83.16 59.94 ;
      RECT 81.52 17.58 81.72 17.78 ;
      RECT 81.52 21.66 81.72 21.86 ;
      RECT 81.52 25.74 81.72 25.94 ;
      RECT 81.52 29.82 81.72 30.02 ;
      RECT 81.52 33.9 81.72 34.1 ;
      RECT 81.52 37.98 81.72 38.18 ;
      RECT 81.52 42.06 81.72 42.26 ;
      RECT 81.52 46.14 81.72 46.34 ;
      RECT 81.52 50.22 81.72 50.42 ;
      RECT 81.52 54.3 81.72 54.5 ;
      RECT 81.52 58.38 81.72 58.58 ;
      RECT 81.12 17.58 81.32 17.78 ;
      RECT 81.12 21.66 81.32 21.86 ;
      RECT 81.12 25.74 81.32 25.94 ;
      RECT 81.12 29.82 81.32 30.02 ;
      RECT 81.12 33.9 81.32 34.1 ;
      RECT 81.12 37.98 81.32 38.18 ;
      RECT 81.12 42.06 81.32 42.26 ;
      RECT 81.12 46.14 81.32 46.34 ;
      RECT 81.12 50.22 81.32 50.42 ;
      RECT 81.12 54.3 81.32 54.5 ;
      RECT 81.12 58.38 81.32 58.58 ;
      RECT 77.84 18.94 78.04 19.14 ;
      RECT 77.84 23.02 78.04 23.22 ;
      RECT 77.84 27.1 78.04 27.3 ;
      RECT 77.84 31.18 78.04 31.38 ;
      RECT 77.84 35.26 78.04 35.46 ;
      RECT 77.84 39.34 78.04 39.54 ;
      RECT 77.84 43.42 78.04 43.62 ;
      RECT 77.84 47.5 78.04 47.7 ;
      RECT 77.84 51.58 78.04 51.78 ;
      RECT 77.84 55.66 78.04 55.86 ;
      RECT 77.84 59.74 78.04 59.94 ;
      RECT 77.44 18.94 77.64 19.14 ;
      RECT 77.44 23.02 77.64 23.22 ;
      RECT 77.44 27.1 77.64 27.3 ;
      RECT 77.44 31.18 77.64 31.38 ;
      RECT 77.44 35.26 77.64 35.46 ;
      RECT 77.44 39.34 77.64 39.54 ;
      RECT 77.44 43.42 77.64 43.62 ;
      RECT 77.44 47.5 77.64 47.7 ;
      RECT 77.44 51.58 77.64 51.78 ;
      RECT 77.44 55.66 77.64 55.86 ;
      RECT 77.44 59.74 77.64 59.94 ;
      RECT 76 17.58 76.2 17.78 ;
      RECT 76 21.66 76.2 21.86 ;
      RECT 76 25.74 76.2 25.94 ;
      RECT 76 29.82 76.2 30.02 ;
      RECT 76 33.9 76.2 34.1 ;
      RECT 76 37.98 76.2 38.18 ;
      RECT 76 42.06 76.2 42.26 ;
      RECT 76 46.14 76.2 46.34 ;
      RECT 76 50.22 76.2 50.42 ;
      RECT 76 54.3 76.2 54.5 ;
      RECT 76 58.38 76.2 58.58 ;
      RECT 75.6 17.58 75.8 17.78 ;
      RECT 75.6 21.66 75.8 21.86 ;
      RECT 75.6 25.74 75.8 25.94 ;
      RECT 75.6 29.82 75.8 30.02 ;
      RECT 75.6 33.9 75.8 34.1 ;
      RECT 75.6 37.98 75.8 38.18 ;
      RECT 75.6 42.06 75.8 42.26 ;
      RECT 75.6 46.14 75.8 46.34 ;
      RECT 75.6 50.22 75.8 50.42 ;
      RECT 75.6 54.3 75.8 54.5 ;
      RECT 75.6 58.38 75.8 58.58 ;
      RECT 74.42 16.64 74.62 16.84 ;
      RECT 74.42 19.69 74.62 19.89 ;
      RECT 72.32 18.94 72.52 19.14 ;
      RECT 72.32 23.02 72.52 23.22 ;
      RECT 72.32 27.1 72.52 27.3 ;
      RECT 72.32 31.18 72.52 31.38 ;
      RECT 72.32 35.26 72.52 35.46 ;
      RECT 72.32 39.34 72.52 39.54 ;
      RECT 72.32 43.42 72.52 43.62 ;
      RECT 72.32 47.5 72.52 47.7 ;
      RECT 72.32 51.58 72.52 51.78 ;
      RECT 72.32 55.66 72.52 55.86 ;
      RECT 72.32 59.74 72.52 59.94 ;
      RECT 71.92 18.94 72.12 19.14 ;
      RECT 71.92 23.02 72.12 23.22 ;
      RECT 71.92 27.1 72.12 27.3 ;
      RECT 71.92 31.18 72.12 31.38 ;
      RECT 71.92 35.26 72.12 35.46 ;
      RECT 71.92 39.34 72.12 39.54 ;
      RECT 71.92 43.42 72.12 43.62 ;
      RECT 71.92 47.5 72.12 47.7 ;
      RECT 71.92 51.58 72.12 51.78 ;
      RECT 71.92 55.66 72.12 55.86 ;
      RECT 71.92 59.74 72.12 59.94 ;
      RECT 70.48 17.58 70.68 17.78 ;
      RECT 70.48 21.66 70.68 21.86 ;
      RECT 70.48 25.74 70.68 25.94 ;
      RECT 70.48 29.82 70.68 30.02 ;
      RECT 70.48 33.9 70.68 34.1 ;
      RECT 70.48 37.98 70.68 38.18 ;
      RECT 70.48 42.06 70.68 42.26 ;
      RECT 70.48 46.14 70.68 46.34 ;
      RECT 70.48 50.22 70.68 50.42 ;
      RECT 70.48 54.3 70.68 54.5 ;
      RECT 70.48 58.38 70.68 58.58 ;
      RECT 70.08 17.58 70.28 17.78 ;
      RECT 70.08 21.66 70.28 21.86 ;
      RECT 70.08 25.74 70.28 25.94 ;
      RECT 70.08 29.82 70.28 30.02 ;
      RECT 70.08 33.9 70.28 34.1 ;
      RECT 70.08 37.98 70.28 38.18 ;
      RECT 70.08 42.06 70.28 42.26 ;
      RECT 70.08 46.14 70.28 46.34 ;
      RECT 70.08 50.22 70.28 50.42 ;
      RECT 70.08 54.3 70.28 54.5 ;
      RECT 70.08 58.38 70.28 58.58 ;
      RECT 66.8 18.94 67 19.14 ;
      RECT 66.8 23.02 67 23.22 ;
      RECT 66.8 27.1 67 27.3 ;
      RECT 66.8 31.18 67 31.38 ;
      RECT 66.8 35.26 67 35.46 ;
      RECT 66.8 39.34 67 39.54 ;
      RECT 66.8 43.42 67 43.62 ;
      RECT 66.8 47.5 67 47.7 ;
      RECT 66.8 51.58 67 51.78 ;
      RECT 66.8 55.66 67 55.86 ;
      RECT 66.8 59.74 67 59.94 ;
      RECT 66.4 18.94 66.6 19.14 ;
      RECT 66.4 23.02 66.6 23.22 ;
      RECT 66.4 27.1 66.6 27.3 ;
      RECT 66.4 31.18 66.6 31.38 ;
      RECT 66.4 35.26 66.6 35.46 ;
      RECT 66.4 39.34 66.6 39.54 ;
      RECT 66.4 43.42 66.6 43.62 ;
      RECT 66.4 47.5 66.6 47.7 ;
      RECT 66.4 51.58 66.6 51.78 ;
      RECT 66.4 55.66 66.6 55.86 ;
      RECT 66.4 59.74 66.6 59.94 ;
      RECT 64.96 17.58 65.16 17.78 ;
      RECT 64.96 21.66 65.16 21.86 ;
      RECT 64.96 25.74 65.16 25.94 ;
      RECT 64.96 29.82 65.16 30.02 ;
      RECT 64.96 33.9 65.16 34.1 ;
      RECT 64.96 37.98 65.16 38.18 ;
      RECT 64.96 42.06 65.16 42.26 ;
      RECT 64.96 46.14 65.16 46.34 ;
      RECT 64.96 50.22 65.16 50.42 ;
      RECT 64.96 54.3 65.16 54.5 ;
      RECT 64.96 58.38 65.16 58.58 ;
      RECT 64.56 17.58 64.76 17.78 ;
      RECT 64.56 21.66 64.76 21.86 ;
      RECT 64.56 25.74 64.76 25.94 ;
      RECT 64.56 29.82 64.76 30.02 ;
      RECT 64.56 33.9 64.76 34.1 ;
      RECT 64.56 37.98 64.76 38.18 ;
      RECT 64.56 42.06 64.76 42.26 ;
      RECT 64.56 46.14 64.76 46.34 ;
      RECT 64.56 50.22 64.76 50.42 ;
      RECT 64.56 54.3 64.76 54.5 ;
      RECT 64.56 58.38 64.76 58.58 ;
      RECT 61.28 18.94 61.48 19.14 ;
      RECT 61.28 23.02 61.48 23.22 ;
      RECT 61.28 27.1 61.48 27.3 ;
      RECT 61.28 31.18 61.48 31.38 ;
      RECT 61.28 35.26 61.48 35.46 ;
      RECT 61.28 39.34 61.48 39.54 ;
      RECT 61.28 43.42 61.48 43.62 ;
      RECT 61.28 47.5 61.48 47.7 ;
      RECT 61.28 51.58 61.48 51.78 ;
      RECT 61.28 55.66 61.48 55.86 ;
      RECT 61.28 59.74 61.48 59.94 ;
      RECT 60.88 18.94 61.08 19.14 ;
      RECT 60.88 23.02 61.08 23.22 ;
      RECT 60.88 27.1 61.08 27.3 ;
      RECT 60.88 31.18 61.08 31.38 ;
      RECT 60.88 35.26 61.08 35.46 ;
      RECT 60.88 39.34 61.08 39.54 ;
      RECT 60.88 43.42 61.08 43.62 ;
      RECT 60.88 47.5 61.08 47.7 ;
      RECT 60.88 51.58 61.08 51.78 ;
      RECT 60.88 55.66 61.08 55.86 ;
      RECT 60.88 59.74 61.08 59.94 ;
      RECT 59.44 17.58 59.64 17.78 ;
      RECT 59.44 21.66 59.64 21.86 ;
      RECT 59.44 25.74 59.64 25.94 ;
      RECT 59.44 29.82 59.64 30.02 ;
      RECT 59.44 33.9 59.64 34.1 ;
      RECT 59.44 37.98 59.64 38.18 ;
      RECT 59.44 42.06 59.64 42.26 ;
      RECT 59.44 46.14 59.64 46.34 ;
      RECT 59.44 50.22 59.64 50.42 ;
      RECT 59.44 54.3 59.64 54.5 ;
      RECT 59.44 58.38 59.64 58.58 ;
      RECT 59.04 17.58 59.24 17.78 ;
      RECT 59.04 21.66 59.24 21.86 ;
      RECT 59.04 25.74 59.24 25.94 ;
      RECT 59.04 29.82 59.24 30.02 ;
      RECT 59.04 33.9 59.24 34.1 ;
      RECT 59.04 37.98 59.24 38.18 ;
      RECT 59.04 42.06 59.24 42.26 ;
      RECT 59.04 46.14 59.24 46.34 ;
      RECT 59.04 50.22 59.24 50.42 ;
      RECT 59.04 54.3 59.24 54.5 ;
      RECT 59.04 58.38 59.24 58.58 ;
      RECT 55.76 18.94 55.96 19.14 ;
      RECT 55.76 23.02 55.96 23.22 ;
      RECT 55.76 27.1 55.96 27.3 ;
      RECT 55.76 31.18 55.96 31.38 ;
      RECT 55.76 35.26 55.96 35.46 ;
      RECT 55.76 39.34 55.96 39.54 ;
      RECT 55.76 43.42 55.96 43.62 ;
      RECT 55.76 47.5 55.96 47.7 ;
      RECT 55.76 51.58 55.96 51.78 ;
      RECT 55.76 55.66 55.96 55.86 ;
      RECT 55.76 59.74 55.96 59.94 ;
      RECT 55.36 18.94 55.56 19.14 ;
      RECT 55.36 23.02 55.56 23.22 ;
      RECT 55.36 27.1 55.56 27.3 ;
      RECT 55.36 31.18 55.56 31.38 ;
      RECT 55.36 35.26 55.56 35.46 ;
      RECT 55.36 39.34 55.56 39.54 ;
      RECT 55.36 43.42 55.56 43.62 ;
      RECT 55.36 47.5 55.56 47.7 ;
      RECT 55.36 51.58 55.56 51.78 ;
      RECT 55.36 55.66 55.56 55.86 ;
      RECT 55.36 59.74 55.56 59.94 ;
      RECT 53.92 17.58 54.12 17.78 ;
      RECT 53.92 21.66 54.12 21.86 ;
      RECT 53.92 25.74 54.12 25.94 ;
      RECT 53.92 29.82 54.12 30.02 ;
      RECT 53.92 33.9 54.12 34.1 ;
      RECT 53.92 37.98 54.12 38.18 ;
      RECT 53.92 42.06 54.12 42.26 ;
      RECT 53.92 46.14 54.12 46.34 ;
      RECT 53.92 50.22 54.12 50.42 ;
      RECT 53.92 54.3 54.12 54.5 ;
      RECT 53.92 58.38 54.12 58.58 ;
      RECT 53.52 17.58 53.72 17.78 ;
      RECT 53.52 21.66 53.72 21.86 ;
      RECT 53.52 25.74 53.72 25.94 ;
      RECT 53.52 29.82 53.72 30.02 ;
      RECT 53.52 33.9 53.72 34.1 ;
      RECT 53.52 37.98 53.72 38.18 ;
      RECT 53.52 42.06 53.72 42.26 ;
      RECT 53.52 46.14 53.72 46.34 ;
      RECT 53.52 50.22 53.72 50.42 ;
      RECT 53.52 54.3 53.72 54.5 ;
      RECT 53.52 58.38 53.72 58.58 ;
      RECT 50.24 18.94 50.44 19.14 ;
      RECT 50.24 23.02 50.44 23.22 ;
      RECT 50.24 27.1 50.44 27.3 ;
      RECT 50.24 31.18 50.44 31.38 ;
      RECT 50.24 35.26 50.44 35.46 ;
      RECT 50.24 39.34 50.44 39.54 ;
      RECT 50.24 43.42 50.44 43.62 ;
      RECT 50.24 47.5 50.44 47.7 ;
      RECT 50.24 51.58 50.44 51.78 ;
      RECT 50.24 55.66 50.44 55.86 ;
      RECT 50.24 59.74 50.44 59.94 ;
      RECT 49.84 18.94 50.04 19.14 ;
      RECT 49.84 23.02 50.04 23.22 ;
      RECT 49.84 27.1 50.04 27.3 ;
      RECT 49.84 31.18 50.04 31.38 ;
      RECT 49.84 35.26 50.04 35.46 ;
      RECT 49.84 39.34 50.04 39.54 ;
      RECT 49.84 43.42 50.04 43.62 ;
      RECT 49.84 47.5 50.04 47.7 ;
      RECT 49.84 51.58 50.04 51.78 ;
      RECT 49.84 55.66 50.04 55.86 ;
      RECT 49.84 59.74 50.04 59.94 ;
      RECT 48.4 17.58 48.6 17.78 ;
      RECT 48.4 21.66 48.6 21.86 ;
      RECT 48.4 25.74 48.6 25.94 ;
      RECT 48.4 29.82 48.6 30.02 ;
      RECT 48.4 33.9 48.6 34.1 ;
      RECT 48.4 37.98 48.6 38.18 ;
      RECT 48.4 42.06 48.6 42.26 ;
      RECT 48.4 46.14 48.6 46.34 ;
      RECT 48.4 50.22 48.6 50.42 ;
      RECT 48.4 54.3 48.6 54.5 ;
      RECT 48.4 58.38 48.6 58.58 ;
      RECT 48 17.58 48.2 17.78 ;
      RECT 48 21.66 48.2 21.86 ;
      RECT 48 25.74 48.2 25.94 ;
      RECT 48 29.82 48.2 30.02 ;
      RECT 48 33.9 48.2 34.1 ;
      RECT 48 37.98 48.2 38.18 ;
      RECT 48 42.06 48.2 42.26 ;
      RECT 48 46.14 48.2 46.34 ;
      RECT 48 50.22 48.2 50.42 ;
      RECT 48 54.3 48.2 54.5 ;
      RECT 48 58.38 48.2 58.58 ;
      RECT 44.72 18.94 44.92 19.14 ;
      RECT 44.72 23.02 44.92 23.22 ;
      RECT 44.72 27.1 44.92 27.3 ;
      RECT 44.72 31.18 44.92 31.38 ;
      RECT 44.72 35.26 44.92 35.46 ;
      RECT 44.72 39.34 44.92 39.54 ;
      RECT 44.72 43.42 44.92 43.62 ;
      RECT 44.72 47.5 44.92 47.7 ;
      RECT 44.72 51.58 44.92 51.78 ;
      RECT 44.72 55.66 44.92 55.86 ;
      RECT 44.72 59.74 44.92 59.94 ;
      RECT 44.32 18.94 44.52 19.14 ;
      RECT 44.32 23.02 44.52 23.22 ;
      RECT 44.32 27.1 44.52 27.3 ;
      RECT 44.32 31.18 44.52 31.38 ;
      RECT 44.32 35.26 44.52 35.46 ;
      RECT 44.32 39.34 44.52 39.54 ;
      RECT 44.32 43.42 44.52 43.62 ;
      RECT 44.32 47.5 44.52 47.7 ;
      RECT 44.32 51.58 44.52 51.78 ;
      RECT 44.32 55.66 44.52 55.86 ;
      RECT 44.32 59.74 44.52 59.94 ;
      RECT 42.88 17.58 43.08 17.78 ;
      RECT 42.88 21.66 43.08 21.86 ;
      RECT 42.88 25.74 43.08 25.94 ;
      RECT 42.88 29.82 43.08 30.02 ;
      RECT 42.88 33.9 43.08 34.1 ;
      RECT 42.88 37.98 43.08 38.18 ;
      RECT 42.88 42.06 43.08 42.26 ;
      RECT 42.88 46.14 43.08 46.34 ;
      RECT 42.88 50.22 43.08 50.42 ;
      RECT 42.88 54.3 43.08 54.5 ;
      RECT 42.88 58.38 43.08 58.58 ;
      RECT 42.48 17.58 42.68 17.78 ;
      RECT 42.48 21.66 42.68 21.86 ;
      RECT 42.48 25.74 42.68 25.94 ;
      RECT 42.48 29.82 42.68 30.02 ;
      RECT 42.48 33.9 42.68 34.1 ;
      RECT 42.48 37.98 42.68 38.18 ;
      RECT 42.48 42.06 42.68 42.26 ;
      RECT 42.48 46.14 42.68 46.34 ;
      RECT 42.48 50.22 42.68 50.42 ;
      RECT 42.48 54.3 42.68 54.5 ;
      RECT 42.48 58.38 42.68 58.58 ;
      RECT 39.2 18.94 39.4 19.14 ;
      RECT 39.2 23.02 39.4 23.22 ;
      RECT 39.2 27.1 39.4 27.3 ;
      RECT 39.2 31.18 39.4 31.38 ;
      RECT 39.2 35.26 39.4 35.46 ;
      RECT 39.2 39.34 39.4 39.54 ;
      RECT 39.2 43.42 39.4 43.62 ;
      RECT 39.2 47.5 39.4 47.7 ;
      RECT 39.2 51.58 39.4 51.78 ;
      RECT 39.2 55.66 39.4 55.86 ;
      RECT 39.2 59.74 39.4 59.94 ;
      RECT 38.8 18.94 39 19.14 ;
      RECT 38.8 23.02 39 23.22 ;
      RECT 38.8 27.1 39 27.3 ;
      RECT 38.8 31.18 39 31.38 ;
      RECT 38.8 35.26 39 35.46 ;
      RECT 38.8 39.34 39 39.54 ;
      RECT 38.8 43.42 39 43.62 ;
      RECT 38.8 47.5 39 47.7 ;
      RECT 38.8 51.58 39 51.78 ;
      RECT 38.8 55.66 39 55.86 ;
      RECT 38.8 59.74 39 59.94 ;
      RECT 37.36 17.58 37.56 17.78 ;
      RECT 37.36 21.66 37.56 21.86 ;
      RECT 37.36 25.74 37.56 25.94 ;
      RECT 37.36 29.82 37.56 30.02 ;
      RECT 37.36 33.9 37.56 34.1 ;
      RECT 37.36 37.98 37.56 38.18 ;
      RECT 37.36 42.06 37.56 42.26 ;
      RECT 37.36 46.14 37.56 46.34 ;
      RECT 37.36 50.22 37.56 50.42 ;
      RECT 37.36 54.3 37.56 54.5 ;
      RECT 37.36 58.38 37.56 58.58 ;
      RECT 36.96 17.58 37.16 17.78 ;
      RECT 36.96 21.66 37.16 21.86 ;
      RECT 36.96 25.74 37.16 25.94 ;
      RECT 36.96 29.82 37.16 30.02 ;
      RECT 36.96 33.9 37.16 34.1 ;
      RECT 36.96 37.98 37.16 38.18 ;
      RECT 36.96 42.06 37.16 42.26 ;
      RECT 36.96 46.14 37.16 46.34 ;
      RECT 36.96 50.22 37.16 50.42 ;
      RECT 36.96 54.3 37.16 54.5 ;
      RECT 36.96 58.38 37.16 58.58 ;
      RECT 33.68 18.94 33.88 19.14 ;
      RECT 33.68 23.02 33.88 23.22 ;
      RECT 33.68 27.1 33.88 27.3 ;
      RECT 33.68 31.18 33.88 31.38 ;
      RECT 33.68 35.26 33.88 35.46 ;
      RECT 33.68 39.34 33.88 39.54 ;
      RECT 33.68 43.42 33.88 43.62 ;
      RECT 33.68 47.5 33.88 47.7 ;
      RECT 33.68 51.58 33.88 51.78 ;
      RECT 33.68 55.66 33.88 55.86 ;
      RECT 33.68 59.74 33.88 59.94 ;
      RECT 33.28 18.94 33.48 19.14 ;
      RECT 33.28 23.02 33.48 23.22 ;
      RECT 33.28 27.1 33.48 27.3 ;
      RECT 33.28 31.18 33.48 31.38 ;
      RECT 33.28 35.26 33.48 35.46 ;
      RECT 33.28 39.34 33.48 39.54 ;
      RECT 33.28 43.42 33.48 43.62 ;
      RECT 33.28 47.5 33.48 47.7 ;
      RECT 33.28 51.58 33.48 51.78 ;
      RECT 33.28 55.66 33.48 55.86 ;
      RECT 33.28 59.74 33.48 59.94 ;
      RECT 31.84 17.58 32.04 17.78 ;
      RECT 31.84 21.66 32.04 21.86 ;
      RECT 31.84 25.74 32.04 25.94 ;
      RECT 31.84 29.82 32.04 30.02 ;
      RECT 31.84 33.9 32.04 34.1 ;
      RECT 31.84 37.98 32.04 38.18 ;
      RECT 31.84 42.06 32.04 42.26 ;
      RECT 31.84 46.14 32.04 46.34 ;
      RECT 31.84 50.22 32.04 50.42 ;
      RECT 31.84 54.3 32.04 54.5 ;
      RECT 31.84 58.38 32.04 58.58 ;
      RECT 31.44 17.58 31.64 17.78 ;
      RECT 31.44 21.66 31.64 21.86 ;
      RECT 31.44 25.74 31.64 25.94 ;
      RECT 31.44 29.82 31.64 30.02 ;
      RECT 31.44 33.9 31.64 34.1 ;
      RECT 31.44 37.98 31.64 38.18 ;
      RECT 31.44 42.06 31.64 42.26 ;
      RECT 31.44 46.14 31.64 46.34 ;
      RECT 31.44 50.22 31.64 50.42 ;
      RECT 31.44 54.3 31.64 54.5 ;
      RECT 31.44 58.38 31.64 58.58 ;
      RECT 28.16 18.94 28.36 19.14 ;
      RECT 28.16 23.02 28.36 23.22 ;
      RECT 28.16 27.1 28.36 27.3 ;
      RECT 28.16 31.18 28.36 31.38 ;
      RECT 28.16 35.26 28.36 35.46 ;
      RECT 28.16 39.34 28.36 39.54 ;
      RECT 28.16 43.42 28.36 43.62 ;
      RECT 28.16 47.5 28.36 47.7 ;
      RECT 28.16 51.58 28.36 51.78 ;
      RECT 28.16 55.66 28.36 55.86 ;
      RECT 28.16 59.74 28.36 59.94 ;
      RECT 27.76 18.94 27.96 19.14 ;
      RECT 27.76 23.02 27.96 23.22 ;
      RECT 27.76 27.1 27.96 27.3 ;
      RECT 27.76 31.18 27.96 31.38 ;
      RECT 27.76 35.26 27.96 35.46 ;
      RECT 27.76 39.34 27.96 39.54 ;
      RECT 27.76 43.42 27.96 43.62 ;
      RECT 27.76 47.5 27.96 47.7 ;
      RECT 27.76 51.58 27.96 51.78 ;
      RECT 27.76 55.66 27.96 55.86 ;
      RECT 27.76 59.74 27.96 59.94 ;
      RECT 26.32 17.58 26.52 17.78 ;
      RECT 26.32 21.66 26.52 21.86 ;
      RECT 26.32 25.74 26.52 25.94 ;
      RECT 26.32 29.82 26.52 30.02 ;
      RECT 26.32 33.9 26.52 34.1 ;
      RECT 26.32 37.98 26.52 38.18 ;
      RECT 26.32 42.06 26.52 42.26 ;
      RECT 26.32 46.14 26.52 46.34 ;
      RECT 26.32 50.22 26.52 50.42 ;
      RECT 26.32 54.3 26.52 54.5 ;
      RECT 26.32 58.38 26.52 58.58 ;
      RECT 25.92 17.58 26.12 17.78 ;
      RECT 25.92 21.66 26.12 21.86 ;
      RECT 25.92 25.74 26.12 25.94 ;
      RECT 25.92 29.82 26.12 30.02 ;
      RECT 25.92 33.9 26.12 34.1 ;
      RECT 25.92 37.98 26.12 38.18 ;
      RECT 25.92 42.06 26.12 42.26 ;
      RECT 25.92 46.14 26.12 46.34 ;
      RECT 25.92 50.22 26.12 50.42 ;
      RECT 25.92 54.3 26.12 54.5 ;
      RECT 25.92 58.38 26.12 58.58 ;
      RECT 22.64 18.94 22.84 19.14 ;
      RECT 22.64 23.02 22.84 23.22 ;
      RECT 22.64 27.1 22.84 27.3 ;
      RECT 22.64 31.18 22.84 31.38 ;
      RECT 22.64 35.26 22.84 35.46 ;
      RECT 22.64 39.34 22.84 39.54 ;
      RECT 22.64 43.42 22.84 43.62 ;
      RECT 22.64 47.5 22.84 47.7 ;
      RECT 22.64 51.58 22.84 51.78 ;
      RECT 22.64 55.66 22.84 55.86 ;
      RECT 22.64 59.74 22.84 59.94 ;
      RECT 22.24 18.94 22.44 19.14 ;
      RECT 22.24 23.02 22.44 23.22 ;
      RECT 22.24 27.1 22.44 27.3 ;
      RECT 22.24 31.18 22.44 31.38 ;
      RECT 22.24 35.26 22.44 35.46 ;
      RECT 22.24 39.34 22.44 39.54 ;
      RECT 22.24 43.42 22.44 43.62 ;
      RECT 22.24 47.5 22.44 47.7 ;
      RECT 22.24 51.58 22.44 51.78 ;
      RECT 22.24 55.66 22.44 55.86 ;
      RECT 22.24 59.74 22.44 59.94 ;
      RECT 20.8 17.58 21 17.78 ;
      RECT 20.8 21.66 21 21.86 ;
      RECT 20.8 25.74 21 25.94 ;
      RECT 20.8 29.82 21 30.02 ;
      RECT 20.8 33.9 21 34.1 ;
      RECT 20.8 37.98 21 38.18 ;
      RECT 20.8 42.06 21 42.26 ;
      RECT 20.8 46.14 21 46.34 ;
      RECT 20.8 50.22 21 50.42 ;
      RECT 20.8 54.3 21 54.5 ;
      RECT 20.8 58.38 21 58.58 ;
      RECT 20.4 17.58 20.6 17.78 ;
      RECT 20.4 21.66 20.6 21.86 ;
      RECT 20.4 25.74 20.6 25.94 ;
      RECT 20.4 29.82 20.6 30.02 ;
      RECT 20.4 33.9 20.6 34.1 ;
      RECT 20.4 37.98 20.6 38.18 ;
      RECT 20.4 42.06 20.6 42.26 ;
      RECT 20.4 46.14 20.6 46.34 ;
      RECT 20.4 50.22 20.6 50.42 ;
      RECT 20.4 54.3 20.6 54.5 ;
      RECT 20.4 58.38 20.6 58.58 ;
    LAYER met4 ;
      RECT 187.67 9.86 188.61 60.18 ;
      RECT 187.43 44.56 188.85 46.56 ;
      RECT 187.43 24.16 188.85 26.16 ;
      RECT 185.83 9.86 186.77 60.18 ;
      RECT 185.59 58.16 187.01 60.16 ;
      RECT 185.59 37.76 187.01 39.76 ;
      RECT 185.59 17.36 187.01 19.36 ;
      RECT 182.15 9.86 183.09 60.18 ;
      RECT 181.91 44.56 183.33 46.56 ;
      RECT 181.91 24.16 183.33 26.16 ;
      RECT 180.31 9.86 181.25 60.18 ;
      RECT 180.07 58.16 181.49 60.16 ;
      RECT 180.07 37.76 181.49 39.76 ;
      RECT 180.07 17.36 181.49 19.36 ;
      RECT 176.63 9.86 177.57 60.18 ;
      RECT 176.39 44.56 177.81 46.56 ;
      RECT 176.39 24.16 177.81 26.16 ;
      RECT 174.79 9.86 175.73 60.18 ;
      RECT 174.55 58.16 175.97 60.16 ;
      RECT 174.55 37.76 175.97 39.76 ;
      RECT 174.55 17.36 175.97 19.36 ;
      RECT 171.11 9.86 172.05 60.18 ;
      RECT 170.87 44.56 172.29 46.56 ;
      RECT 170.87 24.16 172.29 26.16 ;
      RECT 169.27 9.86 170.21 60.18 ;
      RECT 169.03 58.16 170.45 60.16 ;
      RECT 169.03 37.76 170.45 39.76 ;
      RECT 169.03 17.36 170.45 19.36 ;
      RECT 165.59 9.86 166.53 60.18 ;
      RECT 165.35 44.56 166.77 46.56 ;
      RECT 165.35 24.16 166.77 26.16 ;
      RECT 163.75 9.86 164.69 60.18 ;
      RECT 163.51 58.16 164.93 60.16 ;
      RECT 163.51 37.76 164.93 39.76 ;
      RECT 163.51 17.36 164.93 19.36 ;
      RECT 160.07 9.86 161.01 60.18 ;
      RECT 159.83 44.56 161.25 46.56 ;
      RECT 159.83 24.16 161.25 26.16 ;
      RECT 158.23 9.86 159.17 60.18 ;
      RECT 157.99 58.16 159.41 60.16 ;
      RECT 157.99 37.76 159.41 39.76 ;
      RECT 157.99 17.36 159.41 19.36 ;
      RECT 154.55 9.86 155.49 60.18 ;
      RECT 154.31 44.56 155.73 46.56 ;
      RECT 154.31 24.16 155.73 26.16 ;
      RECT 152.71 9.86 153.65 60.18 ;
      RECT 152.47 58.16 153.89 60.16 ;
      RECT 152.47 37.76 153.89 39.76 ;
      RECT 152.47 17.36 153.89 19.36 ;
      RECT 149.03 9.86 149.97 60.18 ;
      RECT 148.79 44.56 150.21 46.56 ;
      RECT 148.79 24.16 150.21 26.16 ;
      RECT 147.19 9.86 148.13 60.18 ;
      RECT 146.95 58.16 148.37 60.16 ;
      RECT 146.95 37.76 148.37 39.76 ;
      RECT 146.95 17.36 148.37 19.36 ;
      RECT 146.115 24.505 146.445 24.835 ;
      RECT 146.13 20.845 146.43 24.835 ;
      RECT 146.115 20.845 146.445 21.175 ;
      RECT 143.51 9.86 144.45 60.18 ;
      RECT 143.27 44.56 144.69 46.56 ;
      RECT 143.27 24.16 144.69 26.16 ;
      RECT 141.67 9.86 142.61 60.18 ;
      RECT 141.43 58.16 142.85 60.16 ;
      RECT 141.43 37.76 142.85 39.76 ;
      RECT 141.43 17.36 142.85 19.36 ;
      RECT 139.905 28.775 140.235 29.105 ;
      RECT 139.92 24.505 140.22 29.105 ;
      RECT 139.905 24.505 140.235 24.835 ;
      RECT 137.99 9.86 138.93 60.18 ;
      RECT 137.75 44.56 139.17 46.56 ;
      RECT 137.75 24.16 139.17 26.16 ;
      RECT 136.15 9.86 137.09 60.18 ;
      RECT 135.91 58.16 137.33 60.16 ;
      RECT 135.91 37.76 137.33 39.76 ;
      RECT 135.91 17.36 137.33 19.36 ;
      RECT 135.075 23.895 135.405 24.225 ;
      RECT 135.09 22.08 135.39 24.225 ;
      RECT 134.4 22.08 135.39 22.38 ;
      RECT 134.4 17.2 134.7 22.38 ;
      RECT 134.4 17.2 135.39 17.5 ;
      RECT 135.09 15.355 135.39 17.5 ;
      RECT 135.075 15.355 135.405 15.685 ;
      RECT 132.47 9.86 133.41 60.18 ;
      RECT 132.23 44.56 133.65 46.56 ;
      RECT 132.23 24.16 133.65 26.16 ;
      RECT 130.63 9.86 131.57 60.18 ;
      RECT 130.39 58.16 131.81 60.16 ;
      RECT 130.39 37.76 131.81 39.76 ;
      RECT 130.39 17.36 131.81 19.36 ;
      RECT 126.95 9.86 127.89 60.18 ;
      RECT 126.71 44.56 128.13 46.56 ;
      RECT 126.71 24.16 128.13 26.16 ;
      RECT 125.11 9.86 126.05 60.18 ;
      RECT 124.87 58.16 126.29 60.16 ;
      RECT 124.87 37.76 126.29 39.76 ;
      RECT 124.87 17.36 126.29 19.36 ;
      RECT 121.43 9.86 122.37 60.18 ;
      RECT 121.19 44.56 122.61 46.56 ;
      RECT 121.19 24.16 122.61 26.16 ;
      RECT 119.59 9.86 120.53 60.18 ;
      RECT 119.35 58.16 120.77 60.16 ;
      RECT 119.35 37.76 120.77 39.76 ;
      RECT 119.35 17.36 120.77 19.36 ;
      RECT 118.515 28.165 118.845 28.495 ;
      RECT 118.53 20.845 118.83 28.495 ;
      RECT 118.515 20.845 118.845 21.175 ;
      RECT 115.91 9.86 116.85 60.18 ;
      RECT 115.67 44.56 117.09 46.56 ;
      RECT 115.67 24.16 117.09 26.16 ;
      RECT 114.07 9.86 115.01 60.18 ;
      RECT 113.83 58.16 115.25 60.16 ;
      RECT 113.83 37.76 115.25 39.76 ;
      RECT 113.83 17.36 115.25 19.36 ;
      RECT 110.39 9.86 111.33 60.18 ;
      RECT 110.15 44.56 111.57 46.56 ;
      RECT 110.15 24.16 111.57 26.16 ;
      RECT 108.55 9.86 109.49 60.18 ;
      RECT 108.31 58.16 109.73 60.16 ;
      RECT 108.31 37.76 109.73 39.76 ;
      RECT 108.31 17.36 109.73 19.36 ;
      RECT 104.87 9.86 105.81 60.18 ;
      RECT 104.63 44.56 106.05 46.56 ;
      RECT 104.63 24.16 106.05 26.16 ;
      RECT 103.03 9.86 103.97 60.18 ;
      RECT 102.79 58.16 104.21 60.16 ;
      RECT 102.79 37.76 104.21 39.76 ;
      RECT 102.79 17.36 104.21 19.36 ;
      RECT 99.35 9.86 100.29 60.18 ;
      RECT 99.11 44.56 100.53 46.56 ;
      RECT 99.11 24.16 100.53 26.16 ;
      RECT 97.51 9.86 98.45 60.18 ;
      RECT 97.27 58.16 98.69 60.16 ;
      RECT 97.27 37.76 98.69 39.76 ;
      RECT 97.27 17.36 98.69 19.36 ;
      RECT 95.745 20.845 96.075 21.175 ;
      RECT 95.76 16.575 96.06 21.175 ;
      RECT 95.745 16.575 96.075 16.905 ;
      RECT 93.83 9.86 94.77 60.18 ;
      RECT 93.59 44.56 95.01 46.56 ;
      RECT 93.59 24.16 95.01 26.16 ;
      RECT 91.99 9.86 92.93 60.18 ;
      RECT 91.75 58.16 93.17 60.16 ;
      RECT 91.75 37.76 93.17 39.76 ;
      RECT 91.75 17.36 93.17 19.36 ;
      RECT 88.31 9.86 89.25 60.18 ;
      RECT 88.07 44.56 89.49 46.56 ;
      RECT 88.07 24.16 89.49 26.16 ;
      RECT 86.47 9.86 87.41 60.18 ;
      RECT 86.23 58.16 87.65 60.16 ;
      RECT 86.23 37.76 87.65 39.76 ;
      RECT 86.23 17.36 87.65 19.36 ;
      RECT 82.79 9.86 83.73 60.18 ;
      RECT 82.55 44.56 83.97 46.56 ;
      RECT 82.55 24.16 83.97 26.16 ;
      RECT 80.95 9.86 81.89 60.18 ;
      RECT 80.71 58.16 82.13 60.16 ;
      RECT 80.71 37.76 82.13 39.76 ;
      RECT 80.71 17.36 82.13 19.36 ;
      RECT 77.27 9.86 78.21 60.18 ;
      RECT 77.03 44.56 78.45 46.56 ;
      RECT 77.03 24.16 78.45 26.16 ;
      RECT 75.43 9.86 76.37 60.18 ;
      RECT 75.19 58.16 76.61 60.16 ;
      RECT 75.19 37.76 76.61 39.76 ;
      RECT 75.19 17.36 76.61 19.36 ;
      RECT 74.355 19.625 74.685 19.955 ;
      RECT 74.37 16.575 74.67 19.955 ;
      RECT 74.355 16.575 74.685 16.905 ;
      RECT 71.75 9.86 72.69 60.18 ;
      RECT 71.51 44.56 72.93 46.56 ;
      RECT 71.51 24.16 72.93 26.16 ;
      RECT 69.91 9.86 70.85 60.18 ;
      RECT 69.67 58.16 71.09 60.16 ;
      RECT 69.67 37.76 71.09 39.76 ;
      RECT 69.67 17.36 71.09 19.36 ;
      RECT 66.23 9.86 67.17 60.18 ;
      RECT 65.99 44.56 67.41 46.56 ;
      RECT 65.99 24.16 67.41 26.16 ;
      RECT 64.39 9.86 65.33 60.18 ;
      RECT 64.15 58.16 65.57 60.16 ;
      RECT 64.15 37.76 65.57 39.76 ;
      RECT 64.15 17.36 65.57 19.36 ;
      RECT 60.71 9.86 61.65 60.18 ;
      RECT 60.47 44.56 61.89 46.56 ;
      RECT 60.47 24.16 61.89 26.16 ;
      RECT 58.87 9.86 59.81 60.18 ;
      RECT 58.63 58.16 60.05 60.16 ;
      RECT 58.63 37.76 60.05 39.76 ;
      RECT 58.63 17.36 60.05 19.36 ;
      RECT 55.19 9.86 56.13 60.18 ;
      RECT 54.95 44.56 56.37 46.56 ;
      RECT 54.95 24.16 56.37 26.16 ;
      RECT 53.35 9.86 54.29 60.18 ;
      RECT 53.11 58.16 54.53 60.16 ;
      RECT 53.11 37.76 54.53 39.76 ;
      RECT 53.11 17.36 54.53 19.36 ;
      RECT 49.67 9.86 50.61 60.18 ;
      RECT 49.43 44.56 50.85 46.56 ;
      RECT 49.43 24.16 50.85 26.16 ;
      RECT 47.83 9.86 48.77 60.18 ;
      RECT 47.59 58.16 49.01 60.16 ;
      RECT 47.59 37.76 49.01 39.76 ;
      RECT 47.59 17.36 49.01 19.36 ;
      RECT 44.15 9.86 45.09 60.18 ;
      RECT 43.91 44.56 45.33 46.56 ;
      RECT 43.91 24.16 45.33 26.16 ;
      RECT 42.31 9.86 43.25 60.18 ;
      RECT 42.07 58.16 43.49 60.16 ;
      RECT 42.07 37.76 43.49 39.76 ;
      RECT 42.07 17.36 43.49 19.36 ;
      RECT 38.63 9.86 39.57 60.18 ;
      RECT 38.39 44.56 39.81 46.56 ;
      RECT 38.39 24.16 39.81 26.16 ;
      RECT 36.79 9.86 37.73 60.18 ;
      RECT 36.55 58.16 37.97 60.16 ;
      RECT 36.55 37.76 37.97 39.76 ;
      RECT 36.55 17.36 37.97 19.36 ;
      RECT 33.11 9.86 34.05 60.18 ;
      RECT 32.87 44.56 34.29 46.56 ;
      RECT 32.87 24.16 34.29 26.16 ;
      RECT 31.27 9.86 32.21 60.18 ;
      RECT 31.03 58.16 32.45 60.16 ;
      RECT 31.03 37.76 32.45 39.76 ;
      RECT 31.03 17.36 32.45 19.36 ;
      RECT 27.59 9.86 28.53 60.18 ;
      RECT 27.35 44.56 28.77 46.56 ;
      RECT 27.35 24.16 28.77 26.16 ;
      RECT 25.75 9.86 26.69 60.18 ;
      RECT 25.51 58.16 26.93 60.16 ;
      RECT 25.51 37.76 26.93 39.76 ;
      RECT 25.51 17.36 26.93 19.36 ;
      RECT 22.07 9.86 23.01 60.18 ;
      RECT 21.83 44.56 23.25 46.56 ;
      RECT 21.83 24.16 23.25 26.16 ;
      RECT 20.23 9.86 21.17 60.18 ;
      RECT 19.99 58.16 21.41 60.16 ;
      RECT 19.99 37.76 21.41 39.76 ;
      RECT 19.99 17.36 21.41 19.36 ;
    LAYER via4 ;
      RECT 187.74 24.76 188.54 25.56 ;
      RECT 187.74 45.16 188.54 45.96 ;
      RECT 185.9 17.96 186.7 18.76 ;
      RECT 185.9 38.36 186.7 39.16 ;
      RECT 185.9 58.76 186.7 59.56 ;
      RECT 182.22 24.76 183.02 25.56 ;
      RECT 182.22 45.16 183.02 45.96 ;
      RECT 180.38 17.96 181.18 18.76 ;
      RECT 180.38 38.36 181.18 39.16 ;
      RECT 180.38 58.76 181.18 59.56 ;
      RECT 176.7 24.76 177.5 25.56 ;
      RECT 176.7 45.16 177.5 45.96 ;
      RECT 174.86 17.96 175.66 18.76 ;
      RECT 174.86 38.36 175.66 39.16 ;
      RECT 174.86 58.76 175.66 59.56 ;
      RECT 171.18 24.76 171.98 25.56 ;
      RECT 171.18 45.16 171.98 45.96 ;
      RECT 169.34 17.96 170.14 18.76 ;
      RECT 169.34 38.36 170.14 39.16 ;
      RECT 169.34 58.76 170.14 59.56 ;
      RECT 165.66 24.76 166.46 25.56 ;
      RECT 165.66 45.16 166.46 45.96 ;
      RECT 163.82 17.96 164.62 18.76 ;
      RECT 163.82 38.36 164.62 39.16 ;
      RECT 163.82 58.76 164.62 59.56 ;
      RECT 160.14 24.76 160.94 25.56 ;
      RECT 160.14 45.16 160.94 45.96 ;
      RECT 158.3 17.96 159.1 18.76 ;
      RECT 158.3 38.36 159.1 39.16 ;
      RECT 158.3 58.76 159.1 59.56 ;
      RECT 154.62 24.76 155.42 25.56 ;
      RECT 154.62 45.16 155.42 45.96 ;
      RECT 152.78 17.96 153.58 18.76 ;
      RECT 152.78 38.36 153.58 39.16 ;
      RECT 152.78 58.76 153.58 59.56 ;
      RECT 149.1 24.76 149.9 25.56 ;
      RECT 149.1 45.16 149.9 45.96 ;
      RECT 147.26 17.96 148.06 18.76 ;
      RECT 147.26 38.36 148.06 39.16 ;
      RECT 147.26 58.76 148.06 59.56 ;
      RECT 143.58 24.76 144.38 25.56 ;
      RECT 143.58 45.16 144.38 45.96 ;
      RECT 141.74 17.96 142.54 18.76 ;
      RECT 141.74 38.36 142.54 39.16 ;
      RECT 141.74 58.76 142.54 59.56 ;
      RECT 138.06 24.76 138.86 25.56 ;
      RECT 138.06 45.16 138.86 45.96 ;
      RECT 136.22 17.96 137.02 18.76 ;
      RECT 136.22 38.36 137.02 39.16 ;
      RECT 136.22 58.76 137.02 59.56 ;
      RECT 132.54 24.76 133.34 25.56 ;
      RECT 132.54 45.16 133.34 45.96 ;
      RECT 130.7 17.96 131.5 18.76 ;
      RECT 130.7 38.36 131.5 39.16 ;
      RECT 130.7 58.76 131.5 59.56 ;
      RECT 127.02 24.76 127.82 25.56 ;
      RECT 127.02 45.16 127.82 45.96 ;
      RECT 125.18 17.96 125.98 18.76 ;
      RECT 125.18 38.36 125.98 39.16 ;
      RECT 125.18 58.76 125.98 59.56 ;
      RECT 121.5 24.76 122.3 25.56 ;
      RECT 121.5 45.16 122.3 45.96 ;
      RECT 119.66 17.96 120.46 18.76 ;
      RECT 119.66 38.36 120.46 39.16 ;
      RECT 119.66 58.76 120.46 59.56 ;
      RECT 115.98 24.76 116.78 25.56 ;
      RECT 115.98 45.16 116.78 45.96 ;
      RECT 114.14 17.96 114.94 18.76 ;
      RECT 114.14 38.36 114.94 39.16 ;
      RECT 114.14 58.76 114.94 59.56 ;
      RECT 110.46 24.76 111.26 25.56 ;
      RECT 110.46 45.16 111.26 45.96 ;
      RECT 108.62 17.96 109.42 18.76 ;
      RECT 108.62 38.36 109.42 39.16 ;
      RECT 108.62 58.76 109.42 59.56 ;
      RECT 104.94 24.76 105.74 25.56 ;
      RECT 104.94 45.16 105.74 45.96 ;
      RECT 103.1 17.96 103.9 18.76 ;
      RECT 103.1 38.36 103.9 39.16 ;
      RECT 103.1 58.76 103.9 59.56 ;
      RECT 99.42 24.76 100.22 25.56 ;
      RECT 99.42 45.16 100.22 45.96 ;
      RECT 97.58 17.96 98.38 18.76 ;
      RECT 97.58 38.36 98.38 39.16 ;
      RECT 97.58 58.76 98.38 59.56 ;
      RECT 93.9 24.76 94.7 25.56 ;
      RECT 93.9 45.16 94.7 45.96 ;
      RECT 92.06 17.96 92.86 18.76 ;
      RECT 92.06 38.36 92.86 39.16 ;
      RECT 92.06 58.76 92.86 59.56 ;
      RECT 88.38 24.76 89.18 25.56 ;
      RECT 88.38 45.16 89.18 45.96 ;
      RECT 86.54 17.96 87.34 18.76 ;
      RECT 86.54 38.36 87.34 39.16 ;
      RECT 86.54 58.76 87.34 59.56 ;
      RECT 82.86 24.76 83.66 25.56 ;
      RECT 82.86 45.16 83.66 45.96 ;
      RECT 81.02 17.96 81.82 18.76 ;
      RECT 81.02 38.36 81.82 39.16 ;
      RECT 81.02 58.76 81.82 59.56 ;
      RECT 77.34 24.76 78.14 25.56 ;
      RECT 77.34 45.16 78.14 45.96 ;
      RECT 75.5 17.96 76.3 18.76 ;
      RECT 75.5 38.36 76.3 39.16 ;
      RECT 75.5 58.76 76.3 59.56 ;
      RECT 71.82 24.76 72.62 25.56 ;
      RECT 71.82 45.16 72.62 45.96 ;
      RECT 69.98 17.96 70.78 18.76 ;
      RECT 69.98 38.36 70.78 39.16 ;
      RECT 69.98 58.76 70.78 59.56 ;
      RECT 66.3 24.76 67.1 25.56 ;
      RECT 66.3 45.16 67.1 45.96 ;
      RECT 64.46 17.96 65.26 18.76 ;
      RECT 64.46 38.36 65.26 39.16 ;
      RECT 64.46 58.76 65.26 59.56 ;
      RECT 60.78 24.76 61.58 25.56 ;
      RECT 60.78 45.16 61.58 45.96 ;
      RECT 58.94 17.96 59.74 18.76 ;
      RECT 58.94 38.36 59.74 39.16 ;
      RECT 58.94 58.76 59.74 59.56 ;
      RECT 55.26 24.76 56.06 25.56 ;
      RECT 55.26 45.16 56.06 45.96 ;
      RECT 53.42 17.96 54.22 18.76 ;
      RECT 53.42 38.36 54.22 39.16 ;
      RECT 53.42 58.76 54.22 59.56 ;
      RECT 49.74 24.76 50.54 25.56 ;
      RECT 49.74 45.16 50.54 45.96 ;
      RECT 47.9 17.96 48.7 18.76 ;
      RECT 47.9 38.36 48.7 39.16 ;
      RECT 47.9 58.76 48.7 59.56 ;
      RECT 44.22 24.76 45.02 25.56 ;
      RECT 44.22 45.16 45.02 45.96 ;
      RECT 42.38 17.96 43.18 18.76 ;
      RECT 42.38 38.36 43.18 39.16 ;
      RECT 42.38 58.76 43.18 59.56 ;
      RECT 38.7 24.76 39.5 25.56 ;
      RECT 38.7 45.16 39.5 45.96 ;
      RECT 36.86 17.96 37.66 18.76 ;
      RECT 36.86 38.36 37.66 39.16 ;
      RECT 36.86 58.76 37.66 59.56 ;
      RECT 33.18 24.76 33.98 25.56 ;
      RECT 33.18 45.16 33.98 45.96 ;
      RECT 31.34 17.96 32.14 18.76 ;
      RECT 31.34 38.36 32.14 39.16 ;
      RECT 31.34 58.76 32.14 59.56 ;
      RECT 27.66 24.76 28.46 25.56 ;
      RECT 27.66 45.16 28.46 45.96 ;
      RECT 25.82 17.96 26.62 18.76 ;
      RECT 25.82 38.36 26.62 39.16 ;
      RECT 25.82 58.76 26.62 59.56 ;
      RECT 22.14 24.76 22.94 25.56 ;
      RECT 22.14 45.16 22.94 45.96 ;
      RECT 20.3 17.96 21.1 18.76 ;
      RECT 20.3 38.36 21.1 39.16 ;
      RECT 20.3 58.76 21.1 59.56 ;
    LAYER met5 ;
      RECT 10.12 17.36 189.98 19.36 ;
      RECT 10.12 24.16 189.98 26.16 ;
      RECT 10.12 37.76 189.98 39.76 ;
      RECT 10.12 44.56 189.98 46.56 ;
      RECT 10.12 58.16 189.98 60.16 ;
    LAYER li1 ;
      RECT 188.455 9.775 188.975 11.575 ;
      RECT 176.035 9.775 176.555 11.575 ;
      RECT 161.315 9.775 161.835 11.575 ;
      RECT 146.595 9.775 147.115 11.575 ;
      RECT 116.235 9.775 116.755 11.575 ;
      RECT 76.675 9.775 77.195 11.575 ;
      RECT 66.555 9.775 67.075 11.575 ;
      RECT 45.395 9.775 45.915 11.575 ;
      RECT 14.115 9.775 14.635 11.575 ;
      RECT 185.905 9.775 187.595 11.555 ;
      RECT 174.425 9.775 175.175 11.555 ;
      RECT 159.705 9.775 160.455 11.555 ;
      RECT 150.495 9.775 153.09 11.555 ;
      RECT 144.985 9.775 145.735 11.555 ;
      RECT 141.295 9.775 143.89 11.555 ;
      RECT 131.185 9.775 132.395 11.555 ;
      RECT 89.785 9.775 90.535 11.555 ;
      RECT 75.065 9.775 75.815 11.555 ;
      RECT 57.585 9.775 58.795 11.555 ;
      RECT 54.345 9.775 56.035 11.555 ;
      RECT 43.325 9.775 44.075 11.555 ;
      RECT 31.805 9.775 33.495 11.555 ;
      RECT 22.625 9.775 23.835 11.555 ;
      RECT 12.045 9.775 13.255 11.555 ;
      RECT 189.605 9.775 189.895 11.11 ;
      RECT 189.145 9.775 189.435 11.11 ;
      RECT 176.725 9.775 177.015 11.11 ;
      RECT 162.005 9.775 162.295 11.11 ;
      RECT 147.285 9.775 147.575 11.11 ;
      RECT 132.565 9.775 132.855 11.11 ;
      RECT 117.845 9.775 118.135 11.11 ;
      RECT 103.125 9.775 103.415 11.11 ;
      RECT 88.405 9.775 88.695 11.11 ;
      RECT 73.685 9.775 73.975 11.11 ;
      RECT 58.965 9.775 59.255 11.11 ;
      RECT 44.245 9.775 44.535 11.11 ;
      RECT 29.525 9.775 29.815 11.11 ;
      RECT 14.805 9.775 15.095 11.11 ;
      RECT 10.205 9.775 10.495 11.11 ;
      RECT 181.815 9.775 182.145 11.095 ;
      RECT 172.615 9.775 172.945 11.095 ;
      RECT 167.095 9.775 167.425 11.095 ;
      RECT 157.895 9.775 158.225 11.095 ;
      RECT 137.655 9.775 137.985 11.095 ;
      RECT 128.915 9.775 129.245 11.095 ;
      RECT 122.935 9.775 123.265 11.095 ;
      RECT 110.415 9.775 110.745 11.095 ;
      RECT 108.215 9.775 108.545 11.095 ;
      RECT 101.775 9.775 102.105 11.095 ;
      RECT 95.335 9.775 95.665 11.095 ;
      RECT 87.515 9.775 87.845 11.095 ;
      RECT 81.995 9.775 82.325 11.095 ;
      RECT 72.795 9.775 73.125 11.095 ;
      RECT 64.975 9.775 65.305 11.095 ;
      RECT 51.635 9.775 51.965 11.095 ;
      RECT 41.515 9.775 41.845 11.095 ;
      RECT 28.635 9.775 28.965 11.095 ;
      RECT 20.355 9.775 20.685 11.095 ;
      RECT 187.765 9.775 188.975 11.035 ;
      RECT 184.085 9.775 187.595 11.035 ;
      RECT 175.345 9.775 176.555 11.035 ;
      RECT 173.505 9.775 175.175 11.035 ;
      RECT 160.625 9.775 161.835 11.035 ;
      RECT 158.785 9.775 160.455 11.035 ;
      RECT 147.745 9.775 153.09 11.035 ;
      RECT 145.905 9.775 147.115 11.035 ;
      RECT 144.065 9.775 145.735 11.035 ;
      RECT 138.545 9.775 143.89 11.035 ;
      RECT 129.805 9.775 132.395 11.035 ;
      RECT 115.545 9.775 116.755 11.035 ;
      RECT 88.865 9.775 90.535 11.035 ;
      RECT 75.985 9.775 77.195 11.035 ;
      RECT 74.145 9.775 75.815 11.035 ;
      RECT 65.865 9.775 67.075 11.035 ;
      RECT 56.205 9.775 58.795 11.035 ;
      RECT 52.525 9.775 56.035 11.035 ;
      RECT 44.705 9.775 45.915 11.035 ;
      RECT 42.405 9.775 44.075 11.035 ;
      RECT 29.985 9.775 33.495 11.035 ;
      RECT 21.245 9.775 23.835 11.035 ;
      RECT 13.425 9.775 14.635 11.035 ;
      RECT 10.665 9.775 13.255 11.035 ;
      RECT 180.975 9.775 181.305 10.745 ;
      RECT 180.135 9.775 180.465 10.745 ;
      RECT 179.295 9.775 179.625 10.745 ;
      RECT 178.535 9.775 178.705 10.745 ;
      RECT 177.695 9.775 177.865 10.745 ;
      RECT 171.775 9.775 172.105 10.745 ;
      RECT 170.935 9.775 171.265 10.745 ;
      RECT 170.095 9.775 170.425 10.745 ;
      RECT 169.335 9.775 169.505 10.745 ;
      RECT 168.495 9.775 168.665 10.745 ;
      RECT 166.255 9.775 166.585 10.745 ;
      RECT 165.415 9.775 165.745 10.745 ;
      RECT 164.575 9.775 164.905 10.745 ;
      RECT 163.815 9.775 163.985 10.745 ;
      RECT 162.975 9.775 163.145 10.745 ;
      RECT 157.055 9.775 157.385 10.745 ;
      RECT 156.215 9.775 156.545 10.745 ;
      RECT 155.375 9.775 155.705 10.745 ;
      RECT 154.615 9.775 154.785 10.745 ;
      RECT 153.775 9.775 153.945 10.745 ;
      RECT 136.815 9.775 137.145 10.745 ;
      RECT 135.975 9.775 136.305 10.745 ;
      RECT 135.135 9.775 135.465 10.745 ;
      RECT 134.375 9.775 134.545 10.745 ;
      RECT 133.535 9.775 133.705 10.745 ;
      RECT 128.075 9.775 128.405 10.745 ;
      RECT 127.235 9.775 127.565 10.745 ;
      RECT 126.395 9.775 126.725 10.745 ;
      RECT 125.635 9.775 125.805 10.745 ;
      RECT 124.795 9.775 124.965 10.745 ;
      RECT 122.095 9.775 122.425 10.745 ;
      RECT 121.255 9.775 121.585 10.745 ;
      RECT 120.415 9.775 120.745 10.745 ;
      RECT 119.655 9.775 119.825 10.745 ;
      RECT 118.815 9.775 118.985 10.745 ;
      RECT 114.695 9.775 114.865 10.745 ;
      RECT 113.855 9.775 114.025 10.745 ;
      RECT 112.935 9.775 113.265 10.745 ;
      RECT 112.095 9.775 112.425 10.745 ;
      RECT 111.255 9.775 111.585 10.745 ;
      RECT 107.375 9.775 107.705 10.745 ;
      RECT 106.535 9.775 106.865 10.745 ;
      RECT 105.695 9.775 106.025 10.745 ;
      RECT 104.935 9.775 105.105 10.745 ;
      RECT 104.095 9.775 104.265 10.745 ;
      RECT 100.935 9.775 101.265 10.745 ;
      RECT 100.095 9.775 100.425 10.745 ;
      RECT 99.255 9.775 99.585 10.745 ;
      RECT 98.495 9.775 98.665 10.745 ;
      RECT 97.655 9.775 97.825 10.745 ;
      RECT 94.495 9.775 94.825 10.745 ;
      RECT 93.655 9.775 93.985 10.745 ;
      RECT 92.815 9.775 93.145 10.745 ;
      RECT 92.055 9.775 92.225 10.745 ;
      RECT 91.215 9.775 91.385 10.745 ;
      RECT 86.675 9.775 87.005 10.745 ;
      RECT 85.835 9.775 86.165 10.745 ;
      RECT 84.995 9.775 85.325 10.745 ;
      RECT 84.235 9.775 84.405 10.745 ;
      RECT 83.395 9.775 83.565 10.745 ;
      RECT 81.155 9.775 81.485 10.745 ;
      RECT 80.315 9.775 80.645 10.745 ;
      RECT 79.475 9.775 79.805 10.745 ;
      RECT 78.715 9.775 78.885 10.745 ;
      RECT 77.875 9.775 78.045 10.745 ;
      RECT 71.955 9.775 72.285 10.745 ;
      RECT 71.115 9.775 71.445 10.745 ;
      RECT 70.275 9.775 70.605 10.745 ;
      RECT 69.515 9.775 69.685 10.745 ;
      RECT 68.675 9.775 68.845 10.745 ;
      RECT 64.135 9.775 64.465 10.745 ;
      RECT 63.295 9.775 63.625 10.745 ;
      RECT 62.455 9.775 62.785 10.745 ;
      RECT 61.695 9.775 61.865 10.745 ;
      RECT 60.855 9.775 61.025 10.745 ;
      RECT 50.795 9.775 51.125 10.745 ;
      RECT 49.955 9.775 50.285 10.745 ;
      RECT 49.115 9.775 49.445 10.745 ;
      RECT 48.355 9.775 48.525 10.745 ;
      RECT 47.515 9.775 47.685 10.745 ;
      RECT 40.675 9.775 41.005 10.745 ;
      RECT 39.835 9.775 40.165 10.745 ;
      RECT 38.995 9.775 39.325 10.745 ;
      RECT 38.235 9.775 38.405 10.745 ;
      RECT 37.395 9.775 37.565 10.745 ;
      RECT 34.155 9.775 34.435 10.745 ;
      RECT 27.795 9.775 28.125 10.745 ;
      RECT 26.955 9.775 27.285 10.745 ;
      RECT 26.115 9.775 26.445 10.745 ;
      RECT 25.355 9.775 25.525 10.745 ;
      RECT 24.515 9.775 24.685 10.745 ;
      RECT 19.515 9.775 19.845 10.745 ;
      RECT 18.675 9.775 19.005 10.745 ;
      RECT 17.835 9.775 18.165 10.745 ;
      RECT 17.075 9.775 17.245 10.745 ;
      RECT 16.235 9.775 16.405 10.745 ;
      RECT 183.145 9.775 183.475 10.705 ;
      RECT 10.12 9.775 189.98 9.945 ;
      RECT 186.385 11.725 187.595 13.955 ;
      RECT 182.705 12.495 184.355 13.955 ;
      RECT 177.185 12.495 179.765 13.955 ;
      RECT 174.885 12.495 175.635 13.955 ;
      RECT 172.125 12.495 173.335 13.955 ;
      RECT 167.985 12.495 169.195 13.955 ;
      RECT 162.465 12.495 165.045 13.955 ;
      RECT 160.625 11.205 161.145 13.955 ;
      RECT 158.785 11.205 159.535 13.955 ;
      RECT 153.265 12.495 155.845 13.955 ;
      RECT 147.745 11.205 150.325 13.955 ;
      RECT 145.905 11.205 146.425 13.955 ;
      RECT 144.065 11.205 144.815 13.955 ;
      RECT 133.025 12.495 135.605 13.955 ;
      RECT 118.305 12.495 118.825 13.955 ;
      RECT 112.785 12.495 113.305 13.955 ;
      RECT 109.105 12.495 110.755 13.955 ;
      RECT 103.585 12.495 106.165 13.955 ;
      RECT 101.745 12.495 102.265 13.955 ;
      RECT 99.905 12.495 100.655 13.955 ;
      RECT 94.385 12.495 96.965 13.955 ;
      RECT 88.865 12.495 91.445 13.955 ;
      RECT 87.025 12.495 87.545 13.955 ;
      RECT 85.185 12.495 85.935 13.955 ;
      RECT 79.665 12.495 82.245 13.955 ;
      RECT 74.145 12.495 76.725 13.955 ;
      RECT 70.925 12.495 72.135 13.955 ;
      RECT 67.245 12.495 68.895 13.955 ;
      RECT 62.185 12.495 62.705 13.955 ;
      RECT 59.425 12.495 60.635 13.955 ;
      RECT 56.205 11.205 57.415 13.955 ;
      RECT 49.765 12.495 50.975 13.955 ;
      RECT 44.705 11.205 45.225 13.955 ;
      RECT 38.725 12.495 41.305 13.955 ;
      RECT 33.665 12.495 34.185 13.955 ;
      RECT 29.985 11.205 31.635 13.955 ;
      RECT 28.145 12.495 28.665 13.955 ;
      RECT 26.305 12.495 27.055 13.955 ;
      RECT 20.785 12.495 23.365 13.955 ;
      RECT 15.265 12.495 17.845 13.955 ;
      RECT 13.425 11.205 13.945 13.955 ;
      RECT 10.665 11.205 11.875 13.955 ;
      RECT 143.175 11.725 143.505 13.465 ;
      RECT 186.385 12.495 188.975 13.435 ;
      RECT 187.765 11.745 188.975 13.435 ;
      RECT 182.705 12.495 186.215 13.435 ;
      RECT 177.185 12.495 182.53 13.435 ;
      RECT 175.345 11.745 176.555 13.435 ;
      RECT 172.125 12.495 174.715 13.435 ;
      RECT 167.985 12.495 170.575 13.435 ;
      RECT 162.465 12.495 167.81 13.435 ;
      RECT 158.785 11.725 160.455 13.435 ;
      RECT 153.265 12.495 158.61 13.435 ;
      RECT 147.745 11.725 153.09 13.435 ;
      RECT 144.065 11.725 145.735 13.435 ;
      RECT 133.025 12.495 138.37 13.435 ;
      RECT 109.105 12.495 112.615 13.435 ;
      RECT 103.585 12.495 108.93 13.435 ;
      RECT 99.905 12.495 101.575 13.435 ;
      RECT 94.385 12.495 99.73 13.435 ;
      RECT 88.865 12.495 94.21 13.435 ;
      RECT 85.185 12.495 86.855 13.435 ;
      RECT 79.665 12.495 85.01 13.435 ;
      RECT 74.145 12.495 79.49 13.435 ;
      RECT 70.925 12.495 73.515 13.435 ;
      RECT 67.245 12.495 70.755 13.435 ;
      RECT 59.425 12.495 62.015 13.435 ;
      RECT 56.205 11.725 58.795 13.435 ;
      RECT 49.765 12.495 52.355 13.435 ;
      RECT 38.725 12.495 44.07 13.435 ;
      RECT 29.985 11.725 33.495 13.435 ;
      RECT 26.305 12.495 27.975 13.435 ;
      RECT 20.785 12.495 26.13 13.435 ;
      RECT 15.265 12.495 20.61 13.435 ;
      RECT 10.665 11.725 13.255 13.435 ;
      RECT 160.625 11.745 161.835 13.415 ;
      RECT 145.905 11.745 147.115 13.415 ;
      RECT 118.305 12.495 119.515 13.415 ;
      RECT 112.785 12.495 113.995 13.415 ;
      RECT 101.745 12.495 102.955 13.415 ;
      RECT 87.025 12.495 88.235 13.415 ;
      RECT 62.185 12.495 63.395 13.415 ;
      RECT 44.705 11.745 45.915 13.415 ;
      RECT 33.665 12.495 34.875 13.415 ;
      RECT 28.145 12.495 29.355 13.415 ;
      RECT 13.425 11.745 14.635 13.415 ;
      RECT 189.605 11.77 189.895 13.39 ;
      RECT 189.145 11.77 189.435 13.39 ;
      RECT 176.725 11.77 177.015 13.39 ;
      RECT 162.005 11.77 162.295 13.39 ;
      RECT 147.285 11.77 147.575 13.39 ;
      RECT 132.565 11.77 132.855 13.39 ;
      RECT 117.845 11.77 118.135 13.39 ;
      RECT 103.125 11.77 103.415 13.39 ;
      RECT 88.405 11.77 88.695 13.39 ;
      RECT 73.685 11.77 73.975 13.39 ;
      RECT 58.965 11.77 59.255 13.39 ;
      RECT 44.245 11.77 44.535 13.39 ;
      RECT 29.525 11.77 29.815 13.39 ;
      RECT 14.805 11.77 15.095 13.39 ;
      RECT 10.205 11.77 10.495 13.39 ;
      RECT 129.45 12.495 129.715 13.19 ;
      RECT 128.59 12.495 128.855 13.19 ;
      RECT 127.73 12.495 127.995 13.19 ;
      RECT 126.87 12.495 127.095 13.19 ;
      RECT 126.01 12.495 126.275 13.19 ;
      RECT 124.985 12.495 125.25 13.19 ;
      RECT 124.1 12.495 124.365 13.19 ;
      RECT 123.24 12.495 123.505 13.19 ;
      RECT 122.375 12.495 122.645 13.19 ;
      RECT 142.335 11.725 142.665 13.145 ;
      RECT 141.495 11.725 141.825 13.145 ;
      RECT 140.655 11.205 140.985 13.145 ;
      RECT 139.815 11.205 140.145 13.145 ;
      RECT 138.975 11.205 139.305 13.145 ;
      RECT 116.855 12.495 117.185 13.145 ;
      RECT 114.595 12.495 114.925 13.145 ;
      RECT 66.255 11.745 66.585 13.145 ;
      RECT 63.995 12.495 64.325 13.145 ;
      RECT 55.275 11.725 55.605 13.145 ;
      RECT 53.015 11.205 53.345 13.145 ;
      RECT 48.775 12.495 49.105 13.145 ;
      RECT 46.515 12.495 46.845 13.145 ;
      RECT 37.735 12.495 38.065 13.145 ;
      RECT 35.475 12.495 35.805 13.145 ;
      RECT 171.185 12.495 171.515 13.045 ;
      RECT 10.12 12.495 189.98 12.665 ;
      RECT 184.085 11.725 187.595 12.665 ;
      RECT 183.145 12.115 183.475 13.955 ;
      RECT 181.815 11.695 182.145 13.435 ;
      RECT 180.975 12.015 181.305 13.435 ;
      RECT 180.135 12.015 180.465 13.435 ;
      RECT 179.295 12.015 179.625 13.955 ;
      RECT 178.455 12.015 178.785 13.955 ;
      RECT 177.615 12.015 177.945 13.955 ;
      RECT 173.505 11.725 175.175 12.665 ;
      RECT 172.615 11.695 172.945 13.955 ;
      RECT 171.775 12.015 172.105 12.665 ;
      RECT 170.935 12.015 171.265 12.665 ;
      RECT 170.095 12.015 170.425 13.435 ;
      RECT 169.255 12.015 169.585 13.435 ;
      RECT 168.415 12.015 168.745 13.955 ;
      RECT 167.095 11.695 167.425 13.435 ;
      RECT 166.255 12.015 166.585 13.435 ;
      RECT 165.415 12.015 165.745 13.435 ;
      RECT 164.575 12.015 164.905 13.955 ;
      RECT 163.735 12.015 164.065 13.955 ;
      RECT 162.895 12.015 163.225 13.955 ;
      RECT 157.895 11.695 158.225 13.435 ;
      RECT 157.055 12.015 157.385 13.435 ;
      RECT 156.215 12.015 156.545 13.435 ;
      RECT 155.375 12.015 155.705 13.955 ;
      RECT 154.535 12.015 154.865 13.955 ;
      RECT 153.695 12.015 154.025 13.955 ;
      RECT 138.545 11.725 143.89 12.665 ;
      RECT 137.655 11.695 137.985 13.435 ;
      RECT 136.815 12.015 137.145 13.435 ;
      RECT 135.975 12.015 136.305 13.435 ;
      RECT 135.135 12.015 135.465 13.955 ;
      RECT 134.295 12.015 134.625 13.955 ;
      RECT 133.455 12.015 133.785 13.955 ;
      RECT 129.805 11.725 132.395 12.665 ;
      RECT 128.915 11.695 129.245 12.665 ;
      RECT 128.075 12.015 128.405 12.665 ;
      RECT 127.235 12.015 127.565 12.665 ;
      RECT 126.395 12.015 126.725 12.665 ;
      RECT 125.555 12.015 125.885 12.665 ;
      RECT 124.715 12.015 125.045 12.665 ;
      RECT 122.935 11.695 123.265 12.665 ;
      RECT 122.095 12.015 122.425 12.665 ;
      RECT 121.255 12.015 121.585 12.665 ;
      RECT 120.415 12.015 120.745 12.665 ;
      RECT 119.575 12.015 119.905 12.665 ;
      RECT 118.735 12.015 119.065 13.415 ;
      RECT 115.545 11.745 116.755 12.665 ;
      RECT 114.615 12.015 114.945 12.665 ;
      RECT 113.775 12.015 114.105 12.665 ;
      RECT 112.935 12.015 113.265 13.955 ;
      RECT 112.095 12.015 112.425 13.435 ;
      RECT 111.255 12.015 111.585 13.435 ;
      RECT 110.415 11.695 110.745 13.955 ;
      RECT 108.215 11.695 108.545 13.435 ;
      RECT 107.375 12.015 107.705 13.435 ;
      RECT 106.535 12.015 106.865 13.435 ;
      RECT 105.695 12.015 106.025 13.955 ;
      RECT 104.855 12.015 105.185 13.955 ;
      RECT 104.015 12.015 104.345 13.955 ;
      RECT 101.775 11.695 102.105 13.955 ;
      RECT 100.935 12.015 101.265 13.435 ;
      RECT 100.095 12.015 100.425 13.955 ;
      RECT 99.255 12.015 99.585 13.435 ;
      RECT 98.415 12.015 98.745 13.435 ;
      RECT 97.575 12.015 97.905 13.435 ;
      RECT 95.335 11.695 95.665 13.955 ;
      RECT 94.495 12.015 94.825 13.955 ;
      RECT 93.655 12.015 93.985 13.435 ;
      RECT 92.815 12.015 93.145 13.435 ;
      RECT 91.975 12.015 92.305 13.435 ;
      RECT 91.135 12.015 91.465 13.435 ;
      RECT 88.865 11.725 90.535 13.955 ;
      RECT 87.515 11.695 87.845 13.415 ;
      RECT 86.675 12.015 87.005 12.665 ;
      RECT 85.835 12.015 86.165 13.435 ;
      RECT 84.995 12.015 85.325 12.665 ;
      RECT 84.155 12.015 84.485 13.435 ;
      RECT 83.315 12.015 83.645 13.435 ;
      RECT 81.995 11.695 82.325 13.435 ;
      RECT 81.155 12.015 81.485 13.955 ;
      RECT 80.315 12.015 80.645 13.955 ;
      RECT 79.475 12.015 79.805 12.665 ;
      RECT 78.635 12.015 78.965 13.435 ;
      RECT 77.795 12.015 78.125 13.435 ;
      RECT 75.985 11.745 77.195 13.435 ;
      RECT 74.145 11.725 75.815 13.955 ;
      RECT 72.795 11.695 73.125 13.435 ;
      RECT 71.955 12.015 72.285 13.435 ;
      RECT 71.115 12.015 71.445 13.955 ;
      RECT 70.275 12.015 70.605 13.435 ;
      RECT 69.435 12.015 69.765 13.435 ;
      RECT 68.595 12.015 68.925 13.435 ;
      RECT 65.865 11.745 67.075 12.665 ;
      RECT 64.975 11.695 65.305 12.665 ;
      RECT 64.135 12.015 64.465 12.665 ;
      RECT 63.295 12.015 63.625 12.665 ;
      RECT 62.455 12.015 62.785 13.415 ;
      RECT 61.615 12.015 61.945 13.435 ;
      RECT 60.775 12.015 61.105 13.435 ;
      RECT 52.525 11.725 56.035 12.665 ;
      RECT 51.635 11.695 51.965 13.435 ;
      RECT 50.795 12.015 51.125 13.435 ;
      RECT 49.955 12.015 50.285 13.955 ;
      RECT 49.115 12.015 49.445 12.665 ;
      RECT 48.275 12.015 48.605 12.665 ;
      RECT 47.435 12.015 47.765 12.665 ;
      RECT 42.405 11.725 44.075 12.665 ;
      RECT 41.515 11.695 41.845 13.435 ;
      RECT 40.675 12.015 41.005 13.955 ;
      RECT 39.835 12.015 40.165 13.955 ;
      RECT 38.995 12.015 39.325 13.955 ;
      RECT 38.155 12.015 38.485 12.665 ;
      RECT 37.315 12.015 37.645 12.665 ;
      RECT 35.025 12.095 35.355 12.665 ;
      RECT 34.135 12.095 34.515 13.415 ;
      RECT 28.635 11.695 28.965 13.415 ;
      RECT 27.795 12.015 28.125 12.665 ;
      RECT 26.955 12.015 27.285 13.435 ;
      RECT 26.115 12.015 26.445 12.665 ;
      RECT 25.275 12.015 25.605 13.435 ;
      RECT 24.435 12.015 24.765 13.435 ;
      RECT 21.245 11.725 23.835 13.435 ;
      RECT 20.355 11.695 20.685 12.665 ;
      RECT 19.515 12.015 19.845 13.435 ;
      RECT 18.675 12.015 19.005 13.435 ;
      RECT 17.835 12.015 18.165 13.435 ;
      RECT 16.995 12.015 17.325 13.955 ;
      RECT 16.155 12.015 16.485 13.955 ;
      RECT 187.765 11.205 188.285 13.435 ;
      RECT 175.345 11.205 175.865 13.435 ;
      RECT 115.545 11.205 116.065 12.665 ;
      RECT 75.985 11.205 76.505 13.955 ;
      RECT 65.865 11.205 66.385 12.665 ;
      RECT 184.085 11.205 185.735 13.435 ;
      RECT 173.505 11.205 174.255 13.435 ;
      RECT 138.545 11.205 141.125 12.665 ;
      RECT 129.805 11.205 131.015 12.665 ;
      RECT 88.865 11.205 89.615 13.955 ;
      RECT 74.145 11.205 74.895 13.955 ;
      RECT 52.525 11.205 54.175 12.665 ;
      RECT 42.405 11.205 43.155 13.435 ;
      RECT 21.245 11.205 22.455 13.955 ;
      RECT 176.035 13.605 176.555 17.015 ;
      RECT 161.315 13.585 161.835 17.015 ;
      RECT 146.595 13.585 147.115 17.015 ;
      RECT 131.875 15.215 132.395 17.015 ;
      RECT 117.155 15.215 117.675 17.015 ;
      RECT 93.235 13.605 93.755 17.015 ;
      RECT 80.355 14.125 80.875 17.015 ;
      RECT 60.115 14.125 60.635 17.015 ;
      RECT 50.915 14.125 51.435 17.015 ;
      RECT 32.515 13.605 33.035 17.015 ;
      RECT 28.835 13.585 29.355 17.015 ;
      RECT 14.115 13.585 14.635 17.015 ;
      RECT 188.225 13.605 188.975 16.995 ;
      RECT 185.925 15.215 187.135 16.995 ;
      RECT 174.425 15.215 175.175 16.995 ;
      RECT 157.855 15.215 160.45 16.995 ;
      RECT 143.135 15.215 145.73 16.995 ;
      RECT 128.415 15.215 131.01 16.995 ;
      RECT 111.865 13.605 112.615 16.995 ;
      RECT 102.205 14.125 102.955 16.995 ;
      RECT 102.435 13.585 102.955 16.995 ;
      RECT 90.685 14.125 92.375 16.995 ;
      RECT 76.895 13.605 79.49 16.995 ;
      RECT 47.455 15.215 50.05 16.995 ;
      RECT 42.385 15.215 44.075 16.995 ;
      RECT 30.905 14.125 31.655 16.995 ;
      RECT 27.225 13.605 27.975 16.995 ;
      RECT 23.535 13.605 26.13 16.995 ;
      RECT 18.015 13.605 20.61 16.995 ;
      RECT 12.045 13.605 13.255 16.995 ;
      RECT 189.605 14.05 189.895 16.55 ;
      RECT 189.145 14.05 189.435 16.55 ;
      RECT 176.725 14.05 177.015 16.55 ;
      RECT 162.005 14.05 162.295 16.55 ;
      RECT 147.285 14.05 147.575 16.55 ;
      RECT 132.565 14.05 132.855 16.55 ;
      RECT 117.845 14.05 118.135 16.55 ;
      RECT 103.125 14.05 103.415 16.55 ;
      RECT 88.405 14.05 88.695 16.55 ;
      RECT 73.685 14.05 73.975 16.55 ;
      RECT 58.965 14.05 59.255 16.55 ;
      RECT 44.245 14.05 44.535 16.55 ;
      RECT 29.525 14.05 29.815 16.55 ;
      RECT 14.805 14.05 15.095 16.55 ;
      RECT 10.205 14.05 10.495 16.55 ;
      RECT 61.195 13.605 61.525 16.535 ;
      RECT 187.305 14.125 188.975 16.475 ;
      RECT 187.765 13.605 188.975 16.475 ;
      RECT 184.545 15.215 187.135 16.475 ;
      RECT 175.345 14.125 176.555 16.475 ;
      RECT 175.805 13.605 176.555 16.475 ;
      RECT 173.505 13.605 174.715 16.475 ;
      RECT 160.625 14.125 161.835 16.475 ;
      RECT 155.105 15.215 160.45 16.475 ;
      RECT 156.015 13.605 158.61 16.475 ;
      RECT 145.905 14.125 147.115 16.475 ;
      RECT 140.385 15.215 145.73 16.475 ;
      RECT 131.185 15.215 132.395 16.475 ;
      RECT 125.665 15.215 131.01 16.475 ;
      RECT 116.465 15.215 117.675 16.475 ;
      RECT 116.9 14.455 117.23 16.475 ;
      RECT 110.945 13.605 112.615 16.475 ;
      RECT 101.285 15.215 102.955 16.475 ;
      RECT 101.745 14.125 102.955 16.475 ;
      RECT 92.545 13.605 93.755 16.475 ;
      RECT 88.865 14.125 92.375 16.475 ;
      RECT 79.665 14.125 80.875 16.475 ;
      RECT 74.145 14.125 79.49 16.475 ;
      RECT 59.425 14.125 60.635 16.475 ;
      RECT 50.225 14.125 51.435 16.475 ;
      RECT 44.705 15.215 50.05 16.475 ;
      RECT 40.565 15.215 44.075 16.475 ;
      RECT 41.475 13.605 44.07 16.475 ;
      RECT 31.825 13.605 33.035 16.475 ;
      RECT 29.985 14.125 31.655 16.475 ;
      RECT 28.145 14.125 29.355 16.475 ;
      RECT 26.305 14.125 27.975 16.475 ;
      RECT 20.785 14.125 26.13 16.475 ;
      RECT 15.265 14.125 20.61 16.475 ;
      RECT 13.425 14.125 14.635 16.475 ;
      RECT 10.665 14.125 13.255 16.475 ;
      RECT 183.645 14.125 183.815 16.395 ;
      RECT 168.925 14.125 169.095 16.395 ;
      RECT 154.205 14.125 154.375 16.395 ;
      RECT 139.485 15.215 139.655 16.395 ;
      RECT 124.765 15.215 124.935 16.395 ;
      RECT 110.045 14.125 110.215 16.395 ;
      RECT 100.385 14.125 100.555 16.395 ;
      RECT 87.505 14.125 87.675 16.395 ;
      RECT 72.785 13.605 72.955 16.395 ;
      RECT 58.065 13.605 58.235 16.395 ;
      RECT 39.665 14.125 39.835 16.395 ;
      RECT 180.71 13.605 180.88 16.185 ;
      RECT 165.99 13.605 166.16 16.185 ;
      RECT 151.27 13.605 151.44 16.185 ;
      RECT 136.55 13.605 136.72 16.185 ;
      RECT 121.83 15.215 122 16.185 ;
      RECT 107.11 13.605 107.28 16.185 ;
      RECT 97.45 13.605 97.62 16.185 ;
      RECT 84.57 13.605 84.74 16.185 ;
      RECT 69.85 13.605 70.02 16.185 ;
      RECT 65.475 14.795 65.645 16.185 ;
      RECT 64.635 15.215 64.805 16.185 ;
      RECT 63.715 15.215 64.045 16.185 ;
      RECT 62.875 13.585 63.205 16.185 ;
      RECT 62.035 15.215 62.365 16.185 ;
      RECT 55.13 15.215 55.3 16.185 ;
      RECT 36.73 15.215 36.9 16.185 ;
      RECT 115.52 15.215 115.85 16.145 ;
      RECT 182.59 15.215 182.905 15.885 ;
      RECT 177.615 14.125 177.945 15.885 ;
      RECT 167.87 15.215 168.185 15.885 ;
      RECT 162.895 14.125 163.225 15.885 ;
      RECT 153.15 15.215 153.465 15.885 ;
      RECT 148.175 14.125 148.505 15.885 ;
      RECT 138.43 15.215 138.745 15.885 ;
      RECT 133.455 14.125 133.785 15.885 ;
      RECT 123.71 15.215 124.025 15.885 ;
      RECT 118.735 14.125 119.065 15.885 ;
      RECT 108.99 15.215 109.305 15.885 ;
      RECT 104.015 14.125 104.345 15.885 ;
      RECT 99.33 13.605 99.645 15.885 ;
      RECT 94.355 15.215 94.685 15.885 ;
      RECT 86.45 13.605 86.765 15.885 ;
      RECT 81.475 14.125 81.805 15.885 ;
      RECT 71.73 14.125 72.045 15.885 ;
      RECT 66.755 15.215 67.085 15.885 ;
      RECT 57.01 14.125 57.325 15.885 ;
      RECT 52.035 15.215 52.365 15.885 ;
      RECT 38.61 15.215 38.925 15.885 ;
      RECT 33.635 15.215 33.965 15.885 ;
      RECT 178.54 14.125 178.805 15.845 ;
      RECT 172.275 14.125 172.6 15.845 ;
      RECT 170.855 15.215 171.125 15.845 ;
      RECT 163.82 14.125 164.085 15.845 ;
      RECT 149.1 14.125 149.365 15.845 ;
      RECT 134.38 14.125 134.645 15.845 ;
      RECT 119.66 15.215 119.925 15.845 ;
      RECT 104.94 14.125 105.205 15.845 ;
      RECT 95.28 14.125 95.545 15.845 ;
      RECT 82.4 14.125 82.665 15.845 ;
      RECT 67.68 14.125 67.945 15.845 ;
      RECT 52.96 15.215 53.225 15.845 ;
      RECT 34.56 13.585 34.825 15.845 ;
      RECT 114.575 15.215 114.93 15.805 ;
      RECT 10.12 15.215 189.98 15.385 ;
      RECT 186.385 14.125 188.975 15.385 ;
      RECT 182.705 14.125 186.215 15.385 ;
      RECT 184.525 13.605 186.215 15.385 ;
      RECT 177.185 14.125 182.53 15.385 ;
      RECT 179.935 13.605 182.53 15.385 ;
      RECT 174.885 14.125 176.555 15.385 ;
      RECT 172.125 14.125 174.715 15.385 ;
      RECT 171.185 14.455 171.515 15.385 ;
      RECT 167.985 14.125 170.575 15.385 ;
      RECT 169.365 13.605 170.575 15.385 ;
      RECT 162.465 14.125 167.81 15.385 ;
      RECT 165.215 13.605 167.81 15.385 ;
      RECT 158.785 14.125 160.455 15.385 ;
      RECT 159.705 13.605 160.455 15.385 ;
      RECT 153.265 14.125 158.61 15.385 ;
      RECT 147.745 14.125 153.09 15.385 ;
      RECT 150.495 13.605 153.09 15.385 ;
      RECT 144.065 14.125 145.735 15.385 ;
      RECT 144.985 13.605 145.735 15.385 ;
      RECT 143.175 14.065 143.505 16.995 ;
      RECT 142.335 14.415 142.665 16.475 ;
      RECT 141.495 14.415 141.825 16.475 ;
      RECT 140.655 14.415 140.985 16.475 ;
      RECT 139.895 14.415 140.065 15.385 ;
      RECT 139.055 14.415 139.225 15.385 ;
      RECT 133.025 14.125 138.37 15.385 ;
      RECT 135.775 13.605 138.37 15.385 ;
      RECT 131.17 14.415 131.43 15.385 ;
      RECT 130.315 14.415 130.57 16.995 ;
      RECT 129.455 14.415 129.71 16.995 ;
      RECT 128.595 14.415 128.85 16.995 ;
      RECT 127.735 14.415 127.99 16.475 ;
      RECT 126.875 14.415 127.13 16.475 ;
      RECT 126.01 14.7 126.27 16.475 ;
      RECT 124.985 14.415 125.24 15.385 ;
      RECT 124.105 14.415 124.36 15.385 ;
      RECT 123.24 14.415 123.5 15.385 ;
      RECT 122.385 14.415 122.64 15.385 ;
      RECT 121.52 14.415 121.78 15.385 ;
      RECT 120.66 14.075 120.925 15.385 ;
      RECT 118.305 14.125 119.515 15.385 ;
      RECT 118.995 13.585 119.515 15.385 ;
      RECT 115.955 14.795 116.31 15.385 ;
      RECT 112.785 14.125 113.995 15.385 ;
      RECT 113.475 13.585 113.995 15.385 ;
      RECT 109.105 14.125 112.615 15.385 ;
      RECT 110.925 13.605 112.615 15.385 ;
      RECT 103.585 14.125 108.93 15.385 ;
      RECT 106.335 13.605 108.93 15.385 ;
      RECT 99.905 14.125 101.575 15.385 ;
      RECT 94.385 14.125 99.73 15.385 ;
      RECT 97.135 13.605 99.73 15.385 ;
      RECT 91.615 13.605 94.21 15.385 ;
      RECT 87.025 14.125 88.235 15.385 ;
      RECT 87.715 13.585 88.235 15.385 ;
      RECT 85.185 14.125 86.855 15.385 ;
      RECT 86.105 13.605 86.855 15.385 ;
      RECT 79.665 14.125 85.01 15.385 ;
      RECT 82.415 13.605 85.01 15.385 ;
      RECT 70.925 14.125 73.515 15.385 ;
      RECT 72.305 13.605 73.515 15.385 ;
      RECT 67.245 14.125 70.755 15.385 ;
      RECT 69.065 13.605 70.755 15.385 ;
      RECT 66.3 14.455 66.63 15.385 ;
      RECT 65.355 14.795 65.71 15.385 ;
      RECT 62.185 14.125 63.395 15.385 ;
      RECT 62.875 13.585 63.395 15.385 ;
      RECT 59.425 14.125 62.015 15.385 ;
      RECT 60.805 13.605 62.015 15.385 ;
      RECT 56.205 14.125 58.795 15.385 ;
      RECT 57.585 13.605 58.795 15.385 ;
      RECT 53.89 14.795 54.245 15.385 ;
      RECT 52.97 14.455 53.3 15.385 ;
      RECT 49.765 14.125 52.355 15.385 ;
      RECT 48.82 14.455 49.15 16.995 ;
      RECT 47.875 14.795 48.23 16.995 ;
      RECT 44.705 14.125 45.915 16.475 ;
      RECT 45.395 13.585 45.915 16.475 ;
      RECT 38.725 14.125 44.07 15.385 ;
      RECT 37.78 14.455 38.11 15.385 ;
      RECT 36.835 14.795 37.19 15.385 ;
      RECT 33.665 14.125 34.875 15.385 ;
      RECT 34.355 13.585 34.875 15.385 ;
      RECT 29.985 14.125 33.495 15.385 ;
      RECT 31.805 13.605 33.495 15.385 ;
      RECT 126.01 14.415 126.265 16.475 ;
      RECT 100.825 13.605 101.575 15.385 ;
      RECT 51.145 13.605 52.355 15.385 ;
      RECT 186.385 17.935 187.595 19.395 ;
      RECT 182.705 17.935 184.355 19.395 ;
      RECT 177.185 17.935 179.765 19.395 ;
      RECT 174.885 17.935 175.635 19.395 ;
      RECT 166.145 17.935 167.355 19.395 ;
      RECT 162.465 17.935 164.115 19.395 ;
      RECT 156.485 17.165 159.065 19.395 ;
      RECT 151.425 17.935 151.945 19.395 ;
      RECT 145.905 16.645 146.425 19.395 ;
      RECT 140.385 16.645 142.965 19.395 ;
      RECT 131.185 16.645 131.705 19.395 ;
      RECT 127.505 17.165 129.155 19.395 ;
      RECT 121.525 17.935 122.735 19.395 ;
      RECT 108.645 17.935 109.165 19.395 ;
      RECT 103.585 17.935 104.105 19.395 ;
      RECT 101.285 16.645 102.035 19.395 ;
      RECT 98.525 17.935 99.735 19.395 ;
      RECT 93.465 17.935 93.985 19.395 ;
      RECT 91.625 17.165 92.375 19.395 ;
      RECT 88.865 16.645 90.075 19.395 ;
      RECT 87.025 17.935 87.545 19.395 ;
      RECT 81.505 17.935 82.255 19.395 ;
      RECT 68.165 17.935 68.685 19.395 ;
      RECT 63.105 17.935 63.625 19.395 ;
      RECT 57.125 17.935 57.875 19.395 ;
      RECT 54.365 17.935 55.575 19.395 ;
      RECT 44.705 16.645 45.225 19.395 ;
      RECT 42.865 17.165 43.385 19.395 ;
      RECT 41.025 16.645 41.775 19.395 ;
      RECT 29.985 17.165 31.635 19.395 ;
      RECT 25.845 17.935 27.495 19.395 ;
      RECT 18.945 17.165 19.465 19.395 ;
      RECT 15.265 16.645 16.915 19.395 ;
      RECT 13.425 16.645 13.945 19.395 ;
      RECT 10.665 16.645 11.875 19.395 ;
      RECT 24.955 17.165 25.285 18.905 ;
      RECT 187.305 17.165 188.975 18.875 ;
      RECT 182.705 17.935 186.215 18.875 ;
      RECT 177.185 17.935 182.53 18.875 ;
      RECT 175.345 17.185 176.555 18.875 ;
      RECT 166.145 17.935 168.735 18.875 ;
      RECT 162.465 17.935 165.975 18.875 ;
      RECT 156.485 17.935 161.83 18.875 ;
      RECT 140.385 17.165 145.73 18.875 ;
      RECT 127.505 17.935 131.015 18.875 ;
      RECT 121.525 17.935 124.115 18.875 ;
      RECT 101.285 17.165 102.955 18.875 ;
      RECT 98.525 17.935 101.115 18.875 ;
      RECT 91.625 17.935 93.295 18.875 ;
      RECT 88.865 17.165 91.455 18.875 ;
      RECT 81.505 17.935 83.175 18.875 ;
      RECT 57.125 17.935 58.795 18.875 ;
      RECT 54.365 17.935 56.955 18.875 ;
      RECT 41.025 17.165 42.695 18.875 ;
      RECT 29.985 17.935 33.495 18.875 ;
      RECT 25.845 17.935 29.355 18.875 ;
      RECT 28.145 17.185 29.355 18.875 ;
      RECT 15.265 17.165 18.775 18.875 ;
      RECT 10.665 17.165 13.255 18.875 ;
      RECT 151.425 17.935 152.635 18.855 ;
      RECT 145.905 17.185 147.115 18.855 ;
      RECT 131.185 17.185 132.395 18.855 ;
      RECT 108.645 17.935 109.855 18.855 ;
      RECT 103.585 17.935 104.795 18.855 ;
      RECT 93.465 17.935 94.675 18.855 ;
      RECT 87.025 17.935 88.235 18.855 ;
      RECT 68.165 17.935 69.375 18.855 ;
      RECT 63.105 17.935 64.315 18.855 ;
      RECT 44.705 16.645 45.915 18.855 ;
      RECT 42.865 17.165 44.075 18.855 ;
      RECT 18.945 17.165 20.155 18.855 ;
      RECT 13.425 17.185 14.635 18.855 ;
      RECT 168.925 17.935 169.215 18.835 ;
      RECT 189.605 17.21 189.895 18.83 ;
      RECT 189.145 17.21 189.435 18.83 ;
      RECT 176.725 17.21 177.015 18.83 ;
      RECT 162.005 17.21 162.295 18.83 ;
      RECT 147.285 17.21 147.575 18.83 ;
      RECT 132.565 17.21 132.855 18.83 ;
      RECT 117.845 17.21 118.135 18.83 ;
      RECT 103.125 17.21 103.415 18.83 ;
      RECT 88.405 17.21 88.695 18.83 ;
      RECT 73.685 17.21 73.975 18.83 ;
      RECT 58.965 17.21 59.255 18.83 ;
      RECT 44.245 17.21 44.535 18.83 ;
      RECT 29.525 17.21 29.815 18.83 ;
      RECT 14.805 17.21 15.095 18.83 ;
      RECT 10.205 17.21 10.495 18.83 ;
      RECT 139.495 17.325 139.665 18.715 ;
      RECT 116.495 16.645 116.665 18.715 ;
      RECT 80.615 17.185 80.785 18.715 ;
      RECT 53.475 17.935 53.645 18.715 ;
      RECT 40.135 17.935 40.305 18.715 ;
      RECT 138.525 17.405 138.735 18.635 ;
      RECT 115.525 17.455 115.735 18.635 ;
      RECT 79.645 17.935 79.855 18.635 ;
      RECT 52.505 17.935 52.715 18.635 ;
      RECT 39.165 17.935 39.375 18.635 ;
      RECT 136.34 17.435 136.71 18.605 ;
      RECT 113.34 17.935 113.71 18.605 ;
      RECT 77.46 17.165 77.83 18.605 ;
      RECT 50.32 16.645 50.69 18.605 ;
      RECT 36.98 17.935 37.35 18.605 ;
      RECT 155.495 16.645 155.825 18.585 ;
      RECT 153.235 17.935 153.565 18.585 ;
      RECT 150.435 17.935 150.765 18.585 ;
      RECT 148.175 17.555 148.505 18.585 ;
      RECT 107.715 17.935 108.045 18.585 ;
      RECT 105.455 17.935 105.785 18.585 ;
      RECT 97.535 17.935 97.865 18.585 ;
      RECT 95.275 17.935 95.605 18.585 ;
      RECT 86.095 17.935 86.425 18.585 ;
      RECT 83.835 17.935 84.165 18.585 ;
      RECT 67.175 17.935 67.505 18.585 ;
      RECT 64.915 17.935 65.245 18.585 ;
      RECT 24.115 17.165 24.445 18.585 ;
      RECT 23.275 17.165 23.605 18.585 ;
      RECT 22.435 16.645 22.765 18.585 ;
      RECT 21.595 16.645 21.925 18.585 ;
      RECT 20.755 17.935 21.085 18.585 ;
      RECT 126.515 16.645 126.815 18.575 ;
      RECT 125.66 17.935 125.92 18.575 ;
      RECT 124.765 17.935 125.06 18.575 ;
      RECT 120.535 17.935 120.835 18.575 ;
      RECT 119.68 17.935 119.94 18.575 ;
      RECT 118.785 17.935 119.08 18.575 ;
      RECT 72.695 17.935 72.995 18.575 ;
      RECT 71.84 17.935 72.1 18.575 ;
      RECT 70.945 17.935 71.24 18.575 ;
      RECT 62.115 17.935 62.415 18.575 ;
      RECT 61.26 17.135 61.52 18.575 ;
      RECT 60.365 17.935 60.66 18.575 ;
      RECT 173.655 16.645 173.98 18.565 ;
      RECT 172.235 17.935 172.505 18.565 ;
      RECT 134.395 17.475 134.645 18.565 ;
      RECT 111.395 16.645 111.645 18.565 ;
      RECT 75.515 16.645 75.765 18.565 ;
      RECT 48.375 17.165 48.625 18.565 ;
      RECT 35.035 17.935 35.285 18.565 ;
      RECT 133.455 17.555 133.785 18.485 ;
      RECT 110.455 17.935 110.785 18.485 ;
      RECT 74.575 16.645 74.905 18.485 ;
      RECT 47.435 17.165 47.765 18.485 ;
      RECT 34.095 17.935 34.425 18.485 ;
      RECT 170.295 17.935 170.965 18.475 ;
      RECT 10.12 17.935 189.98 18.105 ;
      RECT 184.545 17.165 187.135 18.105 ;
      RECT 183.655 17.325 183.825 19.395 ;
      RECT 182.685 17.405 182.895 18.105 ;
      RECT 180.5 17.435 180.87 18.875 ;
      RECT 178.555 17.475 178.805 19.395 ;
      RECT 177.615 17.555 177.945 19.395 ;
      RECT 173.505 17.165 175.175 18.105 ;
      RECT 172.275 17.475 172.6 18.105 ;
      RECT 170.855 17.475 171.125 18.105 ;
      RECT 168.935 17.325 169.105 18.835 ;
      RECT 167.965 17.405 168.175 18.875 ;
      RECT 165.78 17.435 166.15 18.105 ;
      RECT 163.835 17.475 164.085 19.395 ;
      RECT 162.895 17.555 163.225 19.395 ;
      RECT 160.625 17.185 161.835 18.105 ;
      RECT 155.105 17.165 160.45 18.105 ;
      RECT 154.215 17.325 154.385 18.105 ;
      RECT 153.245 17.405 153.455 18.585 ;
      RECT 151.06 17.435 151.43 18.105 ;
      RECT 149.115 17.475 149.365 18.105 ;
      RECT 125.665 17.165 131.01 18.105 ;
      RECT 124.775 17.325 124.945 18.575 ;
      RECT 123.805 17.405 124.015 18.875 ;
      RECT 121.62 17.435 121.99 19.395 ;
      RECT 119.675 17.475 119.925 18.105 ;
      RECT 118.735 17.555 119.065 18.105 ;
      RECT 116.465 17.185 117.675 18.105 ;
      RECT 115.475 17.455 115.805 18.105 ;
      RECT 113.215 17.455 113.545 18.105 ;
      RECT 110.945 17.165 112.615 18.105 ;
      RECT 110.055 17.325 110.225 18.105 ;
      RECT 109.085 17.405 109.295 18.855 ;
      RECT 106.9 17.435 107.27 18.105 ;
      RECT 104.955 17.475 105.205 18.105 ;
      RECT 104.015 17.555 104.345 18.855 ;
      RECT 100.395 17.325 100.565 18.875 ;
      RECT 99.425 17.405 99.635 19.395 ;
      RECT 97.24 17.435 97.61 18.105 ;
      RECT 95.295 17.475 95.545 18.585 ;
      RECT 94.355 17.555 94.685 18.105 ;
      RECT 92.545 17.185 93.755 18.105 ;
      RECT 88.865 17.165 92.375 18.105 ;
      RECT 87.515 17.325 87.685 18.855 ;
      RECT 86.545 17.405 86.755 18.105 ;
      RECT 84.36 17.435 84.73 18.105 ;
      RECT 82.415 17.475 82.665 18.875 ;
      RECT 81.475 17.555 81.805 18.105 ;
      RECT 79.665 17.185 80.875 18.105 ;
      RECT 74.145 17.165 79.49 18.105 ;
      RECT 72.795 17.325 72.965 18.575 ;
      RECT 71.825 17.405 72.035 18.105 ;
      RECT 69.64 17.435 70.01 18.105 ;
      RECT 67.695 17.475 67.945 18.105 ;
      RECT 66.755 17.555 67.085 18.105 ;
      RECT 65.395 17.455 65.725 18.105 ;
      RECT 64.555 17.455 64.885 18.105 ;
      RECT 63.715 17.455 64.045 18.855 ;
      RECT 62.875 17.455 63.205 18.105 ;
      RECT 62.035 17.455 62.365 18.105 ;
      RECT 61.195 17.135 61.525 18.105 ;
      RECT 59.425 17.185 60.635 18.105 ;
      RECT 58.075 17.325 58.245 18.875 ;
      RECT 57.105 17.405 57.315 18.105 ;
      RECT 54.92 17.435 55.29 19.395 ;
      RECT 52.975 17.475 53.225 18.105 ;
      RECT 52.035 17.555 52.365 18.105 ;
      RECT 50.225 17.185 51.435 18.105 ;
      RECT 44.705 17.165 50.05 18.105 ;
      RECT 40.565 17.165 44.075 18.105 ;
      RECT 39.675 17.325 39.845 18.105 ;
      RECT 38.705 17.405 38.915 18.105 ;
      RECT 36.52 17.435 36.89 18.105 ;
      RECT 34.575 17.475 34.825 18.105 ;
      RECT 33.635 17.555 33.965 18.105 ;
      RECT 31.825 17.185 33.035 18.875 ;
      RECT 29.985 17.165 31.655 18.875 ;
      RECT 26.305 17.165 27.975 18.875 ;
      RECT 20.785 17.165 26.13 18.105 ;
      RECT 15.265 17.165 20.61 18.105 ;
      RECT 175.345 16.645 175.865 18.875 ;
      RECT 160.625 16.645 161.145 18.875 ;
      RECT 116.465 16.645 116.985 18.105 ;
      RECT 92.545 16.645 93.065 18.875 ;
      RECT 79.665 16.645 80.185 18.105 ;
      RECT 59.425 16.645 59.945 18.105 ;
      RECT 50.225 16.645 50.745 18.105 ;
      RECT 31.825 16.645 32.345 18.875 ;
      RECT 28.145 16.645 28.665 18.875 ;
      RECT 187.305 16.645 188.055 18.875 ;
      RECT 184.545 16.645 185.755 18.875 ;
      RECT 173.505 16.645 174.255 18.105 ;
      RECT 155.105 16.645 157.685 18.105 ;
      RECT 125.665 16.645 128.245 18.105 ;
      RECT 110.945 16.645 111.695 18.105 ;
      RECT 88.865 16.645 90.515 18.875 ;
      RECT 74.145 16.645 76.725 18.105 ;
      RECT 44.705 16.645 47.285 18.105 ;
      RECT 40.565 16.645 42.215 18.105 ;
      RECT 29.985 16.645 30.735 19.395 ;
      RECT 26.305 16.645 27.055 19.395 ;
      RECT 20.785 16.645 23.365 18.105 ;
      RECT 15.265 16.645 17.845 18.875 ;
      RECT 170.515 20.655 171.035 22.455 ;
      RECT 146.595 19.025 147.115 22.455 ;
      RECT 107.955 20.655 108.475 22.455 ;
      RECT 101.515 19.565 102.035 22.455 ;
      RECT 72.995 20.655 73.515 22.455 ;
      RECT 73.13 19.82 73.515 22.455 ;
      RECT 58.275 19.045 58.795 22.455 ;
      RECT 15.955 19.565 16.475 22.455 ;
      RECT 14.115 19.025 14.635 22.455 ;
      RECT 187.765 19.045 188.975 22.435 ;
      RECT 184.525 19.045 186.215 22.435 ;
      RECT 179.935 19.045 182.53 22.435 ;
      RECT 168.905 20.655 169.655 22.435 ;
      RECT 165.215 20.655 167.81 22.435 ;
      RECT 160.625 20.655 161.835 22.435 ;
      RECT 157.385 19.565 159.075 22.435 ;
      RECT 140.365 20.655 142.055 22.435 ;
      RECT 133.945 20.655 134.695 22.435 ;
      RECT 119.685 20.655 120.895 22.435 ;
      RECT 113.245 20.655 113.995 22.435 ;
      RECT 105.405 20.655 107.095 22.435 ;
      RECT 92.545 19.045 93.295 22.435 ;
      RECT 90.245 19.045 91.455 22.435 ;
      RECT 81.045 20.655 82.255 22.435 ;
      RECT 76.895 20.655 79.49 22.435 ;
      RECT 70.445 20.655 72.135 22.435 ;
      RECT 62.175 20.655 64.77 22.435 ;
      RECT 56.665 20.655 57.415 22.435 ;
      RECT 52.975 20.655 55.57 22.435 ;
      RECT 47.455 20.655 50.05 22.435 ;
      RECT 36.885 20.655 38.095 22.435 ;
      RECT 28.145 19.045 29.355 22.435 ;
      RECT 24.905 20.655 26.595 22.435 ;
      RECT 12.045 19.045 13.255 22.435 ;
      RECT 189.605 19.49 189.895 21.99 ;
      RECT 189.145 19.49 189.435 21.99 ;
      RECT 176.725 19.49 177.015 21.99 ;
      RECT 162.005 19.49 162.295 21.99 ;
      RECT 147.285 19.49 147.575 21.99 ;
      RECT 132.565 19.49 132.855 21.99 ;
      RECT 117.845 19.49 118.135 21.99 ;
      RECT 103.125 19.49 103.415 21.99 ;
      RECT 88.405 19.49 88.695 21.99 ;
      RECT 73.685 19.49 73.975 21.99 ;
      RECT 58.965 19.49 59.255 21.99 ;
      RECT 44.245 19.49 44.535 21.99 ;
      RECT 29.525 19.49 29.815 21.99 ;
      RECT 14.805 19.49 15.095 21.99 ;
      RECT 10.205 19.49 10.495 21.99 ;
      RECT 175.835 19.045 176.165 21.975 ;
      RECT 150.435 20.655 150.765 21.975 ;
      RECT 145.47 19.045 145.73 21.975 ;
      RECT 143.63 19.045 143.89 21.975 ;
      RECT 82.815 19.045 83.145 21.975 ;
      RECT 38.655 20.655 38.985 21.975 ;
      RECT 30.375 19.565 30.705 21.975 ;
      RECT 22.195 20.655 22.525 21.975 ;
      RECT 149.145 20.655 149.355 21.965 ;
      RECT 148.245 20.655 148.475 21.965 ;
      RECT 186.385 19.565 188.975 21.915 ;
      RECT 182.705 19.565 186.215 21.915 ;
      RECT 177.185 19.565 182.53 21.915 ;
      RECT 169.825 20.655 171.035 21.915 ;
      RECT 167.985 20.655 169.655 21.915 ;
      RECT 164.285 19.045 165.975 21.915 ;
      RECT 159.245 20.655 161.835 21.915 ;
      RECT 155.565 20.655 159.075 21.915 ;
      RECT 145.905 19.565 147.115 21.915 ;
      RECT 138.545 20.655 142.055 21.915 ;
      RECT 133.025 20.655 134.695 21.915 ;
      RECT 118.305 20.655 120.895 21.915 ;
      RECT 112.325 20.655 113.995 21.915 ;
      RECT 107.265 20.655 108.475 21.915 ;
      RECT 103.585 20.655 107.095 21.915 ;
      RECT 100.825 20.655 102.035 21.915 ;
      RECT 91.625 19.565 93.295 21.915 ;
      RECT 88.865 19.565 91.455 21.915 ;
      RECT 79.665 20.655 82.255 21.915 ;
      RECT 74.145 20.655 79.49 21.915 ;
      RECT 72.305 20.655 73.515 21.915 ;
      RECT 68.625 20.655 72.135 21.915 ;
      RECT 59.425 20.655 64.77 21.915 ;
      RECT 57.585 19.565 58.795 21.915 ;
      RECT 58.045 19.045 58.795 21.915 ;
      RECT 55.745 19.045 56.955 21.915 ;
      RECT 50.225 20.655 55.57 21.915 ;
      RECT 44.705 20.655 50.05 21.915 ;
      RECT 47.435 20.155 47.765 21.915 ;
      RECT 35.505 20.655 38.095 21.915 ;
      RECT 26.765 19.565 29.355 21.915 ;
      RECT 27.665 19.045 29.355 21.915 ;
      RECT 23.085 20.655 26.595 21.915 ;
      RECT 15.265 19.565 16.475 21.915 ;
      RECT 13.425 19.565 14.635 21.915 ;
      RECT 10.665 19.565 13.255 21.915 ;
      RECT 127.525 19.565 127.695 21.835 ;
      RECT 99.925 19.045 100.095 21.835 ;
      RECT 174.995 19.565 175.325 21.625 ;
      RECT 174.155 20.655 174.485 21.625 ;
      RECT 173.315 20.655 173.645 21.625 ;
      RECT 172.555 20.655 172.725 21.625 ;
      RECT 171.715 20.655 171.885 21.625 ;
      RECT 154.715 20.235 154.885 21.625 ;
      RECT 153.875 20.655 154.045 21.625 ;
      RECT 152.955 20.655 153.285 21.625 ;
      RECT 152.115 19.025 152.445 21.625 ;
      RECT 151.275 20.655 151.605 21.625 ;
      RECT 124.59 20.655 124.76 21.625 ;
      RECT 96.99 20.655 97.16 21.625 ;
      RECT 87.095 19.565 87.265 21.625 ;
      RECT 86.255 20.655 86.425 21.625 ;
      RECT 85.335 20.655 85.665 21.625 ;
      RECT 84.495 20.655 84.825 21.625 ;
      RECT 83.655 20.655 83.985 21.625 ;
      RECT 42.935 19.565 43.105 21.625 ;
      RECT 42.095 19.045 42.265 21.625 ;
      RECT 41.175 19.565 41.505 21.625 ;
      RECT 40.335 20.655 40.665 21.625 ;
      RECT 39.495 20.655 39.825 21.625 ;
      RECT 34.655 20.655 34.825 21.625 ;
      RECT 33.815 20.655 33.985 21.625 ;
      RECT 32.895 19.045 33.225 21.625 ;
      RECT 32.055 19.045 32.385 21.625 ;
      RECT 31.215 19.565 31.545 21.625 ;
      RECT 21.355 20.655 21.685 21.625 ;
      RECT 20.515 20.655 20.845 21.625 ;
      RECT 19.675 19.025 20.005 21.625 ;
      RECT 18.915 20.655 19.085 21.625 ;
      RECT 18.075 19.045 18.245 21.625 ;
      RECT 144.54 19.045 144.87 21.585 ;
      RECT 142.7 19.565 143.03 21.585 ;
      RECT 135.31 20.655 135.64 21.585 ;
      RECT 131.16 20.655 131.49 21.585 ;
      RECT 116.9 20.655 117.23 21.585 ;
      RECT 109.09 19.565 109.42 21.585 ;
      RECT 67.68 20.655 68.01 21.585 ;
      RECT 126.47 20.655 126.785 21.325 ;
      RECT 121.495 20.655 121.825 21.325 ;
      RECT 98.87 19.565 99.185 21.325 ;
      RECT 93.895 19.565 94.225 21.325 ;
      RECT 122.42 19.565 122.685 21.285 ;
      RECT 94.82 20.655 95.085 21.285 ;
      RECT 136.23 20.655 136.585 21.245 ;
      RECT 130.215 19.045 130.57 21.245 ;
      RECT 115.955 20.655 116.31 21.245 ;
      RECT 110.01 20.655 110.365 21.245 ;
      RECT 66.735 20.655 67.09 21.245 ;
      RECT 10.12 20.655 189.98 20.825 ;
      RECT 174.885 19.565 176.555 20.825 ;
      RECT 175.805 19.045 176.555 20.825 ;
      RECT 173.655 20.195 173.98 20.825 ;
      RECT 172.235 20.195 172.505 20.825 ;
      RECT 170.715 19.925 171.055 20.825 ;
      RECT 169.355 19.945 169.685 20.825 ;
      RECT 166.145 19.565 168.735 20.825 ;
      RECT 162.465 19.565 165.975 21.915 ;
      RECT 156.485 19.565 161.83 20.825 ;
      RECT 159.235 19.045 161.83 20.825 ;
      RECT 155.54 19.895 155.87 20.825 ;
      RECT 154.595 20.235 154.95 20.825 ;
      RECT 151.425 19.565 152.635 20.825 ;
      RECT 152.115 19.025 152.635 20.825 ;
      RECT 150.48 19.895 150.81 20.825 ;
      RECT 149.535 20.235 149.89 20.825 ;
      RECT 140.385 19.565 145.73 20.825 ;
      RECT 143.135 19.045 145.73 20.825 ;
      RECT 139.485 19.645 139.655 21.915 ;
      RECT 138.43 20.155 138.745 20.825 ;
      RECT 136.55 19.855 136.72 20.825 ;
      RECT 134.38 20.195 134.645 22.435 ;
      RECT 133.455 20.155 133.785 21.915 ;
      RECT 131.185 19.565 132.395 20.825 ;
      RECT 131.875 19.025 132.395 20.825 ;
      RECT 127.505 19.565 131.015 20.825 ;
      RECT 129.325 19.045 131.015 20.825 ;
      RECT 126.95 19.82 127.335 20.825 ;
      RECT 126.09 19.82 126.35 20.825 ;
      RECT 125.23 19.82 125.49 20.825 ;
      RECT 124.285 19.82 124.63 20.825 ;
      RECT 121.525 19.565 124.115 20.825 ;
      RECT 122.905 19.045 124.115 20.825 ;
      RECT 120.97 19.82 121.355 20.825 ;
      RECT 120.11 19.82 120.37 22.435 ;
      RECT 119.25 19.82 119.51 21.915 ;
      RECT 118.305 19.82 118.65 21.915 ;
      RECT 116.485 19.645 116.655 20.825 ;
      RECT 115.43 20.155 115.745 20.825 ;
      RECT 113.55 19.855 113.72 22.435 ;
      RECT 111.38 20.195 111.645 20.825 ;
      RECT 110.455 20.155 110.785 20.825 ;
      RECT 108.645 19.565 109.855 20.825 ;
      RECT 109.335 19.025 109.855 20.825 ;
      RECT 106.33 20.235 106.685 22.435 ;
      RECT 105.41 19.895 105.74 22.435 ;
      RECT 103.585 19.565 104.795 21.915 ;
      RECT 104.275 19.025 104.795 21.915 ;
      RECT 101.285 19.565 102.955 20.825 ;
      RECT 102.205 19.045 102.955 20.825 ;
      RECT 98.525 19.565 101.115 20.825 ;
      RECT 97.58 19.895 97.91 20.825 ;
      RECT 96.635 20.235 96.99 20.825 ;
      RECT 93.465 19.565 94.675 20.825 ;
      RECT 94.155 19.025 94.675 20.825 ;
      RECT 87.025 19.565 88.235 20.825 ;
      RECT 87.715 19.025 88.235 20.825 ;
      RECT 84.71 20.235 85.065 20.825 ;
      RECT 83.79 19.895 84.12 20.825 ;
      RECT 81.505 19.565 83.175 20.825 ;
      RECT 82.425 19.045 83.175 20.825 ;
      RECT 80.605 19.645 80.775 21.915 ;
      RECT 79.55 20.155 79.865 20.825 ;
      RECT 77.67 19.855 77.84 22.435 ;
      RECT 75.5 20.195 75.765 21.915 ;
      RECT 74.575 20.155 74.905 21.915 ;
      RECT 72.27 19.82 72.53 20.825 ;
      RECT 71.41 19.82 71.67 22.435 ;
      RECT 70.465 19.82 70.81 22.435 ;
      RECT 68.165 19.565 69.375 20.825 ;
      RECT 68.855 19.025 69.375 21.915 ;
      RECT 67.22 19.895 67.55 20.825 ;
      RECT 66.275 20.235 66.63 20.825 ;
      RECT 63.105 19.565 64.315 22.435 ;
      RECT 63.795 19.025 64.315 22.435 ;
      RECT 62.55 19.82 62.935 22.435 ;
      RECT 61.69 19.82 61.95 21.915 ;
      RECT 60.83 19.82 61.09 21.915 ;
      RECT 59.885 19.82 60.23 21.915 ;
      RECT 57.125 19.565 58.795 20.825 ;
      RECT 54.365 19.565 56.955 20.825 ;
      RECT 53.465 19.645 53.635 22.435 ;
      RECT 52.41 20.155 52.725 21.915 ;
      RECT 50.53 19.855 50.7 21.915 ;
      RECT 48.36 20.195 48.625 22.435 ;
      RECT 44.705 19.565 45.915 21.915 ;
      RECT 45.395 19.025 45.915 21.915 ;
      RECT 42.865 19.565 44.075 20.825 ;
      RECT 43.555 19.025 44.075 20.825 ;
      RECT 41.025 19.565 42.695 20.825 ;
      RECT 41.945 19.045 42.695 20.825 ;
      RECT 40.125 19.645 40.295 20.825 ;
      RECT 39.07 20.155 39.385 20.825 ;
      RECT 37.19 19.855 37.36 22.435 ;
      RECT 35.02 20.195 35.285 20.825 ;
      RECT 34.095 20.155 34.425 20.825 ;
      RECT 29.985 19.565 33.495 20.825 ;
      RECT 31.805 19.045 33.495 20.825 ;
      RECT 25.845 19.565 29.355 20.825 ;
      RECT 24.955 19.505 25.285 22.435 ;
      RECT 24.115 19.855 24.445 21.915 ;
      RECT 23.275 19.855 23.605 21.915 ;
      RECT 22.435 19.855 22.765 20.825 ;
      RECT 21.675 19.855 21.845 20.825 ;
      RECT 20.835 19.855 21.005 20.825 ;
      RECT 18.945 19.565 20.155 20.825 ;
      RECT 19.635 19.025 20.155 20.825 ;
      RECT 15.265 19.565 18.775 20.825 ;
      RECT 17.085 19.045 18.775 20.825 ;
      RECT 167.525 19.045 168.735 20.825 ;
      RECT 99.905 19.045 101.115 20.825 ;
      RECT 186.385 22.085 187.595 24.835 ;
      RECT 182.705 22.085 184.355 24.835 ;
      RECT 177.185 22.085 179.765 24.835 ;
      RECT 175.345 23.375 175.865 24.835 ;
      RECT 173.505 23.375 174.255 24.835 ;
      RECT 167.985 23.375 170.565 24.835 ;
      RECT 162.465 22.085 165.045 24.835 ;
      RECT 160.625 22.605 161.145 24.835 ;
      RECT 158.785 23.375 159.535 24.835 ;
      RECT 153.265 23.375 155.845 24.835 ;
      RECT 147.745 23.375 150.325 24.835 ;
      RECT 144.525 23.375 145.735 24.835 ;
      RECT 138.085 23.375 139.295 24.835 ;
      RECT 133.025 22.085 133.545 24.835 ;
      RECT 131.185 23.375 131.705 24.835 ;
      RECT 129.345 23.375 130.095 24.835 ;
      RECT 123.825 23.375 126.405 24.835 ;
      RECT 118.305 22.605 120.885 24.835 ;
      RECT 110.945 23.375 111.465 24.835 ;
      RECT 109.105 23.375 109.855 24.835 ;
      RECT 103.585 22.605 106.165 24.835 ;
      RECT 101.285 22.625 102.035 24.835 ;
      RECT 98.525 23.375 99.735 24.835 ;
      RECT 93.465 23.375 93.985 24.835 ;
      RECT 91.625 22.085 92.375 24.835 ;
      RECT 88.865 22.085 90.075 24.835 ;
      RECT 85.645 23.375 86.855 24.835 ;
      RECT 79.205 23.375 80.415 24.835 ;
      RECT 74.145 22.085 74.665 24.835 ;
      RECT 70.925 22.605 72.135 24.835 ;
      RECT 65.865 23.375 66.385 24.835 ;
      RECT 63.105 22.605 64.315 24.835 ;
      RECT 59.425 22.085 61.075 24.835 ;
      RECT 56.205 22.605 57.415 24.835 ;
      RECT 50.685 22.605 53.265 24.835 ;
      RECT 38.725 23.375 41.305 24.835 ;
      RECT 33.665 23.375 34.185 24.835 ;
      RECT 29.985 23.375 31.635 24.835 ;
      RECT 28.145 22.605 28.665 24.835 ;
      RECT 26.305 23.375 27.055 24.835 ;
      RECT 20.785 23.375 23.365 24.835 ;
      RECT 15.265 23.375 17.845 24.835 ;
      RECT 13.425 22.085 13.945 24.835 ;
      RECT 10.665 22.085 11.875 24.835 ;
      RECT 116.955 23.375 117.285 24.345 ;
      RECT 45.555 22.085 45.885 24.345 ;
      RECT 186.385 22.605 188.975 24.315 ;
      RECT 182.705 22.605 186.215 24.315 ;
      RECT 177.185 22.605 182.53 24.315 ;
      RECT 173.505 23.375 175.175 24.315 ;
      RECT 167.985 23.375 173.33 24.315 ;
      RECT 162.465 22.605 167.81 24.315 ;
      RECT 159.245 22.085 160.455 24.315 ;
      RECT 153.265 23.375 158.61 24.315 ;
      RECT 147.745 23.375 153.09 24.315 ;
      RECT 144.525 23.375 147.115 24.315 ;
      RECT 145.905 22.625 147.115 24.315 ;
      RECT 138.085 23.375 140.675 24.315 ;
      RECT 129.345 23.375 131.015 24.315 ;
      RECT 123.825 23.375 129.17 24.315 ;
      RECT 118.305 23.375 123.65 24.315 ;
      RECT 109.105 23.375 110.775 24.315 ;
      RECT 103.585 23.375 108.93 24.315 ;
      RECT 101.285 23.375 102.955 24.315 ;
      RECT 98.525 23.375 101.115 24.315 ;
      RECT 91.625 22.605 93.295 24.315 ;
      RECT 88.865 22.605 91.455 24.315 ;
      RECT 85.645 23.375 88.235 24.315 ;
      RECT 79.205 23.375 81.795 24.315 ;
      RECT 70.925 23.375 73.515 24.315 ;
      RECT 72.305 22.625 73.515 24.315 ;
      RECT 63.105 23.375 65.695 24.315 ;
      RECT 59.425 22.605 62.935 24.315 ;
      RECT 56.205 23.375 58.795 24.315 ;
      RECT 57.585 22.625 58.795 24.315 ;
      RECT 50.685 23.375 56.03 24.315 ;
      RECT 38.725 23.375 44.07 24.315 ;
      RECT 29.985 23.375 33.495 24.315 ;
      RECT 26.765 22.085 27.975 24.315 ;
      RECT 20.785 23.375 26.13 24.315 ;
      RECT 15.265 23.375 20.61 24.315 ;
      RECT 10.665 22.605 13.255 24.315 ;
      RECT 175.345 23.375 176.555 24.295 ;
      RECT 160.625 22.605 161.835 24.295 ;
      RECT 133.025 22.605 134.235 24.295 ;
      RECT 131.185 23.375 132.395 24.295 ;
      RECT 110.945 23.375 112.155 24.295 ;
      RECT 93.465 23.375 94.675 24.295 ;
      RECT 74.145 22.085 75.355 24.295 ;
      RECT 65.865 23.375 67.075 24.295 ;
      RECT 33.665 23.375 34.875 24.295 ;
      RECT 28.145 22.605 29.355 24.295 ;
      RECT 13.425 22.625 14.635 24.295 ;
      RECT 189.605 22.65 189.895 24.27 ;
      RECT 189.145 22.65 189.435 24.27 ;
      RECT 176.725 22.65 177.015 24.27 ;
      RECT 162.005 22.65 162.295 24.27 ;
      RECT 147.285 22.65 147.575 24.27 ;
      RECT 132.565 22.65 132.855 24.27 ;
      RECT 117.845 22.65 118.135 24.27 ;
      RECT 103.125 22.65 103.415 24.27 ;
      RECT 88.405 22.65 88.695 24.27 ;
      RECT 73.685 22.65 73.975 24.27 ;
      RECT 58.965 22.65 59.255 24.27 ;
      RECT 44.245 22.65 44.535 24.27 ;
      RECT 29.525 22.65 29.815 24.27 ;
      RECT 14.805 22.65 15.095 24.27 ;
      RECT 10.205 22.65 10.495 24.27 ;
      RECT 143.595 23.375 143.925 24.025 ;
      RECT 141.335 22.605 141.665 24.025 ;
      RECT 137.155 23.375 137.485 24.025 ;
      RECT 134.895 23.375 135.225 24.025 ;
      RECT 116.115 23.375 116.445 24.025 ;
      RECT 115.275 23.375 115.605 24.025 ;
      RECT 114.435 23.375 114.765 24.025 ;
      RECT 113.595 22.605 113.925 24.025 ;
      RECT 112.755 22.605 113.085 24.025 ;
      RECT 97.535 23.375 97.865 24.025 ;
      RECT 95.275 23.375 95.605 24.025 ;
      RECT 84.715 23.375 85.045 24.025 ;
      RECT 82.455 23.375 82.785 24.025 ;
      RECT 78.275 22.605 78.605 24.025 ;
      RECT 76.015 22.085 76.345 24.025 ;
      RECT 69.995 22.605 70.325 24.025 ;
      RECT 67.735 23.375 68.065 24.025 ;
      RECT 49.755 23.375 50.085 24.025 ;
      RECT 48.915 22.605 49.245 24.025 ;
      RECT 48.075 22.605 48.405 24.025 ;
      RECT 47.235 22.605 47.565 24.025 ;
      RECT 46.395 22.085 46.725 24.025 ;
      RECT 37.735 22.605 38.065 24.025 ;
      RECT 35.475 23.375 35.805 24.025 ;
      RECT 10.12 23.375 189.98 23.545 ;
      RECT 175.835 22.575 176.165 24.295 ;
      RECT 174.995 22.895 175.325 23.545 ;
      RECT 174.155 22.895 174.485 24.315 ;
      RECT 173.315 22.895 173.645 23.545 ;
      RECT 172.475 22.895 172.805 24.315 ;
      RECT 171.635 22.895 171.965 24.315 ;
      RECT 169.825 22.625 171.035 24.315 ;
      RECT 167.985 22.605 169.655 24.835 ;
      RECT 159.245 22.605 161.835 23.545 ;
      RECT 155.565 22.605 159.075 23.545 ;
      RECT 154.635 22.895 154.965 24.835 ;
      RECT 153.795 22.895 154.125 24.835 ;
      RECT 152.955 22.895 153.285 23.545 ;
      RECT 152.115 22.895 152.445 24.315 ;
      RECT 151.275 22.895 151.605 24.315 ;
      RECT 150.435 22.575 150.765 24.315 ;
      RECT 149.145 22.555 149.355 24.835 ;
      RECT 148.245 22.555 148.475 24.835 ;
      RECT 145.47 22.535 145.73 24.835 ;
      RECT 144.54 22.995 144.87 24.835 ;
      RECT 143.63 22.535 143.89 24.025 ;
      RECT 142.7 22.995 143.03 23.545 ;
      RECT 138.545 22.605 142.055 23.545 ;
      RECT 137.615 22.895 137.945 23.545 ;
      RECT 135.355 22.895 135.685 23.545 ;
      RECT 133.025 22.605 134.695 23.545 ;
      RECT 131.115 22.895 131.445 23.545 ;
      RECT 128.855 22.895 129.185 23.545 ;
      RECT 127.535 22.765 127.705 24.315 ;
      RECT 126.565 22.845 126.775 24.315 ;
      RECT 124.38 22.875 124.75 24.835 ;
      RECT 122.435 22.915 122.685 24.315 ;
      RECT 121.495 22.995 121.825 24.315 ;
      RECT 118.305 22.605 120.895 24.315 ;
      RECT 116.855 22.895 117.185 23.545 ;
      RECT 114.595 22.895 114.925 23.545 ;
      RECT 112.325 22.605 113.995 23.545 ;
      RECT 111.395 22.895 111.725 24.295 ;
      RECT 109.135 22.895 109.465 24.835 ;
      RECT 107.265 22.625 108.475 24.315 ;
      RECT 103.585 22.605 107.095 24.315 ;
      RECT 100.825 22.085 101.345 23.545 ;
      RECT 99.935 22.765 100.105 24.315 ;
      RECT 98.965 22.845 99.175 24.835 ;
      RECT 96.78 22.875 97.15 23.545 ;
      RECT 94.835 22.915 95.085 23.545 ;
      RECT 93.895 22.995 94.225 24.295 ;
      RECT 87.015 22.895 87.345 24.315 ;
      RECT 86.175 22.895 86.505 24.835 ;
      RECT 85.335 22.895 85.665 23.545 ;
      RECT 84.495 22.895 84.825 23.545 ;
      RECT 83.655 22.895 83.985 23.545 ;
      RECT 82.815 22.575 83.145 23.545 ;
      RECT 79.665 22.605 82.255 23.545 ;
      RECT 74.145 22.605 79.49 23.545 ;
      RECT 68.625 22.605 72.135 23.545 ;
      RECT 67.635 22.895 67.965 23.545 ;
      RECT 65.375 22.895 65.705 23.545 ;
      RECT 59.425 22.605 64.77 23.545 ;
      RECT 55.745 22.085 56.495 23.545 ;
      RECT 50.225 22.605 55.57 23.545 ;
      RECT 44.705 22.605 50.05 23.545 ;
      RECT 42.855 22.895 43.185 24.315 ;
      RECT 42.015 22.895 42.345 24.315 ;
      RECT 41.175 22.895 41.505 24.315 ;
      RECT 40.335 22.895 40.665 24.835 ;
      RECT 39.495 22.895 39.825 24.835 ;
      RECT 38.655 22.575 38.985 23.545 ;
      RECT 35.505 22.605 38.095 23.545 ;
      RECT 34.575 22.895 34.905 23.545 ;
      RECT 33.735 22.895 34.065 24.835 ;
      RECT 32.895 22.895 33.225 24.315 ;
      RECT 32.055 22.895 32.385 24.315 ;
      RECT 31.215 22.895 31.545 24.835 ;
      RECT 30.375 22.575 30.705 24.835 ;
      RECT 26.765 22.605 29.355 23.545 ;
      RECT 23.085 22.605 26.595 23.545 ;
      RECT 22.195 22.575 22.525 24.835 ;
      RECT 21.355 22.895 21.685 24.835 ;
      RECT 20.515 22.895 20.845 23.545 ;
      RECT 19.675 22.895 20.005 24.315 ;
      RECT 18.835 22.895 19.165 24.315 ;
      RECT 17.995 22.895 18.325 24.315 ;
      RECT 15.265 22.625 16.475 24.835 ;
      RECT 169.825 22.085 170.345 24.835 ;
      RECT 145.905 22.085 146.425 24.315 ;
      RECT 107.265 22.085 107.785 24.315 ;
      RECT 72.305 22.085 72.825 24.315 ;
      RECT 57.585 22.085 58.105 24.315 ;
      RECT 15.265 22.085 15.785 24.835 ;
      RECT 167.985 22.085 168.735 24.835 ;
      RECT 155.565 22.085 157.215 24.315 ;
      RECT 138.545 22.085 140.195 24.315 ;
      RECT 133.025 22.085 133.775 24.295 ;
      RECT 118.305 22.085 119.515 24.835 ;
      RECT 112.325 22.085 113.075 23.545 ;
      RECT 103.585 22.085 105.235 24.835 ;
      RECT 79.665 22.085 80.875 24.315 ;
      RECT 74.145 22.085 76.725 23.545 ;
      RECT 68.625 22.085 70.275 23.545 ;
      RECT 59.425 22.085 62.005 24.315 ;
      RECT 50.225 22.085 52.805 23.545 ;
      RECT 44.705 22.085 47.285 23.545 ;
      RECT 35.505 22.085 36.715 23.545 ;
      RECT 23.085 22.085 24.735 24.315 ;
      RECT 176.035 24.465 176.555 27.895 ;
      RECT 152.115 24.485 152.635 27.895 ;
      RECT 146.595 24.485 147.115 27.895 ;
      RECT 126.355 25.005 126.875 27.895 ;
      RECT 109.795 25.005 110.315 27.895 ;
      RECT 102.435 24.485 102.955 27.895 ;
      RECT 87.715 24.485 88.235 27.895 ;
      RECT 72.075 25.005 72.595 27.895 ;
      RECT 50.915 25.005 51.435 27.895 ;
      RECT 36.195 26.095 36.715 27.895 ;
      RECT 21.475 25.005 21.995 27.895 ;
      RECT 14.115 24.465 14.635 27.895 ;
      RECT 187.765 24.485 188.975 27.875 ;
      RECT 184.525 24.485 186.215 27.875 ;
      RECT 179.935 24.485 182.53 27.875 ;
      RECT 174.425 24.485 175.175 27.875 ;
      RECT 170.735 24.485 173.33 27.875 ;
      RECT 165.215 24.485 167.81 27.875 ;
      RECT 159.235 26.095 161.83 27.875 ;
      RECT 149.565 25.005 151.255 27.875 ;
      RECT 135.775 26.095 138.37 27.875 ;
      RECT 131.645 25.005 132.395 27.875 ;
      RECT 131.875 24.465 132.395 27.875 ;
      RECT 124.745 25.005 125.495 27.875 ;
      RECT 121.055 24.485 123.65 27.875 ;
      RECT 106.335 24.485 108.93 27.875 ;
      RECT 100.825 26.095 101.575 27.875 ;
      RECT 97.135 26.095 99.73 27.875 ;
      RECT 91.615 26.095 94.21 27.875 ;
      RECT 86.105 25.005 86.855 27.875 ;
      RECT 75.965 26.095 77.655 27.875 ;
      RECT 63.105 25.005 63.855 27.875 ;
      RECT 60.805 25.005 62.015 27.875 ;
      RECT 47.455 26.095 50.05 27.875 ;
      RECT 32.735 26.095 35.33 27.875 ;
      RECT 18.015 24.485 20.61 27.875 ;
      RECT 12.045 24.485 13.255 27.875 ;
      RECT 189.605 24.93 189.895 27.43 ;
      RECT 189.145 24.93 189.435 27.43 ;
      RECT 176.725 24.93 177.015 27.43 ;
      RECT 162.005 24.93 162.295 27.43 ;
      RECT 147.285 24.93 147.575 27.43 ;
      RECT 132.565 24.93 132.855 27.43 ;
      RECT 117.845 24.93 118.135 27.43 ;
      RECT 103.125 24.93 103.415 27.43 ;
      RECT 88.405 24.93 88.695 27.43 ;
      RECT 73.685 24.93 73.975 27.43 ;
      RECT 58.965 24.93 59.255 27.43 ;
      RECT 44.245 24.93 44.535 27.43 ;
      RECT 29.525 24.93 29.815 27.43 ;
      RECT 14.805 24.93 15.095 27.43 ;
      RECT 10.205 24.93 10.495 27.43 ;
      RECT 186.385 25.005 188.975 27.355 ;
      RECT 182.705 25.005 186.215 27.355 ;
      RECT 177.185 25.005 182.53 27.355 ;
      RECT 175.345 25.005 176.555 27.355 ;
      RECT 173.505 25.005 175.175 27.355 ;
      RECT 167.985 25.005 173.33 27.355 ;
      RECT 162.465 25.005 167.81 27.355 ;
      RECT 156.485 26.095 161.83 27.355 ;
      RECT 158.785 25.005 160.455 27.355 ;
      RECT 151.425 24.485 152.635 27.355 ;
      RECT 147.745 25.005 151.255 27.355 ;
      RECT 145.905 24.485 147.115 27.355 ;
      RECT 133.025 26.095 138.37 27.355 ;
      RECT 135.77 25.675 136.125 27.355 ;
      RECT 130.725 26.095 132.395 27.355 ;
      RECT 131.185 25.005 132.395 27.355 ;
      RECT 125.665 25.005 126.875 27.355 ;
      RECT 123.825 25.005 125.495 27.355 ;
      RECT 118.305 25.005 123.65 27.355 ;
      RECT 109.105 25.005 110.315 27.355 ;
      RECT 103.585 25.005 108.93 27.355 ;
      RECT 101.745 25.005 102.955 27.355 ;
      RECT 102.205 24.485 102.955 27.355 ;
      RECT 99.905 24.485 101.115 27.355 ;
      RECT 94.385 26.095 99.73 27.355 ;
      RECT 88.865 26.095 94.21 27.355 ;
      RECT 87.025 24.485 88.235 27.355 ;
      RECT 85.185 26.095 86.855 27.355 ;
      RECT 74.145 26.095 77.655 27.355 ;
      RECT 71.385 25.005 72.595 27.355 ;
      RECT 62.185 26.095 63.855 27.355 ;
      RECT 59.425 25.005 62.015 27.355 ;
      RECT 50.225 26.095 51.435 27.355 ;
      RECT 44.705 26.095 50.05 27.355 ;
      RECT 47.235 25.295 47.565 27.355 ;
      RECT 35.505 26.095 36.715 27.355 ;
      RECT 31.805 24.485 33.495 27.355 ;
      RECT 20.785 25.005 21.995 27.355 ;
      RECT 15.265 25.005 20.61 27.355 ;
      RECT 13.425 25.005 14.635 27.355 ;
      RECT 10.665 25.005 13.255 27.355 ;
      RECT 145.005 25.005 145.175 27.275 ;
      RECT 116.945 26.095 117.115 27.275 ;
      RECT 84.285 26.095 84.455 27.275 ;
      RECT 70.485 26.095 70.655 27.275 ;
      RECT 58.065 24.485 58.235 27.275 ;
      RECT 43.345 24.485 43.515 27.275 ;
      RECT 28.625 25.005 28.795 27.275 ;
      RECT 142.07 26.095 142.24 27.065 ;
      RECT 114.01 26.095 114.18 27.065 ;
      RECT 81.35 24.485 81.52 27.065 ;
      RECT 67.55 26.095 67.72 27.065 ;
      RECT 55.13 24.485 55.3 27.065 ;
      RECT 40.41 25.005 40.58 27.065 ;
      RECT 25.69 24.485 25.86 27.065 ;
      RECT 155.54 25.005 155.87 27.025 ;
      RECT 127.49 24.485 127.82 27.025 ;
      RECT 143.95 26.095 144.265 26.765 ;
      RECT 138.975 25.005 139.305 26.765 ;
      RECT 115.89 26.095 116.205 26.765 ;
      RECT 110.915 26.095 111.245 26.765 ;
      RECT 83.23 26.095 83.545 26.765 ;
      RECT 78.255 26.095 78.585 26.765 ;
      RECT 69.43 26.095 69.745 26.765 ;
      RECT 64.455 25.005 64.785 26.765 ;
      RECT 57.01 25.005 57.325 26.765 ;
      RECT 52.035 25.005 52.365 26.765 ;
      RECT 42.29 24.485 42.605 26.765 ;
      RECT 37.315 26.095 37.645 26.765 ;
      RECT 27.57 24.485 27.885 26.765 ;
      RECT 22.595 25.005 22.925 26.765 ;
      RECT 139.9 24.485 140.165 26.725 ;
      RECT 111.84 24.465 112.105 26.725 ;
      RECT 79.18 26.095 79.445 26.725 ;
      RECT 65.38 24.485 65.645 26.725 ;
      RECT 52.96 25.005 53.225 26.725 ;
      RECT 38.24 26.095 38.505 26.725 ;
      RECT 23.52 25.005 23.785 26.725 ;
      RECT 154.595 25.005 154.95 26.685 ;
      RECT 128.41 24.485 128.765 26.685 ;
      RECT 10.12 26.095 189.98 26.265 ;
      RECT 160.625 25.005 161.835 26.265 ;
      RECT 161.315 24.465 161.835 26.265 ;
      RECT 153.265 25.005 158.61 26.265 ;
      RECT 150.495 24.485 153.09 26.265 ;
      RECT 144.525 25.005 147.115 26.265 ;
      RECT 142.21 25.675 142.565 26.265 ;
      RECT 141.29 25.335 141.62 26.265 ;
      RECT 138.085 25.005 140.675 26.265 ;
      RECT 139.465 24.485 140.675 26.265 ;
      RECT 134.85 25.335 135.18 27.355 ;
      RECT 133.025 25.005 134.235 27.355 ;
      RECT 133.715 24.465 134.235 27.355 ;
      RECT 129.345 25.005 131.015 26.265 ;
      RECT 123.825 25.005 129.17 26.265 ;
      RECT 126.575 24.485 129.17 26.265 ;
      RECT 116.955 24.945 117.285 26.265 ;
      RECT 116.115 25.295 116.445 26.265 ;
      RECT 115.275 25.295 115.605 26.265 ;
      RECT 114.435 25.295 114.765 26.265 ;
      RECT 113.675 25.295 113.845 26.265 ;
      RECT 112.835 25.295 113.005 26.265 ;
      RECT 110.945 25.005 112.155 26.265 ;
      RECT 111.635 24.465 112.155 26.265 ;
      RECT 110.025 24.485 110.775 26.265 ;
      RECT 101.285 25.005 102.955 26.265 ;
      RECT 98.525 25.005 101.115 26.265 ;
      RECT 97.58 25.335 97.91 27.875 ;
      RECT 96.635 25.675 96.99 27.355 ;
      RECT 93.465 25.005 94.675 26.265 ;
      RECT 91.625 25.005 93.295 27.875 ;
      RECT 92.545 24.485 93.295 27.875 ;
      RECT 88.865 25.005 91.455 27.355 ;
      RECT 90.245 24.485 91.455 27.355 ;
      RECT 85.645 25.005 88.235 26.265 ;
      RECT 83.33 25.675 83.685 26.265 ;
      RECT 82.41 25.335 82.74 26.265 ;
      RECT 79.205 25.005 81.795 26.265 ;
      RECT 80.585 24.485 81.795 26.265 ;
      RECT 76.89 25.675 77.245 27.875 ;
      RECT 75.97 25.335 76.3 27.875 ;
      RECT 74.145 25.005 75.355 27.355 ;
      RECT 74.835 24.465 75.355 27.355 ;
      RECT 70.925 25.005 73.515 26.265 ;
      RECT 72.305 24.485 73.515 26.265 ;
      RECT 68.61 25.675 68.965 26.265 ;
      RECT 67.69 25.335 68.02 26.265 ;
      RECT 65.865 25.005 67.075 26.265 ;
      RECT 66.555 24.465 67.075 26.265 ;
      RECT 63.105 25.005 65.695 26.265 ;
      RECT 64.485 24.485 65.695 26.265 ;
      RECT 56.205 25.005 58.795 26.265 ;
      RECT 57.585 24.485 58.795 26.265 ;
      RECT 50.685 25.005 56.03 26.265 ;
      RECT 53.435 24.485 56.03 26.265 ;
      RECT 49.835 25.295 50.005 27.875 ;
      RECT 48.995 25.295 49.165 27.875 ;
      RECT 48.075 25.295 48.405 27.875 ;
      RECT 46.395 25.295 46.725 27.355 ;
      RECT 45.555 24.945 45.885 27.355 ;
      RECT 38.725 25.005 44.07 26.265 ;
      RECT 41.475 24.485 44.07 26.265 ;
      RECT 37.78 25.335 38.11 26.265 ;
      RECT 36.835 25.675 37.19 26.265 ;
      RECT 33.665 25.005 34.875 27.875 ;
      RECT 34.355 24.465 34.875 27.875 ;
      RECT 29.985 25.005 33.495 27.355 ;
      RECT 28.145 25.005 29.355 26.265 ;
      RECT 28.835 24.465 29.355 26.265 ;
      RECT 26.305 25.005 27.975 26.265 ;
      RECT 27.225 24.485 27.975 26.265 ;
      RECT 20.785 25.005 26.13 26.265 ;
      RECT 23.535 24.485 26.13 26.265 ;
      RECT 159.705 24.485 160.455 27.875 ;
      RECT 156.015 24.485 158.61 26.265 ;
      RECT 130.265 24.485 131.015 26.265 ;
      RECT 94.155 24.465 94.675 26.265 ;
      RECT 61.245 24.485 62.935 26.265 ;
      RECT 186.385 27.525 187.595 30.275 ;
      RECT 182.705 27.525 184.355 30.275 ;
      RECT 177.185 27.525 179.765 30.275 ;
      RECT 169.825 27.525 170.345 30.275 ;
      RECT 167.985 27.525 168.735 30.275 ;
      RECT 162.465 27.525 165.045 30.275 ;
      RECT 158.325 28.045 159.975 30.275 ;
      RECT 149.585 28.045 150.105 30.275 ;
      RECT 147.745 27.525 148.495 30.275 ;
      RECT 145.905 27.525 146.425 30.275 ;
      RECT 144.065 28.815 144.815 30.275 ;
      RECT 138.545 28.815 141.125 30.275 ;
      RECT 133.025 27.525 135.605 30.275 ;
      RECT 131.185 28.045 131.705 30.275 ;
      RECT 129.345 28.815 130.095 30.275 ;
      RECT 123.825 28.815 126.405 30.275 ;
      RECT 118.305 27.525 120.885 30.275 ;
      RECT 116.465 28.815 116.985 30.275 ;
      RECT 114.625 28.815 115.375 30.275 ;
      RECT 103.585 27.525 105.235 30.275 ;
      RECT 101.745 27.525 102.265 30.275 ;
      RECT 99.905 27.525 100.655 30.275 ;
      RECT 94.385 27.525 96.965 30.275 ;
      RECT 88.865 27.525 91.445 30.275 ;
      RECT 87.025 27.525 87.545 30.275 ;
      RECT 85.185 27.525 85.935 30.275 ;
      RECT 79.665 28.815 82.245 30.275 ;
      RECT 74.145 28.045 76.725 30.275 ;
      RECT 72.305 28.815 72.825 30.275 ;
      RECT 70.465 28.815 71.215 30.275 ;
      RECT 64.945 28.815 67.525 30.275 ;
      RECT 59.425 28.045 62.005 30.275 ;
      RECT 57.585 28.815 58.105 30.275 ;
      RECT 55.745 28.815 56.495 30.275 ;
      RECT 50.225 28.815 52.805 30.275 ;
      RECT 44.705 27.525 47.285 30.275 ;
      RECT 38.725 28.815 41.305 30.275 ;
      RECT 33.665 28.045 34.185 30.275 ;
      RECT 29.985 27.525 31.635 30.275 ;
      RECT 28.145 28.815 28.665 30.275 ;
      RECT 26.305 28.815 27.055 30.275 ;
      RECT 20.785 28.815 23.365 30.275 ;
      RECT 15.265 27.525 17.845 30.275 ;
      RECT 13.425 27.525 13.945 30.275 ;
      RECT 10.665 27.525 11.875 30.275 ;
      RECT 175.835 28.065 176.165 29.785 ;
      RECT 186.385 28.045 188.975 29.755 ;
      RECT 182.705 28.045 186.215 29.755 ;
      RECT 177.185 28.045 182.53 29.755 ;
      RECT 167.985 27.525 169.655 29.755 ;
      RECT 162.465 28.045 167.81 29.755 ;
      RECT 158.325 28.815 161.835 29.755 ;
      RECT 147.745 28.045 149.415 29.755 ;
      RECT 144.065 28.815 145.735 29.755 ;
      RECT 138.545 28.815 143.89 29.755 ;
      RECT 133.025 28.045 138.37 29.755 ;
      RECT 129.345 28.815 131.015 29.755 ;
      RECT 123.825 28.815 129.17 29.755 ;
      RECT 118.305 28.045 123.65 29.755 ;
      RECT 114.625 28.815 116.295 29.755 ;
      RECT 103.585 28.045 107.095 29.755 ;
      RECT 99.905 28.045 101.575 29.755 ;
      RECT 94.385 28.045 99.73 29.755 ;
      RECT 88.865 28.045 94.21 29.755 ;
      RECT 85.185 28.045 86.855 29.755 ;
      RECT 79.665 28.815 85.01 29.755 ;
      RECT 74.145 28.815 79.49 29.755 ;
      RECT 70.465 28.815 72.135 29.755 ;
      RECT 64.945 28.815 70.29 29.755 ;
      RECT 59.425 28.815 64.77 29.755 ;
      RECT 55.745 28.815 57.415 29.755 ;
      RECT 50.225 28.815 55.57 29.755 ;
      RECT 44.705 28.045 50.05 29.755 ;
      RECT 38.725 28.815 44.07 29.755 ;
      RECT 29.985 28.045 33.495 29.755 ;
      RECT 26.305 28.815 27.975 29.755 ;
      RECT 20.785 28.815 26.13 29.755 ;
      RECT 15.265 28.045 20.61 29.755 ;
      RECT 10.665 28.045 13.255 29.755 ;
      RECT 169.825 28.045 171.035 29.735 ;
      RECT 149.585 28.045 150.795 29.735 ;
      RECT 145.905 28.065 147.115 29.735 ;
      RECT 131.185 28.045 132.395 29.735 ;
      RECT 116.465 28.815 117.675 29.735 ;
      RECT 101.745 28.065 102.955 29.735 ;
      RECT 87.025 28.065 88.235 29.735 ;
      RECT 72.305 28.815 73.515 29.735 ;
      RECT 57.585 28.815 58.795 29.735 ;
      RECT 33.665 28.045 34.875 29.735 ;
      RECT 28.145 28.815 29.355 29.735 ;
      RECT 13.425 28.065 14.635 29.735 ;
      RECT 189.605 28.09 189.895 29.71 ;
      RECT 189.145 28.09 189.435 29.71 ;
      RECT 176.725 28.09 177.015 29.71 ;
      RECT 162.005 28.09 162.295 29.71 ;
      RECT 147.285 28.09 147.575 29.71 ;
      RECT 132.565 28.09 132.855 29.71 ;
      RECT 117.845 28.09 118.135 29.71 ;
      RECT 103.125 28.09 103.415 29.71 ;
      RECT 88.405 28.09 88.695 29.71 ;
      RECT 73.685 28.09 73.975 29.71 ;
      RECT 58.965 28.09 59.255 29.71 ;
      RECT 44.245 28.09 44.535 29.71 ;
      RECT 29.525 28.09 29.815 29.71 ;
      RECT 14.805 28.09 15.095 29.71 ;
      RECT 10.205 28.09 10.495 29.71 ;
      RECT 157.435 27.525 157.605 29.595 ;
      RECT 113.735 28.815 113.905 29.595 ;
      RECT 156.465 28.815 156.675 29.515 ;
      RECT 112.765 28.815 112.975 29.515 ;
      RECT 154.28 28.815 154.65 29.485 ;
      RECT 110.58 28.815 110.95 29.485 ;
      RECT 174.995 28.815 175.325 29.465 ;
      RECT 174.155 28.045 174.485 29.465 ;
      RECT 173.315 28.815 173.645 29.465 ;
      RECT 172.475 28.045 172.805 29.465 ;
      RECT 171.635 28.045 171.965 29.465 ;
      RECT 37.735 28.815 38.065 29.465 ;
      RECT 35.475 28.815 35.805 29.465 ;
      RECT 152.335 28.065 152.585 29.445 ;
      RECT 108.635 28.045 108.885 29.445 ;
      RECT 151.395 28.815 151.725 29.365 ;
      RECT 107.695 28.045 108.025 29.365 ;
      RECT 10.12 28.815 189.98 28.985 ;
      RECT 175.345 28.065 176.555 28.985 ;
      RECT 173.505 28.045 175.175 28.985 ;
      RECT 167.985 28.045 173.33 28.985 ;
      RECT 156.485 28.045 161.83 28.985 ;
      RECT 155.495 28.335 155.825 28.985 ;
      RECT 153.235 28.335 153.565 28.985 ;
      RECT 151.425 28.065 152.635 28.985 ;
      RECT 147.745 28.045 151.255 28.985 ;
      RECT 145.015 28.205 145.185 29.755 ;
      RECT 144.045 28.285 144.255 28.985 ;
      RECT 141.86 28.315 142.23 29.755 ;
      RECT 139.915 28.355 140.165 30.275 ;
      RECT 138.975 28.435 139.305 30.275 ;
      RECT 130.725 27.525 131.475 28.985 ;
      RECT 129.795 28.335 130.125 29.755 ;
      RECT 127.535 28.335 127.865 29.755 ;
      RECT 125.665 28.065 126.875 29.755 ;
      RECT 123.825 28.045 125.495 30.275 ;
      RECT 116.955 28.205 117.125 29.735 ;
      RECT 115.985 28.285 116.195 29.755 ;
      RECT 113.8 28.315 114.17 28.985 ;
      RECT 111.855 28.355 112.105 28.985 ;
      RECT 110.915 28.435 111.245 28.985 ;
      RECT 109.105 28.065 110.315 28.985 ;
      RECT 103.585 28.045 108.93 28.985 ;
      RECT 84.295 28.205 84.465 29.755 ;
      RECT 83.325 28.285 83.535 29.755 ;
      RECT 81.14 28.315 81.51 30.275 ;
      RECT 79.195 28.355 79.445 29.755 ;
      RECT 78.255 28.435 78.585 29.755 ;
      RECT 74.145 28.045 77.655 29.755 ;
      RECT 71.385 28.065 72.595 28.985 ;
      RECT 70.495 28.205 70.665 30.275 ;
      RECT 69.525 28.285 69.735 29.755 ;
      RECT 67.34 28.315 67.71 29.755 ;
      RECT 65.395 28.355 65.645 30.275 ;
      RECT 64.455 28.435 64.785 28.985 ;
      RECT 62.185 28.045 63.855 29.755 ;
      RECT 59.425 28.045 62.015 29.755 ;
      RECT 58.075 28.205 58.245 29.735 ;
      RECT 57.105 28.285 57.315 29.755 ;
      RECT 54.92 28.315 55.29 29.755 ;
      RECT 52.975 28.355 53.225 29.755 ;
      RECT 52.035 28.435 52.365 30.275 ;
      RECT 50.225 28.065 51.435 30.275 ;
      RECT 43.355 28.205 43.525 29.755 ;
      RECT 42.385 28.285 42.595 29.755 ;
      RECT 40.2 28.315 40.57 30.275 ;
      RECT 38.255 28.355 38.505 28.985 ;
      RECT 37.315 28.435 37.645 28.985 ;
      RECT 35.505 28.065 36.715 28.985 ;
      RECT 29.985 28.045 35.33 28.985 ;
      RECT 28.635 28.205 28.805 29.735 ;
      RECT 27.665 28.285 27.875 29.755 ;
      RECT 25.48 28.315 25.85 29.755 ;
      RECT 23.535 28.355 23.785 29.755 ;
      RECT 22.595 28.435 22.925 30.275 ;
      RECT 20.785 28.065 21.995 30.275 ;
      RECT 175.345 27.525 175.865 28.985 ;
      RECT 151.425 27.525 151.945 28.985 ;
      RECT 125.665 27.525 126.185 30.275 ;
      RECT 109.105 27.525 109.625 28.985 ;
      RECT 71.385 27.525 71.905 29.755 ;
      RECT 50.225 27.525 50.745 30.275 ;
      RECT 35.505 27.525 36.025 28.985 ;
      RECT 20.785 27.525 21.305 30.275 ;
      RECT 173.505 27.525 174.255 28.985 ;
      RECT 167.985 27.525 170.565 28.985 ;
      RECT 156.485 27.525 159.065 28.985 ;
      RECT 147.745 27.525 149.395 29.755 ;
      RECT 123.825 27.525 124.575 30.275 ;
      RECT 103.585 27.525 106.165 29.755 ;
      RECT 74.145 27.525 75.795 30.275 ;
      RECT 62.185 27.525 62.935 29.755 ;
      RECT 59.425 27.525 60.635 30.275 ;
      RECT 29.985 27.525 32.565 29.755 ;
      RECT 176.035 31.535 176.555 33.335 ;
      RECT 152.115 31.535 152.635 33.335 ;
      RECT 146.595 29.905 147.115 33.335 ;
      RECT 131.875 29.905 132.395 33.335 ;
      RECT 117.155 29.905 117.675 33.335 ;
      RECT 94.155 31.535 94.675 33.335 ;
      RECT 87.715 29.905 88.235 33.335 ;
      RECT 72.995 29.905 73.515 33.335 ;
      RECT 58.275 29.905 58.795 33.335 ;
      RECT 34.355 29.905 34.875 33.335 ;
      RECT 28.835 29.905 29.355 33.335 ;
      RECT 14.115 29.905 14.635 33.335 ;
      RECT 187.765 29.925 188.975 33.315 ;
      RECT 184.525 29.925 186.215 33.315 ;
      RECT 179.935 29.925 182.53 33.315 ;
      RECT 174.425 31.535 175.175 33.315 ;
      RECT 170.735 31.535 173.33 33.315 ;
      RECT 165.215 29.925 167.81 33.315 ;
      RECT 159.235 30.445 161.83 33.315 ;
      RECT 149.565 31.535 151.255 33.315 ;
      RECT 144.985 29.925 145.735 33.315 ;
      RECT 141.295 29.925 143.89 33.315 ;
      RECT 135.775 29.925 138.37 33.315 ;
      RECT 130.265 29.925 131.015 33.315 ;
      RECT 126.575 29.925 129.17 33.315 ;
      RECT 121.055 29.925 123.65 33.315 ;
      RECT 115.545 29.925 116.295 33.315 ;
      RECT 111.855 31.535 114.45 33.315 ;
      RECT 106.335 31.535 108.93 33.315 ;
      RECT 102.205 30.445 102.955 33.315 ;
      RECT 102.435 29.905 102.955 33.315 ;
      RECT 99.905 30.445 101.115 33.315 ;
      RECT 92.545 29.925 93.295 33.315 ;
      RECT 90.245 30.445 91.455 33.315 ;
      RECT 86.105 29.925 86.855 33.315 ;
      RECT 83.805 31.535 85.015 33.315 ;
      RECT 71.385 29.925 72.135 33.315 ;
      RECT 67.695 29.925 70.29 33.315 ;
      RECT 62.175 29.925 64.77 33.315 ;
      RECT 56.665 29.925 57.415 33.315 ;
      RECT 52.975 29.925 55.57 33.315 ;
      RECT 47.455 29.925 50.05 33.315 ;
      RECT 41.475 29.925 44.07 33.315 ;
      RECT 31.805 29.925 33.495 33.315 ;
      RECT 27.225 29.925 27.975 33.315 ;
      RECT 23.535 29.925 26.13 33.315 ;
      RECT 18.015 29.925 20.61 33.315 ;
      RECT 12.045 29.925 13.255 33.315 ;
      RECT 189.605 30.37 189.895 32.87 ;
      RECT 189.145 30.37 189.435 32.87 ;
      RECT 176.725 30.37 177.015 32.87 ;
      RECT 162.005 30.37 162.295 32.87 ;
      RECT 147.285 30.37 147.575 32.87 ;
      RECT 132.565 30.37 132.855 32.87 ;
      RECT 117.845 30.37 118.135 32.87 ;
      RECT 103.125 30.37 103.415 32.87 ;
      RECT 88.405 30.37 88.695 32.87 ;
      RECT 73.685 30.37 73.975 32.87 ;
      RECT 58.965 30.37 59.255 32.87 ;
      RECT 44.245 30.37 44.535 32.87 ;
      RECT 29.525 30.37 29.815 32.87 ;
      RECT 14.805 30.37 15.095 32.87 ;
      RECT 10.205 30.37 10.495 32.87 ;
      RECT 186.385 30.445 188.975 32.795 ;
      RECT 182.705 30.445 186.215 32.795 ;
      RECT 177.185 30.445 182.53 32.795 ;
      RECT 175.345 31.535 176.555 32.795 ;
      RECT 175.835 30.385 176.165 32.795 ;
      RECT 173.505 31.535 175.175 32.795 ;
      RECT 174.155 30.735 174.485 32.795 ;
      RECT 167.985 31.535 173.33 32.795 ;
      RECT 170.515 29.905 171.035 32.795 ;
      RECT 162.465 30.445 167.81 32.795 ;
      RECT 156.485 31.535 161.83 32.795 ;
      RECT 158.325 30.445 161.83 32.795 ;
      RECT 151.425 31.535 152.635 32.795 ;
      RECT 147.745 31.535 151.255 32.795 ;
      RECT 145.905 30.445 147.115 32.795 ;
      RECT 144.065 30.445 145.735 32.795 ;
      RECT 138.545 30.445 143.89 32.795 ;
      RECT 133.025 30.445 138.37 32.795 ;
      RECT 131.185 30.445 132.395 32.795 ;
      RECT 129.345 30.445 131.015 32.795 ;
      RECT 123.825 30.445 129.17 32.795 ;
      RECT 118.305 30.445 123.65 32.795 ;
      RECT 116.465 30.445 117.675 32.795 ;
      RECT 114.625 30.445 116.295 32.795 ;
      RECT 109.105 31.535 114.45 32.795 ;
      RECT 105.405 29.925 107.095 32.795 ;
      RECT 101.285 31.535 102.955 32.795 ;
      RECT 101.745 30.445 102.955 32.795 ;
      RECT 98.525 31.535 101.115 32.795 ;
      RECT 93.465 31.535 94.675 32.795 ;
      RECT 91.625 29.925 93.295 32.795 ;
      RECT 88.865 30.445 91.455 32.795 ;
      RECT 87.025 30.445 88.235 32.795 ;
      RECT 85.185 30.445 86.855 32.795 ;
      RECT 82.425 31.535 85.015 32.795 ;
      RECT 72.305 30.445 73.515 32.795 ;
      RECT 70.465 30.445 72.135 32.795 ;
      RECT 64.945 30.445 70.29 32.795 ;
      RECT 59.425 30.445 64.77 32.795 ;
      RECT 57.585 30.445 58.795 32.795 ;
      RECT 55.745 30.445 57.415 32.795 ;
      RECT 50.225 30.445 55.57 32.795 ;
      RECT 44.705 30.445 50.05 32.795 ;
      RECT 38.725 30.445 44.07 32.795 ;
      RECT 33.665 30.445 34.875 32.795 ;
      RECT 29.985 30.445 33.495 32.795 ;
      RECT 28.145 30.445 29.355 32.795 ;
      RECT 26.305 30.445 27.975 32.795 ;
      RECT 20.785 30.445 26.13 32.795 ;
      RECT 15.265 30.445 20.61 32.795 ;
      RECT 13.425 30.445 14.635 32.795 ;
      RECT 10.665 30.445 13.255 32.795 ;
      RECT 81.525 30.445 81.695 32.715 ;
      RECT 78.59 29.925 78.76 32.505 ;
      RECT 155.54 31.535 155.87 32.465 ;
      RECT 97.58 29.925 97.91 32.465 ;
      RECT 37.78 30.775 38.11 32.465 ;
      RECT 80.47 30.445 80.785 32.205 ;
      RECT 75.495 30.445 75.825 32.205 ;
      RECT 76.42 30.445 76.685 32.165 ;
      RECT 154.595 31.535 154.95 32.125 ;
      RECT 96.635 30.445 96.99 32.125 ;
      RECT 36.835 31.115 37.19 32.125 ;
      RECT 10.12 31.535 189.98 31.705 ;
      RECT 174.995 30.735 175.325 31.705 ;
      RECT 173.315 30.735 173.645 31.705 ;
      RECT 172.555 30.735 172.725 33.315 ;
      RECT 171.715 30.735 171.885 33.315 ;
      RECT 169.825 30.445 171.035 32.795 ;
      RECT 167.985 30.445 169.655 32.795 ;
      RECT 168.905 29.925 169.655 32.795 ;
      RECT 160.145 29.925 161.835 31.705 ;
      RECT 157.425 30.525 157.595 32.795 ;
      RECT 156.37 31.035 156.685 31.705 ;
      RECT 154.49 30.735 154.66 31.705 ;
      RECT 152.32 31.075 152.585 33.335 ;
      RECT 151.395 31.035 151.725 31.705 ;
      RECT 149.585 30.445 150.795 33.315 ;
      RECT 150.275 29.905 150.795 33.315 ;
      RECT 147.745 30.445 149.415 32.795 ;
      RECT 148.665 29.925 149.415 32.795 ;
      RECT 113.725 30.525 113.895 33.315 ;
      RECT 112.67 31.035 112.985 33.315 ;
      RECT 110.79 30.735 110.96 32.795 ;
      RECT 108.62 31.075 108.885 33.315 ;
      RECT 107.695 31.035 108.025 33.315 ;
      RECT 103.585 30.445 107.095 32.795 ;
      RECT 94.385 30.445 99.73 31.705 ;
      RECT 88.865 30.445 94.21 31.705 ;
      RECT 91.615 29.925 94.21 31.705 ;
      RECT 79.665 30.445 85.01 31.705 ;
      RECT 82.415 29.925 85.01 31.705 ;
      RECT 74.145 30.445 79.49 31.705 ;
      RECT 76.895 29.925 79.49 31.705 ;
      RECT 100.825 29.925 101.575 31.705 ;
      RECT 97.135 29.925 99.73 31.705 ;
      RECT 186.385 32.965 187.595 35.715 ;
      RECT 182.705 32.965 184.355 35.715 ;
      RECT 177.185 32.965 179.765 35.715 ;
      RECT 175.345 32.965 175.865 35.715 ;
      RECT 173.505 32.965 174.255 35.715 ;
      RECT 167.985 32.965 170.565 35.715 ;
      RECT 162.465 32.965 165.045 35.715 ;
      RECT 160.625 33.485 161.145 35.715 ;
      RECT 158.785 33.485 159.535 35.715 ;
      RECT 147.745 32.965 149.395 35.715 ;
      RECT 145.905 32.965 146.425 35.715 ;
      RECT 144.065 32.965 144.815 35.715 ;
      RECT 138.545 32.965 141.125 35.715 ;
      RECT 133.025 32.965 135.605 35.715 ;
      RECT 122.905 33.485 123.425 35.715 ;
      RECT 121.065 33.485 121.815 35.715 ;
      RECT 118.305 32.965 119.515 35.715 ;
      RECT 116.465 32.965 116.985 35.715 ;
      RECT 114.625 32.965 115.375 35.715 ;
      RECT 109.105 32.965 111.685 35.715 ;
      RECT 103.585 32.965 106.165 35.715 ;
      RECT 100.365 34.255 101.575 35.715 ;
      RECT 91.625 32.965 92.145 35.715 ;
      RECT 88.865 32.965 90.075 35.715 ;
      RECT 87.025 32.965 87.545 35.715 ;
      RECT 85.185 32.965 85.935 35.715 ;
      RECT 79.665 34.255 82.245 35.715 ;
      RECT 74.145 34.255 76.725 35.715 ;
      RECT 72.305 32.965 72.825 35.715 ;
      RECT 70.465 32.965 71.215 35.715 ;
      RECT 64.945 32.965 67.525 35.715 ;
      RECT 59.425 32.965 62.005 35.715 ;
      RECT 57.585 32.965 58.105 35.715 ;
      RECT 55.745 32.965 56.495 35.715 ;
      RECT 50.225 32.965 52.805 35.715 ;
      RECT 44.705 32.965 47.285 35.715 ;
      RECT 40.565 33.485 42.215 35.715 ;
      RECT 31.825 33.485 32.345 35.715 ;
      RECT 29.985 32.965 30.735 35.715 ;
      RECT 28.145 32.965 28.665 35.715 ;
      RECT 26.305 32.965 27.055 35.715 ;
      RECT 20.785 32.965 23.365 35.715 ;
      RECT 15.265 32.965 17.845 35.715 ;
      RECT 13.425 32.965 13.945 35.715 ;
      RECT 10.665 32.965 11.875 35.715 ;
      RECT 186.385 33.485 188.975 35.195 ;
      RECT 182.705 33.485 186.215 35.195 ;
      RECT 177.185 33.485 182.53 35.195 ;
      RECT 173.505 33.485 175.175 35.195 ;
      RECT 167.985 33.485 173.33 35.195 ;
      RECT 162.465 33.485 167.81 35.195 ;
      RECT 158.785 33.485 160.455 35.195 ;
      RECT 147.745 33.485 151.255 35.195 ;
      RECT 144.065 33.485 145.735 35.195 ;
      RECT 138.545 33.485 143.89 35.195 ;
      RECT 133.025 33.485 138.37 35.195 ;
      RECT 121.065 33.485 122.735 35.195 ;
      RECT 118.305 33.485 120.895 35.195 ;
      RECT 114.625 33.485 116.295 35.195 ;
      RECT 109.105 33.485 114.45 35.195 ;
      RECT 103.585 33.485 108.93 35.195 ;
      RECT 101.285 33.485 102.955 35.195 ;
      RECT 88.865 33.485 91.455 35.195 ;
      RECT 85.185 33.485 86.855 35.195 ;
      RECT 79.665 34.255 85.01 35.195 ;
      RECT 74.145 34.255 79.49 35.195 ;
      RECT 70.465 33.485 72.135 35.195 ;
      RECT 64.945 33.485 70.29 35.195 ;
      RECT 59.425 33.485 64.77 35.195 ;
      RECT 55.745 33.485 57.415 35.195 ;
      RECT 50.225 33.485 55.57 35.195 ;
      RECT 44.705 33.485 50.05 35.195 ;
      RECT 40.565 34.255 44.075 35.195 ;
      RECT 29.985 33.485 31.655 35.195 ;
      RECT 26.305 33.485 27.975 35.195 ;
      RECT 20.785 33.485 26.13 35.195 ;
      RECT 15.265 33.485 20.61 35.195 ;
      RECT 10.665 33.485 13.255 35.195 ;
      RECT 175.345 33.505 176.555 35.175 ;
      RECT 160.625 34.255 161.835 35.175 ;
      RECT 145.905 33.505 147.115 35.175 ;
      RECT 122.905 34.255 124.115 35.175 ;
      RECT 116.465 33.505 117.675 35.175 ;
      RECT 91.625 33.485 92.835 35.175 ;
      RECT 87.025 33.505 88.235 35.175 ;
      RECT 72.305 33.505 73.515 35.175 ;
      RECT 57.585 33.505 58.795 35.175 ;
      RECT 31.825 33.485 33.035 35.175 ;
      RECT 28.145 33.505 29.355 35.175 ;
      RECT 13.425 33.505 14.635 35.175 ;
      RECT 189.605 33.53 189.895 35.15 ;
      RECT 189.145 33.53 189.435 35.15 ;
      RECT 176.725 33.53 177.015 35.15 ;
      RECT 162.005 33.53 162.295 35.15 ;
      RECT 147.285 33.53 147.575 35.15 ;
      RECT 132.565 33.53 132.855 35.15 ;
      RECT 117.845 33.53 118.135 35.15 ;
      RECT 103.125 33.53 103.415 35.15 ;
      RECT 88.405 33.53 88.695 35.15 ;
      RECT 73.685 33.53 73.975 35.15 ;
      RECT 58.965 33.53 59.255 35.15 ;
      RECT 44.245 33.53 44.535 35.15 ;
      RECT 29.525 33.53 29.815 35.15 ;
      RECT 14.805 33.53 15.095 35.15 ;
      RECT 10.205 33.53 10.495 35.15 ;
      RECT 157.895 32.965 158.065 35.035 ;
      RECT 130.755 33.485 130.925 35.035 ;
      RECT 99.475 32.965 99.645 35.035 ;
      RECT 39.675 32.965 39.845 35.035 ;
      RECT 156.925 32.965 157.135 34.955 ;
      RECT 129.785 32.965 129.995 34.955 ;
      RECT 98.505 34.255 98.715 34.955 ;
      RECT 38.705 34.255 38.915 34.955 ;
      RECT 154.74 34.255 155.11 34.925 ;
      RECT 127.6 33.485 127.97 34.925 ;
      RECT 96.32 34.255 96.69 34.925 ;
      RECT 36.52 34.255 36.89 34.925 ;
      RECT 152.795 34.255 153.045 34.885 ;
      RECT 125.655 32.965 125.905 34.885 ;
      RECT 94.375 33.505 94.625 34.885 ;
      RECT 34.575 33.505 34.825 34.885 ;
      RECT 151.855 33.505 152.185 34.805 ;
      RECT 124.715 32.965 125.045 34.805 ;
      RECT 93.435 34.255 93.765 34.805 ;
      RECT 33.635 34.255 33.965 34.805 ;
      RECT 10.12 34.255 189.98 34.425 ;
      RECT 156.485 33.485 161.83 34.425 ;
      RECT 155.495 33.775 155.825 34.425 ;
      RECT 153.235 33.775 153.565 34.425 ;
      RECT 151.425 33.505 152.635 34.425 ;
      RECT 131.185 33.505 132.395 34.425 ;
      RECT 129.345 33.485 131.015 34.425 ;
      RECT 123.825 33.485 129.17 34.425 ;
      RECT 118.305 33.485 123.65 34.425 ;
      RECT 98.525 33.485 101.115 34.425 ;
      RECT 97.535 33.775 97.865 34.425 ;
      RECT 95.275 33.775 95.605 34.425 ;
      RECT 93.465 33.505 94.675 34.425 ;
      RECT 91.625 33.485 93.295 34.425 ;
      RECT 82.425 33.485 85.015 34.425 ;
      RECT 81.535 33.645 81.705 35.715 ;
      RECT 80.565 33.725 80.775 35.715 ;
      RECT 78.38 33.755 78.75 35.195 ;
      RECT 76.435 33.795 76.685 35.715 ;
      RECT 75.495 33.875 75.825 35.715 ;
      RECT 38.725 33.485 44.07 34.425 ;
      RECT 37.735 33.775 38.065 34.425 ;
      RECT 35.475 33.775 35.805 34.425 ;
      RECT 33.665 33.505 34.875 34.425 ;
      RECT 29.985 33.485 33.495 34.425 ;
      RECT 151.425 32.965 151.945 34.425 ;
      RECT 131.185 32.965 131.705 34.425 ;
      RECT 93.465 32.965 93.985 34.425 ;
      RECT 33.665 32.965 34.185 34.425 ;
      RECT 156.485 32.965 159.065 34.425 ;
      RECT 129.345 32.965 130.095 34.425 ;
      RECT 123.825 32.965 126.405 34.425 ;
      RECT 118.305 32.965 120.885 35.195 ;
      RECT 101.285 32.965 102.035 35.195 ;
      RECT 98.525 32.965 99.735 34.425 ;
      RECT 91.625 32.965 92.375 35.175 ;
      RECT 82.425 32.965 83.635 35.195 ;
      RECT 38.725 32.965 41.305 34.425 ;
      RECT 29.985 32.965 31.635 35.195 ;
      RECT 176.035 35.345 176.555 38.775 ;
      RECT 161.315 35.345 161.835 38.775 ;
      RECT 146.595 35.345 147.115 38.775 ;
      RECT 131.875 36.975 132.395 38.775 ;
      RECT 117.155 35.345 117.675 38.775 ;
      RECT 102.435 35.365 102.955 38.775 ;
      RECT 87.715 35.345 88.235 38.775 ;
      RECT 72.075 36.975 72.595 38.775 ;
      RECT 58.275 35.345 58.795 38.775 ;
      RECT 43.555 35.365 44.075 38.775 ;
      RECT 28.835 35.345 29.355 38.775 ;
      RECT 14.115 35.345 14.635 38.775 ;
      RECT 187.765 35.365 188.975 38.755 ;
      RECT 184.525 35.365 186.215 38.755 ;
      RECT 179.935 35.365 182.53 38.755 ;
      RECT 174.425 35.365 175.175 38.755 ;
      RECT 170.735 35.365 173.33 38.755 ;
      RECT 165.215 35.365 167.81 38.755 ;
      RECT 159.705 35.365 160.455 38.755 ;
      RECT 156.015 36.975 158.61 38.755 ;
      RECT 150.495 36.975 153.09 38.755 ;
      RECT 144.985 35.365 145.735 38.755 ;
      RECT 141.295 35.365 143.89 38.755 ;
      RECT 135.775 35.365 138.37 38.755 ;
      RECT 130.265 36.975 131.015 38.755 ;
      RECT 126.575 36.975 129.17 38.755 ;
      RECT 121.055 36.975 123.65 38.755 ;
      RECT 115.545 35.365 116.295 38.755 ;
      RECT 111.855 35.365 114.45 38.755 ;
      RECT 106.335 35.365 108.93 38.755 ;
      RECT 100.825 35.885 101.575 38.755 ;
      RECT 97.135 36.975 99.73 38.755 ;
      RECT 91.615 36.975 94.21 38.755 ;
      RECT 86.105 35.365 86.855 38.755 ;
      RECT 82.415 35.365 85.01 38.755 ;
      RECT 76.895 35.365 79.49 38.755 ;
      RECT 64.485 36.975 65.695 38.755 ;
      RECT 61.245 35.885 62.935 38.755 ;
      RECT 56.665 35.365 57.415 38.755 ;
      RECT 52.975 35.365 55.57 38.755 ;
      RECT 47.455 35.365 50.05 38.755 ;
      RECT 41.945 35.885 42.695 38.755 ;
      RECT 38.255 36.975 40.85 38.755 ;
      RECT 32.735 36.975 35.33 38.755 ;
      RECT 27.225 35.365 27.975 38.755 ;
      RECT 23.535 35.365 26.13 38.755 ;
      RECT 18.015 35.365 20.61 38.755 ;
      RECT 12.045 35.365 13.255 38.755 ;
      RECT 189.605 35.81 189.895 38.31 ;
      RECT 189.145 35.81 189.435 38.31 ;
      RECT 176.725 35.81 177.015 38.31 ;
      RECT 162.005 35.81 162.295 38.31 ;
      RECT 147.285 35.81 147.575 38.31 ;
      RECT 132.565 35.81 132.855 38.31 ;
      RECT 117.845 35.81 118.135 38.31 ;
      RECT 103.125 35.81 103.415 38.31 ;
      RECT 88.405 35.81 88.695 38.31 ;
      RECT 73.685 35.81 73.975 38.31 ;
      RECT 58.965 35.81 59.255 38.31 ;
      RECT 44.245 35.81 44.535 38.31 ;
      RECT 29.525 35.81 29.815 38.31 ;
      RECT 14.805 35.81 15.095 38.31 ;
      RECT 10.205 35.81 10.495 38.31 ;
      RECT 70.495 35.885 70.825 38.295 ;
      RECT 186.385 35.885 188.975 38.235 ;
      RECT 182.705 35.885 186.215 38.235 ;
      RECT 177.185 35.885 182.53 38.235 ;
      RECT 175.345 35.885 176.555 38.235 ;
      RECT 173.505 35.885 175.175 38.235 ;
      RECT 167.985 35.885 173.33 38.235 ;
      RECT 162.465 35.885 167.81 38.235 ;
      RECT 160.625 35.885 161.835 38.235 ;
      RECT 158.785 35.885 160.455 38.235 ;
      RECT 153.265 36.975 158.61 38.235 ;
      RECT 149.565 35.365 151.255 38.235 ;
      RECT 145.905 35.885 147.115 38.235 ;
      RECT 144.065 35.885 145.735 38.235 ;
      RECT 138.545 35.885 143.89 38.235 ;
      RECT 133.025 35.885 138.37 38.235 ;
      RECT 131.185 36.975 132.395 38.235 ;
      RECT 129.345 36.975 131.015 38.235 ;
      RECT 123.825 36.975 129.17 38.235 ;
      RECT 118.305 36.975 123.65 38.235 ;
      RECT 116.465 35.885 117.675 38.235 ;
      RECT 114.625 35.885 116.295 38.235 ;
      RECT 109.105 35.885 114.45 38.235 ;
      RECT 103.585 35.885 108.93 38.235 ;
      RECT 101.745 35.365 102.955 38.235 ;
      RECT 99.905 36.975 101.575 38.235 ;
      RECT 94.385 36.975 99.73 38.235 ;
      RECT 88.865 36.975 94.21 38.235 ;
      RECT 87.025 35.885 88.235 38.235 ;
      RECT 85.185 35.885 86.855 38.235 ;
      RECT 79.665 35.885 85.01 38.235 ;
      RECT 74.145 35.885 79.49 38.235 ;
      RECT 71.385 35.365 72.135 38.235 ;
      RECT 63.105 36.975 65.695 38.235 ;
      RECT 59.425 35.885 62.935 38.235 ;
      RECT 57.585 35.885 58.795 38.235 ;
      RECT 55.745 35.885 57.415 38.235 ;
      RECT 50.225 35.885 55.57 38.235 ;
      RECT 44.705 35.885 50.05 38.235 ;
      RECT 42.865 35.365 44.075 38.235 ;
      RECT 41.025 35.885 42.695 38.235 ;
      RECT 35.505 36.975 40.85 38.235 ;
      RECT 29.985 36.975 35.33 38.235 ;
      RECT 32.515 35.345 33.035 38.235 ;
      RECT 28.145 35.885 29.355 38.235 ;
      RECT 26.305 35.885 27.975 38.235 ;
      RECT 20.785 35.885 26.13 38.235 ;
      RECT 15.265 35.885 20.61 38.235 ;
      RECT 13.425 35.885 14.635 38.235 ;
      RECT 10.665 35.885 13.255 38.235 ;
      RECT 69.655 35.365 69.985 37.945 ;
      RECT 68.815 35.365 69.145 37.945 ;
      RECT 67.975 35.365 68.305 37.945 ;
      RECT 67.215 35.885 67.385 37.945 ;
      RECT 66.375 35.885 66.545 37.945 ;
      RECT 10.12 36.975 189.98 37.145 ;
      RECT 157.885 35.965 158.055 38.755 ;
      RECT 156.83 36.475 157.145 38.755 ;
      RECT 154.95 36.175 155.12 38.235 ;
      RECT 152.78 36.515 153.045 38.755 ;
      RECT 151.855 36.475 152.185 38.755 ;
      RECT 147.745 35.885 151.255 38.235 ;
      RECT 130.745 35.965 130.915 38.755 ;
      RECT 129.69 36.475 130.005 38.235 ;
      RECT 127.81 36.175 127.98 38.755 ;
      RECT 125.64 36.515 125.905 38.235 ;
      RECT 124.715 36.475 125.045 38.235 ;
      RECT 122.905 35.885 124.115 37.145 ;
      RECT 121.065 35.885 122.735 38.755 ;
      RECT 121.985 35.365 122.735 38.755 ;
      RECT 118.305 35.885 120.895 38.235 ;
      RECT 119.685 35.365 120.895 38.235 ;
      RECT 100.365 35.885 102.955 37.145 ;
      RECT 99.465 35.965 99.635 38.755 ;
      RECT 98.41 36.475 98.725 38.755 ;
      RECT 96.53 36.175 96.7 38.235 ;
      RECT 94.36 36.515 94.625 37.145 ;
      RECT 93.435 36.475 93.765 38.755 ;
      RECT 91.625 35.885 92.835 38.755 ;
      RECT 92.315 35.345 92.835 38.755 ;
      RECT 88.865 35.885 91.455 38.235 ;
      RECT 90.245 35.365 91.455 38.235 ;
      RECT 72.305 35.885 73.515 37.145 ;
      RECT 72.995 35.345 73.515 37.145 ;
      RECT 70.465 35.885 72.135 37.145 ;
      RECT 64.945 35.885 70.29 37.145 ;
      RECT 67.695 35.365 70.29 37.145 ;
      RECT 62.175 35.365 64.77 37.145 ;
      RECT 40.565 35.885 44.075 37.145 ;
      RECT 42.385 35.365 44.075 37.145 ;
      RECT 39.665 35.965 39.835 38.755 ;
      RECT 38.61 36.475 38.925 38.755 ;
      RECT 36.73 36.175 36.9 38.235 ;
      RECT 34.56 36.515 34.825 38.755 ;
      RECT 33.635 36.475 33.965 38.755 ;
      RECT 31.825 35.885 33.035 38.235 ;
      RECT 29.985 35.885 31.655 38.235 ;
      RECT 30.905 35.365 31.655 38.235 ;
      RECT 123.595 35.345 124.115 37.145 ;
      RECT 186.385 38.405 187.595 41.155 ;
      RECT 182.705 38.405 184.355 41.155 ;
      RECT 177.185 38.405 179.765 41.155 ;
      RECT 175.345 38.405 175.865 41.155 ;
      RECT 173.505 38.405 174.255 41.155 ;
      RECT 167.985 38.405 170.565 41.155 ;
      RECT 162.465 38.405 165.045 41.155 ;
      RECT 160.625 38.405 161.145 41.155 ;
      RECT 158.785 38.405 159.535 41.155 ;
      RECT 153.265 38.405 155.845 41.155 ;
      RECT 147.745 38.405 150.325 41.155 ;
      RECT 145.905 38.405 146.425 41.155 ;
      RECT 144.065 38.405 144.815 41.155 ;
      RECT 138.545 38.405 141.125 41.155 ;
      RECT 133.025 38.405 135.605 41.155 ;
      RECT 131.185 38.405 131.705 41.155 ;
      RECT 129.345 38.405 130.095 41.155 ;
      RECT 123.825 38.405 126.405 41.155 ;
      RECT 118.305 38.405 120.885 41.155 ;
      RECT 116.465 38.405 116.985 41.155 ;
      RECT 114.625 38.405 115.375 41.155 ;
      RECT 109.105 38.405 111.685 41.155 ;
      RECT 103.585 38.405 106.165 41.155 ;
      RECT 101.745 38.405 102.265 41.155 ;
      RECT 99.905 38.405 100.655 41.155 ;
      RECT 94.385 38.405 96.965 41.155 ;
      RECT 88.865 38.405 91.445 41.155 ;
      RECT 87.025 38.405 87.545 41.155 ;
      RECT 85.185 38.405 85.935 41.155 ;
      RECT 79.665 38.405 82.245 41.155 ;
      RECT 74.145 38.405 76.725 41.155 ;
      RECT 72.305 39.695 72.825 41.155 ;
      RECT 70.465 39.695 71.215 41.155 ;
      RECT 64.945 39.695 67.525 41.155 ;
      RECT 59.425 38.925 62.005 41.155 ;
      RECT 57.585 38.405 58.105 41.155 ;
      RECT 55.745 38.405 56.495 41.155 ;
      RECT 50.225 38.405 52.805 41.155 ;
      RECT 44.705 38.405 47.285 41.155 ;
      RECT 42.865 38.405 43.385 41.155 ;
      RECT 41.025 38.405 41.775 41.155 ;
      RECT 35.505 38.405 38.085 41.155 ;
      RECT 29.985 38.405 32.565 41.155 ;
      RECT 28.145 38.405 28.665 41.155 ;
      RECT 26.305 38.405 27.055 41.155 ;
      RECT 20.785 38.405 23.365 41.155 ;
      RECT 15.265 38.405 17.845 41.155 ;
      RECT 13.425 38.405 13.945 41.155 ;
      RECT 10.665 38.405 11.875 41.155 ;
      RECT 186.385 38.925 188.975 40.635 ;
      RECT 182.705 38.925 186.215 40.635 ;
      RECT 177.185 38.925 182.53 40.635 ;
      RECT 173.505 38.925 175.175 40.635 ;
      RECT 167.985 38.925 173.33 40.635 ;
      RECT 162.465 38.925 167.81 40.635 ;
      RECT 158.785 38.925 160.455 40.635 ;
      RECT 153.265 38.925 158.61 40.635 ;
      RECT 147.745 38.925 153.09 40.635 ;
      RECT 144.065 38.925 145.735 40.635 ;
      RECT 138.545 38.925 143.89 40.635 ;
      RECT 133.025 38.925 138.37 40.635 ;
      RECT 129.345 38.925 131.015 40.635 ;
      RECT 123.825 38.925 129.17 40.635 ;
      RECT 118.305 38.925 123.65 40.635 ;
      RECT 114.625 38.925 116.295 40.635 ;
      RECT 109.105 38.925 114.45 40.635 ;
      RECT 103.585 38.925 108.93 40.635 ;
      RECT 99.905 38.925 101.575 40.635 ;
      RECT 94.385 38.925 99.73 40.635 ;
      RECT 88.865 38.925 94.21 40.635 ;
      RECT 85.185 38.925 86.855 40.635 ;
      RECT 79.665 38.925 85.01 40.635 ;
      RECT 74.145 38.925 79.49 40.635 ;
      RECT 70.465 39.695 72.135 40.635 ;
      RECT 64.945 39.695 70.29 40.635 ;
      RECT 59.425 39.695 64.77 40.635 ;
      RECT 55.745 38.925 57.415 40.635 ;
      RECT 50.225 38.925 55.57 40.635 ;
      RECT 44.705 38.925 50.05 40.635 ;
      RECT 41.025 38.925 42.695 40.635 ;
      RECT 35.505 38.925 40.85 40.635 ;
      RECT 29.985 38.925 35.33 40.635 ;
      RECT 26.305 38.925 27.975 40.635 ;
      RECT 20.785 38.925 26.13 40.635 ;
      RECT 15.265 38.925 20.61 40.635 ;
      RECT 10.665 38.925 13.255 40.635 ;
      RECT 175.345 38.945 176.555 40.615 ;
      RECT 160.625 38.945 161.835 40.615 ;
      RECT 145.905 38.945 147.115 40.615 ;
      RECT 131.185 38.945 132.395 40.615 ;
      RECT 116.465 38.945 117.675 40.615 ;
      RECT 101.745 38.945 102.955 40.615 ;
      RECT 87.025 38.945 88.235 40.615 ;
      RECT 72.305 39.695 73.515 40.615 ;
      RECT 57.585 38.945 58.795 40.615 ;
      RECT 42.865 38.945 44.075 40.615 ;
      RECT 28.145 38.945 29.355 40.615 ;
      RECT 13.425 38.945 14.635 40.615 ;
      RECT 189.605 38.97 189.895 40.59 ;
      RECT 189.145 38.97 189.435 40.59 ;
      RECT 176.725 38.97 177.015 40.59 ;
      RECT 162.005 38.97 162.295 40.59 ;
      RECT 147.285 38.97 147.575 40.59 ;
      RECT 132.565 38.97 132.855 40.59 ;
      RECT 117.845 38.97 118.135 40.59 ;
      RECT 103.125 38.97 103.415 40.59 ;
      RECT 88.405 38.97 88.695 40.59 ;
      RECT 73.685 38.97 73.975 40.59 ;
      RECT 58.965 38.97 59.255 40.59 ;
      RECT 44.245 38.97 44.535 40.59 ;
      RECT 29.525 38.97 29.815 40.59 ;
      RECT 14.805 38.97 15.095 40.59 ;
      RECT 10.205 38.97 10.495 40.59 ;
      RECT 10.12 39.695 189.98 39.865 ;
      RECT 71.385 38.945 72.595 39.865 ;
      RECT 70.495 38.895 70.825 41.155 ;
      RECT 69.655 39.215 69.985 40.635 ;
      RECT 68.815 39.215 69.145 40.635 ;
      RECT 67.975 39.215 68.305 40.635 ;
      RECT 67.135 39.215 67.465 41.155 ;
      RECT 66.295 39.215 66.625 41.155 ;
      RECT 63.105 38.925 65.695 39.865 ;
      RECT 59.425 38.925 62.935 40.635 ;
      RECT 71.385 38.405 71.905 40.635 ;
      RECT 63.105 38.405 64.315 40.635 ;
      RECT 59.425 38.405 61.075 41.155 ;
      RECT 176.035 40.785 176.555 44.215 ;
      RECT 161.315 40.785 161.835 44.215 ;
      RECT 146.595 40.785 147.115 44.215 ;
      RECT 131.875 40.785 132.395 44.215 ;
      RECT 117.155 40.785 117.675 44.215 ;
      RECT 102.435 40.785 102.955 44.215 ;
      RECT 87.715 40.785 88.235 44.215 ;
      RECT 72.995 40.785 73.515 44.215 ;
      RECT 58.275 40.785 58.795 44.215 ;
      RECT 43.555 40.785 44.075 44.215 ;
      RECT 28.835 40.785 29.355 44.215 ;
      RECT 14.115 40.785 14.635 44.215 ;
      RECT 187.765 40.805 188.975 44.195 ;
      RECT 184.525 40.805 186.215 44.195 ;
      RECT 179.935 40.805 182.53 44.195 ;
      RECT 174.425 40.805 175.175 44.195 ;
      RECT 170.735 40.805 173.33 44.195 ;
      RECT 165.215 40.805 167.81 44.195 ;
      RECT 159.705 40.805 160.455 44.195 ;
      RECT 156.015 40.805 158.61 44.195 ;
      RECT 150.495 40.805 153.09 44.195 ;
      RECT 144.985 40.805 145.735 44.195 ;
      RECT 141.295 40.805 143.89 44.195 ;
      RECT 135.775 40.805 138.37 44.195 ;
      RECT 130.265 40.805 131.015 44.195 ;
      RECT 126.575 40.805 129.17 44.195 ;
      RECT 121.055 40.805 123.65 44.195 ;
      RECT 115.545 40.805 116.295 44.195 ;
      RECT 111.855 40.805 114.45 44.195 ;
      RECT 106.335 40.805 108.93 44.195 ;
      RECT 100.825 40.805 101.575 44.195 ;
      RECT 97.135 40.805 99.73 44.195 ;
      RECT 91.615 40.805 94.21 44.195 ;
      RECT 86.105 40.805 86.855 44.195 ;
      RECT 82.415 40.805 85.01 44.195 ;
      RECT 76.895 40.805 79.49 44.195 ;
      RECT 71.385 40.805 72.135 44.195 ;
      RECT 67.695 40.805 70.29 44.195 ;
      RECT 62.175 40.805 64.77 44.195 ;
      RECT 56.665 40.805 57.415 44.195 ;
      RECT 52.975 40.805 55.57 44.195 ;
      RECT 47.455 40.805 50.05 44.195 ;
      RECT 41.945 40.805 42.695 44.195 ;
      RECT 38.255 40.805 40.85 44.195 ;
      RECT 32.735 40.805 35.33 44.195 ;
      RECT 27.225 40.805 27.975 44.195 ;
      RECT 23.535 40.805 26.13 44.195 ;
      RECT 18.015 40.805 20.61 44.195 ;
      RECT 12.045 40.805 13.255 44.195 ;
      RECT 189.605 41.25 189.895 43.75 ;
      RECT 189.145 41.25 189.435 43.75 ;
      RECT 176.725 41.25 177.015 43.75 ;
      RECT 162.005 41.25 162.295 43.75 ;
      RECT 147.285 41.25 147.575 43.75 ;
      RECT 132.565 41.25 132.855 43.75 ;
      RECT 117.845 41.25 118.135 43.75 ;
      RECT 103.125 41.25 103.415 43.75 ;
      RECT 88.405 41.25 88.695 43.75 ;
      RECT 73.685 41.25 73.975 43.75 ;
      RECT 58.965 41.25 59.255 43.75 ;
      RECT 44.245 41.25 44.535 43.75 ;
      RECT 29.525 41.25 29.815 43.75 ;
      RECT 14.805 41.25 15.095 43.75 ;
      RECT 10.205 41.25 10.495 43.75 ;
      RECT 186.385 41.325 188.975 43.675 ;
      RECT 182.705 41.325 186.215 43.675 ;
      RECT 177.185 41.325 182.53 43.675 ;
      RECT 175.345 41.325 176.555 43.675 ;
      RECT 173.505 41.325 175.175 43.675 ;
      RECT 167.985 41.325 173.33 43.675 ;
      RECT 162.465 41.325 167.81 43.675 ;
      RECT 160.625 41.325 161.835 43.675 ;
      RECT 158.785 41.325 160.455 43.675 ;
      RECT 153.265 41.325 158.61 43.675 ;
      RECT 147.745 41.325 153.09 43.675 ;
      RECT 145.905 41.325 147.115 43.675 ;
      RECT 144.065 41.325 145.735 43.675 ;
      RECT 138.545 41.325 143.89 43.675 ;
      RECT 133.025 41.325 138.37 43.675 ;
      RECT 131.185 41.325 132.395 43.675 ;
      RECT 129.345 41.325 131.015 43.675 ;
      RECT 123.825 41.325 129.17 43.675 ;
      RECT 118.305 41.325 123.65 43.675 ;
      RECT 116.465 41.325 117.675 43.675 ;
      RECT 114.625 41.325 116.295 43.675 ;
      RECT 109.105 41.325 114.45 43.675 ;
      RECT 103.585 41.325 108.93 43.675 ;
      RECT 101.745 41.325 102.955 43.675 ;
      RECT 99.905 41.325 101.575 43.675 ;
      RECT 94.385 41.325 99.73 43.675 ;
      RECT 88.865 41.325 94.21 43.675 ;
      RECT 87.025 41.325 88.235 43.675 ;
      RECT 85.185 41.325 86.855 43.675 ;
      RECT 79.665 41.325 85.01 43.675 ;
      RECT 74.145 41.325 79.49 43.675 ;
      RECT 72.305 41.325 73.515 43.675 ;
      RECT 70.465 41.325 72.135 43.675 ;
      RECT 64.945 41.325 70.29 43.675 ;
      RECT 59.425 41.325 64.77 43.675 ;
      RECT 57.585 41.325 58.795 43.675 ;
      RECT 55.745 41.325 57.415 43.675 ;
      RECT 50.225 41.325 55.57 43.675 ;
      RECT 44.705 41.325 50.05 43.675 ;
      RECT 42.865 41.325 44.075 43.675 ;
      RECT 41.025 41.325 42.695 43.675 ;
      RECT 35.505 41.325 40.85 43.675 ;
      RECT 29.985 41.325 35.33 43.675 ;
      RECT 28.145 41.325 29.355 43.675 ;
      RECT 26.305 41.325 27.975 43.675 ;
      RECT 20.785 41.325 26.13 43.675 ;
      RECT 15.265 41.325 20.61 43.675 ;
      RECT 13.425 41.325 14.635 43.675 ;
      RECT 10.665 41.325 13.255 43.675 ;
      RECT 10.12 42.415 189.98 42.585 ;
      RECT 186.385 43.845 187.595 46.595 ;
      RECT 182.705 43.845 184.355 46.595 ;
      RECT 177.185 43.845 179.765 46.595 ;
      RECT 175.345 43.845 175.865 46.595 ;
      RECT 173.505 43.845 174.255 46.595 ;
      RECT 167.985 43.845 170.565 46.595 ;
      RECT 162.465 43.845 165.045 46.595 ;
      RECT 160.625 43.845 161.145 46.595 ;
      RECT 158.785 43.845 159.535 46.595 ;
      RECT 153.265 43.845 155.845 46.595 ;
      RECT 147.745 43.845 150.325 46.595 ;
      RECT 145.905 43.845 146.425 46.595 ;
      RECT 144.065 43.845 144.815 46.595 ;
      RECT 138.545 43.845 141.125 46.595 ;
      RECT 133.025 43.845 135.605 46.595 ;
      RECT 131.185 43.845 131.705 46.595 ;
      RECT 129.345 43.845 130.095 46.595 ;
      RECT 123.825 43.845 126.405 46.595 ;
      RECT 118.305 43.845 120.885 46.595 ;
      RECT 116.465 43.845 116.985 46.595 ;
      RECT 114.625 43.845 115.375 46.595 ;
      RECT 109.105 43.845 111.685 46.595 ;
      RECT 103.585 43.845 106.165 46.595 ;
      RECT 101.745 43.845 102.265 46.595 ;
      RECT 99.905 43.845 100.655 46.595 ;
      RECT 94.385 43.845 96.965 46.595 ;
      RECT 88.865 43.845 91.445 46.595 ;
      RECT 87.025 43.845 87.545 46.595 ;
      RECT 85.185 43.845 85.935 46.595 ;
      RECT 79.665 43.845 82.245 46.595 ;
      RECT 74.145 43.845 76.725 46.595 ;
      RECT 72.305 43.845 72.825 46.595 ;
      RECT 70.465 43.845 71.215 46.595 ;
      RECT 64.945 43.845 67.525 46.595 ;
      RECT 59.425 43.845 62.005 46.595 ;
      RECT 57.585 43.845 58.105 46.595 ;
      RECT 55.745 43.845 56.495 46.595 ;
      RECT 50.225 43.845 52.805 46.595 ;
      RECT 44.705 43.845 47.285 46.595 ;
      RECT 42.865 43.845 43.385 46.595 ;
      RECT 41.025 43.845 41.775 46.595 ;
      RECT 35.505 43.845 38.085 46.595 ;
      RECT 29.985 43.845 32.565 46.595 ;
      RECT 28.145 43.845 28.665 46.595 ;
      RECT 26.305 43.845 27.055 46.595 ;
      RECT 20.785 43.845 23.365 46.595 ;
      RECT 15.265 43.845 17.845 46.595 ;
      RECT 13.425 43.845 13.945 46.595 ;
      RECT 10.665 43.845 11.875 46.595 ;
      RECT 186.385 44.365 188.975 46.075 ;
      RECT 182.705 44.365 186.215 46.075 ;
      RECT 177.185 44.365 182.53 46.075 ;
      RECT 173.505 44.365 175.175 46.075 ;
      RECT 167.985 44.365 173.33 46.075 ;
      RECT 162.465 44.365 167.81 46.075 ;
      RECT 158.785 44.365 160.455 46.075 ;
      RECT 153.265 44.365 158.61 46.075 ;
      RECT 147.745 44.365 153.09 46.075 ;
      RECT 144.065 44.365 145.735 46.075 ;
      RECT 138.545 44.365 143.89 46.075 ;
      RECT 133.025 44.365 138.37 46.075 ;
      RECT 129.345 44.365 131.015 46.075 ;
      RECT 123.825 44.365 129.17 46.075 ;
      RECT 118.305 44.365 123.65 46.075 ;
      RECT 114.625 44.365 116.295 46.075 ;
      RECT 109.105 44.365 114.45 46.075 ;
      RECT 103.585 44.365 108.93 46.075 ;
      RECT 99.905 44.365 101.575 46.075 ;
      RECT 94.385 44.365 99.73 46.075 ;
      RECT 88.865 44.365 94.21 46.075 ;
      RECT 85.185 44.365 86.855 46.075 ;
      RECT 79.665 44.365 85.01 46.075 ;
      RECT 74.145 44.365 79.49 46.075 ;
      RECT 70.465 44.365 72.135 46.075 ;
      RECT 64.945 44.365 70.29 46.075 ;
      RECT 59.425 44.365 64.77 46.075 ;
      RECT 55.745 44.365 57.415 46.075 ;
      RECT 50.225 44.365 55.57 46.075 ;
      RECT 44.705 44.365 50.05 46.075 ;
      RECT 41.025 44.365 42.695 46.075 ;
      RECT 35.505 44.365 40.85 46.075 ;
      RECT 29.985 44.365 35.33 46.075 ;
      RECT 26.305 44.365 27.975 46.075 ;
      RECT 20.785 44.365 26.13 46.075 ;
      RECT 15.265 44.365 20.61 46.075 ;
      RECT 10.665 44.365 13.255 46.075 ;
      RECT 175.345 44.385 176.555 46.055 ;
      RECT 160.625 44.385 161.835 46.055 ;
      RECT 145.905 44.385 147.115 46.055 ;
      RECT 131.185 44.385 132.395 46.055 ;
      RECT 116.465 44.385 117.675 46.055 ;
      RECT 101.745 44.385 102.955 46.055 ;
      RECT 87.025 44.385 88.235 46.055 ;
      RECT 72.305 44.385 73.515 46.055 ;
      RECT 57.585 44.385 58.795 46.055 ;
      RECT 42.865 44.385 44.075 46.055 ;
      RECT 28.145 44.385 29.355 46.055 ;
      RECT 13.425 44.385 14.635 46.055 ;
      RECT 189.605 44.41 189.895 46.03 ;
      RECT 189.145 44.41 189.435 46.03 ;
      RECT 176.725 44.41 177.015 46.03 ;
      RECT 162.005 44.41 162.295 46.03 ;
      RECT 147.285 44.41 147.575 46.03 ;
      RECT 132.565 44.41 132.855 46.03 ;
      RECT 117.845 44.41 118.135 46.03 ;
      RECT 103.125 44.41 103.415 46.03 ;
      RECT 88.405 44.41 88.695 46.03 ;
      RECT 73.685 44.41 73.975 46.03 ;
      RECT 58.965 44.41 59.255 46.03 ;
      RECT 44.245 44.41 44.535 46.03 ;
      RECT 29.525 44.41 29.815 46.03 ;
      RECT 14.805 44.41 15.095 46.03 ;
      RECT 10.205 44.41 10.495 46.03 ;
      RECT 10.12 45.135 189.98 45.305 ;
      RECT 176.035 46.225 176.555 49.655 ;
      RECT 161.315 46.225 161.835 49.655 ;
      RECT 146.595 46.225 147.115 49.655 ;
      RECT 131.875 46.225 132.395 49.655 ;
      RECT 117.155 46.225 117.675 49.655 ;
      RECT 102.435 46.225 102.955 49.655 ;
      RECT 87.715 46.225 88.235 49.655 ;
      RECT 72.995 46.225 73.515 49.655 ;
      RECT 58.275 46.225 58.795 49.655 ;
      RECT 43.555 46.225 44.075 49.655 ;
      RECT 28.835 46.225 29.355 49.655 ;
      RECT 14.115 46.225 14.635 49.655 ;
      RECT 187.765 46.245 188.975 49.635 ;
      RECT 184.525 46.245 186.215 49.635 ;
      RECT 179.935 46.245 182.53 49.635 ;
      RECT 174.425 46.245 175.175 49.635 ;
      RECT 170.735 46.245 173.33 49.635 ;
      RECT 165.215 46.245 167.81 49.635 ;
      RECT 159.705 46.245 160.455 49.635 ;
      RECT 156.015 46.245 158.61 49.635 ;
      RECT 150.495 46.245 153.09 49.635 ;
      RECT 144.985 46.245 145.735 49.635 ;
      RECT 141.295 46.245 143.89 49.635 ;
      RECT 135.775 46.245 138.37 49.635 ;
      RECT 130.265 46.245 131.015 49.635 ;
      RECT 126.575 46.245 129.17 49.635 ;
      RECT 121.055 46.245 123.65 49.635 ;
      RECT 115.545 46.245 116.295 49.635 ;
      RECT 111.855 46.245 114.45 49.635 ;
      RECT 106.335 46.245 108.93 49.635 ;
      RECT 100.825 46.245 101.575 49.635 ;
      RECT 97.135 46.245 99.73 49.635 ;
      RECT 91.615 46.245 94.21 49.635 ;
      RECT 86.105 46.245 86.855 49.635 ;
      RECT 82.415 46.245 85.01 49.635 ;
      RECT 76.895 46.245 79.49 49.635 ;
      RECT 71.385 46.245 72.135 49.635 ;
      RECT 67.695 46.245 70.29 49.635 ;
      RECT 62.175 46.245 64.77 49.635 ;
      RECT 56.665 46.245 57.415 49.635 ;
      RECT 52.975 46.245 55.57 49.635 ;
      RECT 47.455 46.245 50.05 49.635 ;
      RECT 41.945 46.245 42.695 49.635 ;
      RECT 38.255 46.245 40.85 49.635 ;
      RECT 32.735 46.245 35.33 49.635 ;
      RECT 27.225 46.245 27.975 49.635 ;
      RECT 23.535 46.245 26.13 49.635 ;
      RECT 18.015 46.245 20.61 49.635 ;
      RECT 12.045 46.245 13.255 49.635 ;
      RECT 189.605 46.69 189.895 49.19 ;
      RECT 189.145 46.69 189.435 49.19 ;
      RECT 176.725 46.69 177.015 49.19 ;
      RECT 162.005 46.69 162.295 49.19 ;
      RECT 147.285 46.69 147.575 49.19 ;
      RECT 132.565 46.69 132.855 49.19 ;
      RECT 117.845 46.69 118.135 49.19 ;
      RECT 103.125 46.69 103.415 49.19 ;
      RECT 88.405 46.69 88.695 49.19 ;
      RECT 73.685 46.69 73.975 49.19 ;
      RECT 58.965 46.69 59.255 49.19 ;
      RECT 44.245 46.69 44.535 49.19 ;
      RECT 29.525 46.69 29.815 49.19 ;
      RECT 14.805 46.69 15.095 49.19 ;
      RECT 10.205 46.69 10.495 49.19 ;
      RECT 186.385 46.765 188.975 49.115 ;
      RECT 182.705 46.765 186.215 49.115 ;
      RECT 177.185 46.765 182.53 49.115 ;
      RECT 175.345 46.765 176.555 49.115 ;
      RECT 173.505 46.765 175.175 49.115 ;
      RECT 167.985 46.765 173.33 49.115 ;
      RECT 162.465 46.765 167.81 49.115 ;
      RECT 160.625 46.765 161.835 49.115 ;
      RECT 158.785 46.765 160.455 49.115 ;
      RECT 153.265 46.765 158.61 49.115 ;
      RECT 147.745 46.765 153.09 49.115 ;
      RECT 145.905 46.765 147.115 49.115 ;
      RECT 144.065 46.765 145.735 49.115 ;
      RECT 138.545 46.765 143.89 49.115 ;
      RECT 133.025 46.765 138.37 49.115 ;
      RECT 131.185 46.765 132.395 49.115 ;
      RECT 129.345 46.765 131.015 49.115 ;
      RECT 123.825 46.765 129.17 49.115 ;
      RECT 118.305 46.765 123.65 49.115 ;
      RECT 116.465 46.765 117.675 49.115 ;
      RECT 114.625 46.765 116.295 49.115 ;
      RECT 109.105 46.765 114.45 49.115 ;
      RECT 103.585 46.765 108.93 49.115 ;
      RECT 101.745 46.765 102.955 49.115 ;
      RECT 99.905 46.765 101.575 49.115 ;
      RECT 94.385 46.765 99.73 49.115 ;
      RECT 88.865 46.765 94.21 49.115 ;
      RECT 87.025 46.765 88.235 49.115 ;
      RECT 85.185 46.765 86.855 49.115 ;
      RECT 79.665 46.765 85.01 49.115 ;
      RECT 74.145 46.765 79.49 49.115 ;
      RECT 72.305 46.765 73.515 49.115 ;
      RECT 70.465 46.765 72.135 49.115 ;
      RECT 64.945 46.765 70.29 49.115 ;
      RECT 59.425 46.765 64.77 49.115 ;
      RECT 57.585 46.765 58.795 49.115 ;
      RECT 55.745 46.765 57.415 49.115 ;
      RECT 50.225 46.765 55.57 49.115 ;
      RECT 44.705 46.765 50.05 49.115 ;
      RECT 42.865 46.765 44.075 49.115 ;
      RECT 41.025 46.765 42.695 49.115 ;
      RECT 35.505 46.765 40.85 49.115 ;
      RECT 29.985 46.765 35.33 49.115 ;
      RECT 28.145 46.765 29.355 49.115 ;
      RECT 26.305 46.765 27.975 49.115 ;
      RECT 20.785 46.765 26.13 49.115 ;
      RECT 15.265 46.765 20.61 49.115 ;
      RECT 13.425 46.765 14.635 49.115 ;
      RECT 10.665 46.765 13.255 49.115 ;
      RECT 10.12 47.855 189.98 48.025 ;
      RECT 186.385 49.285 187.595 52.035 ;
      RECT 182.705 49.285 184.355 52.035 ;
      RECT 177.185 49.285 179.765 52.035 ;
      RECT 175.345 49.285 175.865 52.035 ;
      RECT 173.505 49.285 174.255 52.035 ;
      RECT 167.985 49.285 170.565 52.035 ;
      RECT 162.465 49.285 165.045 52.035 ;
      RECT 160.625 49.285 161.145 52.035 ;
      RECT 158.785 49.285 159.535 52.035 ;
      RECT 153.265 49.285 155.845 52.035 ;
      RECT 147.745 49.285 150.325 52.035 ;
      RECT 145.905 49.285 146.425 52.035 ;
      RECT 144.065 49.285 144.815 52.035 ;
      RECT 138.545 49.285 141.125 52.035 ;
      RECT 133.025 49.285 135.605 52.035 ;
      RECT 131.185 49.285 131.705 52.035 ;
      RECT 129.345 49.285 130.095 52.035 ;
      RECT 123.825 49.285 126.405 52.035 ;
      RECT 118.305 49.285 120.885 52.035 ;
      RECT 116.465 49.285 116.985 52.035 ;
      RECT 114.625 49.285 115.375 52.035 ;
      RECT 109.105 49.285 111.685 52.035 ;
      RECT 103.585 49.285 106.165 52.035 ;
      RECT 101.745 49.285 102.265 52.035 ;
      RECT 99.905 49.285 100.655 52.035 ;
      RECT 94.385 49.285 96.965 52.035 ;
      RECT 88.865 49.285 91.445 52.035 ;
      RECT 87.025 49.285 87.545 52.035 ;
      RECT 85.185 49.285 85.935 52.035 ;
      RECT 79.665 49.285 82.245 52.035 ;
      RECT 74.145 49.285 76.725 52.035 ;
      RECT 72.305 49.285 72.825 52.035 ;
      RECT 70.465 49.285 71.215 52.035 ;
      RECT 64.945 49.285 67.525 52.035 ;
      RECT 59.425 49.285 62.005 52.035 ;
      RECT 57.585 49.285 58.105 52.035 ;
      RECT 55.745 49.285 56.495 52.035 ;
      RECT 50.225 49.285 52.805 52.035 ;
      RECT 44.705 49.285 47.285 52.035 ;
      RECT 42.865 49.285 43.385 52.035 ;
      RECT 41.025 49.285 41.775 52.035 ;
      RECT 35.505 49.285 38.085 52.035 ;
      RECT 29.985 49.285 32.565 52.035 ;
      RECT 28.145 49.285 28.665 52.035 ;
      RECT 26.305 49.285 27.055 52.035 ;
      RECT 20.785 49.285 23.365 52.035 ;
      RECT 15.265 49.285 17.845 52.035 ;
      RECT 13.425 49.285 13.945 52.035 ;
      RECT 10.665 49.285 11.875 52.035 ;
      RECT 186.385 49.805 188.975 51.515 ;
      RECT 182.705 49.805 186.215 51.515 ;
      RECT 177.185 49.805 182.53 51.515 ;
      RECT 173.505 49.805 175.175 51.515 ;
      RECT 167.985 49.805 173.33 51.515 ;
      RECT 162.465 49.805 167.81 51.515 ;
      RECT 158.785 49.805 160.455 51.515 ;
      RECT 153.265 49.805 158.61 51.515 ;
      RECT 147.745 49.805 153.09 51.515 ;
      RECT 144.065 49.805 145.735 51.515 ;
      RECT 138.545 49.805 143.89 51.515 ;
      RECT 133.025 49.805 138.37 51.515 ;
      RECT 129.345 49.805 131.015 51.515 ;
      RECT 123.825 49.805 129.17 51.515 ;
      RECT 118.305 49.805 123.65 51.515 ;
      RECT 114.625 49.805 116.295 51.515 ;
      RECT 109.105 49.805 114.45 51.515 ;
      RECT 103.585 49.805 108.93 51.515 ;
      RECT 99.905 49.805 101.575 51.515 ;
      RECT 94.385 49.805 99.73 51.515 ;
      RECT 88.865 49.805 94.21 51.515 ;
      RECT 85.185 49.805 86.855 51.515 ;
      RECT 79.665 49.805 85.01 51.515 ;
      RECT 74.145 49.805 79.49 51.515 ;
      RECT 70.465 49.805 72.135 51.515 ;
      RECT 64.945 49.805 70.29 51.515 ;
      RECT 59.425 49.805 64.77 51.515 ;
      RECT 55.745 49.805 57.415 51.515 ;
      RECT 50.225 49.805 55.57 51.515 ;
      RECT 44.705 49.805 50.05 51.515 ;
      RECT 41.025 49.805 42.695 51.515 ;
      RECT 35.505 49.805 40.85 51.515 ;
      RECT 29.985 49.805 35.33 51.515 ;
      RECT 26.305 49.805 27.975 51.515 ;
      RECT 20.785 49.805 26.13 51.515 ;
      RECT 15.265 49.805 20.61 51.515 ;
      RECT 10.665 49.805 13.255 51.515 ;
      RECT 175.345 49.825 176.555 51.495 ;
      RECT 160.625 49.825 161.835 51.495 ;
      RECT 145.905 49.825 147.115 51.495 ;
      RECT 131.185 49.825 132.395 51.495 ;
      RECT 116.465 49.825 117.675 51.495 ;
      RECT 101.745 49.825 102.955 51.495 ;
      RECT 87.025 49.825 88.235 51.495 ;
      RECT 72.305 49.825 73.515 51.495 ;
      RECT 57.585 49.825 58.795 51.495 ;
      RECT 42.865 49.825 44.075 51.495 ;
      RECT 28.145 49.825 29.355 51.495 ;
      RECT 13.425 49.825 14.635 51.495 ;
      RECT 189.605 49.85 189.895 51.47 ;
      RECT 189.145 49.85 189.435 51.47 ;
      RECT 176.725 49.85 177.015 51.47 ;
      RECT 162.005 49.85 162.295 51.47 ;
      RECT 147.285 49.85 147.575 51.47 ;
      RECT 132.565 49.85 132.855 51.47 ;
      RECT 117.845 49.85 118.135 51.47 ;
      RECT 103.125 49.85 103.415 51.47 ;
      RECT 88.405 49.85 88.695 51.47 ;
      RECT 73.685 49.85 73.975 51.47 ;
      RECT 58.965 49.85 59.255 51.47 ;
      RECT 44.245 49.85 44.535 51.47 ;
      RECT 29.525 49.85 29.815 51.47 ;
      RECT 14.805 49.85 15.095 51.47 ;
      RECT 10.205 49.85 10.495 51.47 ;
      RECT 10.12 50.575 189.98 50.745 ;
      RECT 176.035 51.665 176.555 55.095 ;
      RECT 161.315 51.665 161.835 55.095 ;
      RECT 146.595 51.665 147.115 55.095 ;
      RECT 131.875 51.665 132.395 55.095 ;
      RECT 117.155 51.665 117.675 55.095 ;
      RECT 102.435 51.665 102.955 55.095 ;
      RECT 87.715 51.665 88.235 55.095 ;
      RECT 72.995 51.665 73.515 55.095 ;
      RECT 58.275 51.665 58.795 55.095 ;
      RECT 43.555 51.665 44.075 55.095 ;
      RECT 28.835 51.665 29.355 55.095 ;
      RECT 14.115 51.665 14.635 55.095 ;
      RECT 187.765 51.685 188.975 55.075 ;
      RECT 184.525 51.685 186.215 55.075 ;
      RECT 179.935 51.685 182.53 55.075 ;
      RECT 174.425 51.685 175.175 55.075 ;
      RECT 170.735 51.685 173.33 55.075 ;
      RECT 165.215 51.685 167.81 55.075 ;
      RECT 159.705 51.685 160.455 55.075 ;
      RECT 156.015 51.685 158.61 55.075 ;
      RECT 150.495 51.685 153.09 55.075 ;
      RECT 144.985 51.685 145.735 55.075 ;
      RECT 141.295 51.685 143.89 55.075 ;
      RECT 135.775 51.685 138.37 55.075 ;
      RECT 130.265 51.685 131.015 55.075 ;
      RECT 126.575 51.685 129.17 55.075 ;
      RECT 121.055 51.685 123.65 55.075 ;
      RECT 115.545 51.685 116.295 55.075 ;
      RECT 111.855 51.685 114.45 55.075 ;
      RECT 106.335 51.685 108.93 55.075 ;
      RECT 100.825 51.685 101.575 55.075 ;
      RECT 97.135 51.685 99.73 55.075 ;
      RECT 91.615 51.685 94.21 55.075 ;
      RECT 86.105 51.685 86.855 55.075 ;
      RECT 82.415 51.685 85.01 55.075 ;
      RECT 76.895 51.685 79.49 55.075 ;
      RECT 71.385 51.685 72.135 55.075 ;
      RECT 67.695 51.685 70.29 55.075 ;
      RECT 62.175 51.685 64.77 55.075 ;
      RECT 56.665 51.685 57.415 55.075 ;
      RECT 52.975 51.685 55.57 55.075 ;
      RECT 47.455 51.685 50.05 55.075 ;
      RECT 41.945 51.685 42.695 55.075 ;
      RECT 38.255 51.685 40.85 55.075 ;
      RECT 32.735 51.685 35.33 55.075 ;
      RECT 27.225 51.685 27.975 55.075 ;
      RECT 23.535 51.685 26.13 55.075 ;
      RECT 18.015 51.685 20.61 55.075 ;
      RECT 12.045 51.685 13.255 55.075 ;
      RECT 189.605 52.13 189.895 54.63 ;
      RECT 189.145 52.13 189.435 54.63 ;
      RECT 176.725 52.13 177.015 54.63 ;
      RECT 162.005 52.13 162.295 54.63 ;
      RECT 147.285 52.13 147.575 54.63 ;
      RECT 132.565 52.13 132.855 54.63 ;
      RECT 117.845 52.13 118.135 54.63 ;
      RECT 103.125 52.13 103.415 54.63 ;
      RECT 88.405 52.13 88.695 54.63 ;
      RECT 73.685 52.13 73.975 54.63 ;
      RECT 58.965 52.13 59.255 54.63 ;
      RECT 44.245 52.13 44.535 54.63 ;
      RECT 29.525 52.13 29.815 54.63 ;
      RECT 14.805 52.13 15.095 54.63 ;
      RECT 10.205 52.13 10.495 54.63 ;
      RECT 186.385 52.205 188.975 54.555 ;
      RECT 182.705 52.205 186.215 54.555 ;
      RECT 177.185 52.205 182.53 54.555 ;
      RECT 175.345 52.205 176.555 54.555 ;
      RECT 173.505 52.205 175.175 54.555 ;
      RECT 167.985 52.205 173.33 54.555 ;
      RECT 162.465 52.205 167.81 54.555 ;
      RECT 160.625 52.205 161.835 54.555 ;
      RECT 158.785 52.205 160.455 54.555 ;
      RECT 153.265 52.205 158.61 54.555 ;
      RECT 147.745 52.205 153.09 54.555 ;
      RECT 145.905 52.205 147.115 54.555 ;
      RECT 144.065 52.205 145.735 54.555 ;
      RECT 138.545 52.205 143.89 54.555 ;
      RECT 133.025 52.205 138.37 54.555 ;
      RECT 131.185 52.205 132.395 54.555 ;
      RECT 129.345 52.205 131.015 54.555 ;
      RECT 123.825 52.205 129.17 54.555 ;
      RECT 118.305 52.205 123.65 54.555 ;
      RECT 116.465 52.205 117.675 54.555 ;
      RECT 114.625 52.205 116.295 54.555 ;
      RECT 109.105 52.205 114.45 54.555 ;
      RECT 103.585 52.205 108.93 54.555 ;
      RECT 101.745 52.205 102.955 54.555 ;
      RECT 99.905 52.205 101.575 54.555 ;
      RECT 94.385 52.205 99.73 54.555 ;
      RECT 88.865 52.205 94.21 54.555 ;
      RECT 87.025 52.205 88.235 54.555 ;
      RECT 85.185 52.205 86.855 54.555 ;
      RECT 79.665 52.205 85.01 54.555 ;
      RECT 74.145 52.205 79.49 54.555 ;
      RECT 72.305 52.205 73.515 54.555 ;
      RECT 70.465 52.205 72.135 54.555 ;
      RECT 64.945 52.205 70.29 54.555 ;
      RECT 59.425 52.205 64.77 54.555 ;
      RECT 57.585 52.205 58.795 54.555 ;
      RECT 55.745 52.205 57.415 54.555 ;
      RECT 50.225 52.205 55.57 54.555 ;
      RECT 44.705 52.205 50.05 54.555 ;
      RECT 42.865 52.205 44.075 54.555 ;
      RECT 41.025 52.205 42.695 54.555 ;
      RECT 35.505 52.205 40.85 54.555 ;
      RECT 29.985 52.205 35.33 54.555 ;
      RECT 28.145 52.205 29.355 54.555 ;
      RECT 26.305 52.205 27.975 54.555 ;
      RECT 20.785 52.205 26.13 54.555 ;
      RECT 15.265 52.205 20.61 54.555 ;
      RECT 13.425 52.205 14.635 54.555 ;
      RECT 10.665 52.205 13.255 54.555 ;
      RECT 10.12 53.295 189.98 53.465 ;
      RECT 186.385 54.725 187.595 57.475 ;
      RECT 182.705 54.725 184.355 57.475 ;
      RECT 177.185 54.725 179.765 57.475 ;
      RECT 175.345 54.725 175.865 57.475 ;
      RECT 173.505 54.725 174.255 57.475 ;
      RECT 167.985 54.725 170.565 57.475 ;
      RECT 162.465 54.725 165.045 57.475 ;
      RECT 160.625 54.725 161.145 57.475 ;
      RECT 158.785 54.725 159.535 57.475 ;
      RECT 153.265 54.725 155.845 57.475 ;
      RECT 147.745 54.725 150.325 57.475 ;
      RECT 145.905 54.725 146.425 57.475 ;
      RECT 144.065 54.725 144.815 57.475 ;
      RECT 138.545 54.725 141.125 57.475 ;
      RECT 133.025 54.725 135.605 57.475 ;
      RECT 131.185 54.725 131.705 57.475 ;
      RECT 129.345 54.725 130.095 57.475 ;
      RECT 123.825 54.725 126.405 57.475 ;
      RECT 118.305 54.725 120.885 57.475 ;
      RECT 116.465 54.725 116.985 57.475 ;
      RECT 114.625 54.725 115.375 57.475 ;
      RECT 109.105 54.725 111.685 57.475 ;
      RECT 103.585 54.725 106.165 57.475 ;
      RECT 101.745 54.725 102.265 57.475 ;
      RECT 99.905 54.725 100.655 57.475 ;
      RECT 94.385 54.725 96.965 57.475 ;
      RECT 88.865 54.725 91.445 57.475 ;
      RECT 87.025 54.725 87.545 57.475 ;
      RECT 85.185 54.725 85.935 57.475 ;
      RECT 79.665 54.725 82.245 57.475 ;
      RECT 74.145 54.725 76.725 57.475 ;
      RECT 72.305 54.725 72.825 57.475 ;
      RECT 70.465 54.725 71.215 57.475 ;
      RECT 64.945 54.725 67.525 57.475 ;
      RECT 59.425 54.725 62.005 57.475 ;
      RECT 57.585 54.725 58.105 57.475 ;
      RECT 55.745 54.725 56.495 57.475 ;
      RECT 50.225 54.725 52.805 57.475 ;
      RECT 44.705 54.725 47.285 57.475 ;
      RECT 42.865 54.725 43.385 57.475 ;
      RECT 41.025 54.725 41.775 57.475 ;
      RECT 35.505 54.725 38.085 57.475 ;
      RECT 29.985 54.725 32.565 57.475 ;
      RECT 28.145 54.725 28.665 57.475 ;
      RECT 26.305 54.725 27.055 57.475 ;
      RECT 20.785 54.725 23.365 57.475 ;
      RECT 15.265 54.725 17.845 57.475 ;
      RECT 13.425 54.725 13.945 57.475 ;
      RECT 10.665 54.725 11.875 57.475 ;
      RECT 186.385 55.245 188.975 56.955 ;
      RECT 182.705 55.245 186.215 56.955 ;
      RECT 177.185 55.245 182.53 56.955 ;
      RECT 173.505 55.245 175.175 56.955 ;
      RECT 167.985 55.245 173.33 56.955 ;
      RECT 162.465 55.245 167.81 56.955 ;
      RECT 158.785 55.245 160.455 56.955 ;
      RECT 153.265 55.245 158.61 56.955 ;
      RECT 147.745 55.245 153.09 56.955 ;
      RECT 144.065 55.245 145.735 56.955 ;
      RECT 138.545 55.245 143.89 56.955 ;
      RECT 133.025 55.245 138.37 56.955 ;
      RECT 129.345 55.245 131.015 56.955 ;
      RECT 123.825 55.245 129.17 56.955 ;
      RECT 118.305 55.245 123.65 56.955 ;
      RECT 114.625 55.245 116.295 56.955 ;
      RECT 109.105 55.245 114.45 56.955 ;
      RECT 103.585 55.245 108.93 56.955 ;
      RECT 99.905 55.245 101.575 56.955 ;
      RECT 94.385 55.245 99.73 56.955 ;
      RECT 88.865 55.245 94.21 56.955 ;
      RECT 85.185 55.245 86.855 56.955 ;
      RECT 79.665 55.245 85.01 56.955 ;
      RECT 74.145 55.245 79.49 56.955 ;
      RECT 70.465 55.245 72.135 56.955 ;
      RECT 64.945 55.245 70.29 56.955 ;
      RECT 59.425 55.245 64.77 56.955 ;
      RECT 55.745 55.245 57.415 56.955 ;
      RECT 50.225 55.245 55.57 56.955 ;
      RECT 44.705 55.245 50.05 56.955 ;
      RECT 41.025 55.245 42.695 56.955 ;
      RECT 35.505 55.245 40.85 56.955 ;
      RECT 29.985 55.245 35.33 56.955 ;
      RECT 26.305 55.245 27.975 56.955 ;
      RECT 20.785 55.245 26.13 56.955 ;
      RECT 15.265 55.245 20.61 56.955 ;
      RECT 10.665 55.245 13.255 56.955 ;
      RECT 175.345 55.265 176.555 56.935 ;
      RECT 160.625 55.265 161.835 56.935 ;
      RECT 145.905 55.265 147.115 56.935 ;
      RECT 131.185 55.265 132.395 56.935 ;
      RECT 116.465 55.265 117.675 56.935 ;
      RECT 101.745 55.265 102.955 56.935 ;
      RECT 87.025 55.265 88.235 56.935 ;
      RECT 72.305 55.265 73.515 56.935 ;
      RECT 57.585 55.265 58.795 56.935 ;
      RECT 42.865 55.265 44.075 56.935 ;
      RECT 28.145 55.265 29.355 56.935 ;
      RECT 13.425 55.265 14.635 56.935 ;
      RECT 189.605 55.29 189.895 56.91 ;
      RECT 189.145 55.29 189.435 56.91 ;
      RECT 176.725 55.29 177.015 56.91 ;
      RECT 162.005 55.29 162.295 56.91 ;
      RECT 147.285 55.29 147.575 56.91 ;
      RECT 132.565 55.29 132.855 56.91 ;
      RECT 117.845 55.29 118.135 56.91 ;
      RECT 103.125 55.29 103.415 56.91 ;
      RECT 88.405 55.29 88.695 56.91 ;
      RECT 73.685 55.29 73.975 56.91 ;
      RECT 58.965 55.29 59.255 56.91 ;
      RECT 44.245 55.29 44.535 56.91 ;
      RECT 29.525 55.29 29.815 56.91 ;
      RECT 14.805 55.29 15.095 56.91 ;
      RECT 10.205 55.29 10.495 56.91 ;
      RECT 10.12 56.015 189.98 56.185 ;
      RECT 10.12 58.735 189.98 58.905 ;
      RECT 189.605 57.57 189.895 58.905 ;
      RECT 189.145 57.57 189.435 58.905 ;
      RECT 186.385 57.645 188.975 58.905 ;
      RECT 187.765 57.125 188.975 58.905 ;
      RECT 182.705 57.645 186.215 58.905 ;
      RECT 184.525 57.125 186.215 58.905 ;
      RECT 177.185 57.645 182.53 58.905 ;
      RECT 179.935 57.125 182.53 58.905 ;
      RECT 176.725 57.57 177.015 58.905 ;
      RECT 175.345 57.645 176.555 58.905 ;
      RECT 176.035 57.105 176.555 58.905 ;
      RECT 173.505 57.645 175.175 58.905 ;
      RECT 174.425 57.125 175.175 58.905 ;
      RECT 167.985 57.645 173.33 58.905 ;
      RECT 170.735 57.125 173.33 58.905 ;
      RECT 162.465 57.645 167.81 58.905 ;
      RECT 165.215 57.125 167.81 58.905 ;
      RECT 162.005 57.57 162.295 58.905 ;
      RECT 160.625 57.645 161.835 58.905 ;
      RECT 161.315 57.105 161.835 58.905 ;
      RECT 158.785 57.645 160.455 58.905 ;
      RECT 159.705 57.125 160.455 58.905 ;
      RECT 153.265 57.645 158.61 58.905 ;
      RECT 156.015 57.125 158.61 58.905 ;
      RECT 147.745 57.645 153.09 58.905 ;
      RECT 150.495 57.125 153.09 58.905 ;
      RECT 147.285 57.57 147.575 58.905 ;
      RECT 145.905 57.645 147.115 58.905 ;
      RECT 146.595 57.105 147.115 58.905 ;
      RECT 144.065 57.645 145.735 58.905 ;
      RECT 144.985 57.125 145.735 58.905 ;
      RECT 138.545 57.645 143.89 58.905 ;
      RECT 141.295 57.125 143.89 58.905 ;
      RECT 133.025 57.645 138.37 58.905 ;
      RECT 135.775 57.125 138.37 58.905 ;
      RECT 132.565 57.57 132.855 58.905 ;
      RECT 131.185 57.645 132.395 58.905 ;
      RECT 131.875 57.105 132.395 58.905 ;
      RECT 129.345 57.645 131.015 58.905 ;
      RECT 130.265 57.125 131.015 58.905 ;
      RECT 123.825 57.645 129.17 58.905 ;
      RECT 126.575 57.125 129.17 58.905 ;
      RECT 118.305 57.645 123.65 58.905 ;
      RECT 121.055 57.125 123.65 58.905 ;
      RECT 117.845 57.57 118.135 58.905 ;
      RECT 116.465 57.645 117.675 58.905 ;
      RECT 117.155 57.105 117.675 58.905 ;
      RECT 114.625 57.645 116.295 58.905 ;
      RECT 115.545 57.125 116.295 58.905 ;
      RECT 109.105 57.645 114.45 58.905 ;
      RECT 111.855 57.125 114.45 58.905 ;
      RECT 103.585 57.645 108.93 58.905 ;
      RECT 106.335 57.125 108.93 58.905 ;
      RECT 103.125 57.57 103.415 58.905 ;
      RECT 101.745 57.645 102.955 58.905 ;
      RECT 102.435 57.105 102.955 58.905 ;
      RECT 99.905 57.645 101.575 58.905 ;
      RECT 100.825 57.125 101.575 58.905 ;
      RECT 94.385 57.645 99.73 58.905 ;
      RECT 97.135 57.125 99.73 58.905 ;
      RECT 88.865 57.645 94.21 58.905 ;
      RECT 91.615 57.125 94.21 58.905 ;
      RECT 88.405 57.57 88.695 58.905 ;
      RECT 87.025 57.645 88.235 58.905 ;
      RECT 87.715 57.105 88.235 58.905 ;
      RECT 85.185 57.645 86.855 58.905 ;
      RECT 86.105 57.125 86.855 58.905 ;
      RECT 79.665 57.645 85.01 58.905 ;
      RECT 82.415 57.125 85.01 58.905 ;
      RECT 74.145 57.645 79.49 58.905 ;
      RECT 76.895 57.125 79.49 58.905 ;
      RECT 73.685 57.57 73.975 58.905 ;
      RECT 72.305 57.645 73.515 58.905 ;
      RECT 72.995 57.105 73.515 58.905 ;
      RECT 70.465 57.645 72.135 58.905 ;
      RECT 71.385 57.125 72.135 58.905 ;
      RECT 64.945 57.645 70.29 58.905 ;
      RECT 67.695 57.125 70.29 58.905 ;
      RECT 59.425 57.645 64.77 58.905 ;
      RECT 62.175 57.125 64.77 58.905 ;
      RECT 58.965 57.57 59.255 58.905 ;
      RECT 57.585 57.645 58.795 58.905 ;
      RECT 58.275 57.105 58.795 58.905 ;
      RECT 55.745 57.645 57.415 58.905 ;
      RECT 56.665 57.125 57.415 58.905 ;
      RECT 50.225 57.645 55.57 58.905 ;
      RECT 52.975 57.125 55.57 58.905 ;
      RECT 44.705 57.645 50.05 58.905 ;
      RECT 47.455 57.125 50.05 58.905 ;
      RECT 44.245 57.57 44.535 58.905 ;
      RECT 42.865 57.645 44.075 58.905 ;
      RECT 43.555 57.105 44.075 58.905 ;
      RECT 41.025 57.645 42.695 58.905 ;
      RECT 41.945 57.125 42.695 58.905 ;
      RECT 35.505 57.645 40.85 58.905 ;
      RECT 38.255 57.125 40.85 58.905 ;
      RECT 29.985 57.645 35.33 58.905 ;
      RECT 32.735 57.125 35.33 58.905 ;
      RECT 29.525 57.57 29.815 58.905 ;
      RECT 28.145 57.645 29.355 58.905 ;
      RECT 28.835 57.105 29.355 58.905 ;
      RECT 26.305 57.645 27.975 58.905 ;
      RECT 27.225 57.125 27.975 58.905 ;
      RECT 20.785 57.645 26.13 58.905 ;
      RECT 23.535 57.125 26.13 58.905 ;
      RECT 15.265 57.645 20.61 58.905 ;
      RECT 18.015 57.125 20.61 58.905 ;
      RECT 14.805 57.57 15.095 58.905 ;
      RECT 13.425 57.645 14.635 58.905 ;
      RECT 14.115 57.105 14.635 58.905 ;
      RECT 10.665 57.645 13.255 58.905 ;
      RECT 12.045 57.125 13.255 58.905 ;
      RECT 10.205 57.57 10.495 58.905 ;
      RECT 183.995 17.195 184.325 17.715 ;
      RECT 184.205 16.445 184.375 17.28 ;
      RECT 184.15 17.155 184.375 17.28 ;
      RECT 184.16 16.445 184.375 16.575 ;
      RECT 183.985 15.6 184.315 16.525 ;
      RECT 183.155 17.195 183.485 17.72 ;
      RECT 183.285 16.695 183.485 17.72 ;
      RECT 183.285 16.695 184.035 17.025 ;
      RECT 183.285 15.555 183.475 17.72 ;
      RECT 182.58 16.115 183.475 16.49 ;
      RECT 183.135 15.555 183.475 16.49 ;
      RECT 183.655 11.82 183.915 12.325 ;
      RECT 183.735 10.115 183.915 12.325 ;
      RECT 183.645 10.115 183.915 11.02 ;
      RECT 182.795 11.775 182.965 12.325 ;
      RECT 182.795 11.775 183.46 11.945 ;
      RECT 183.29 10.875 183.46 11.945 ;
      RECT 183.29 11.19 183.565 11.52 ;
      RECT 182.785 10.875 183.46 11.045 ;
      RECT 182.785 10.115 182.965 11.045 ;
      RECT 181.625 17.485 182.41 17.655 ;
      RECT 182.24 15.685 182.41 17.655 ;
      RECT 182.24 16.695 183.115 17.025 ;
      RECT 181.525 15.685 182.41 15.855 ;
      RECT 181.605 16.985 182.07 17.315 ;
      RECT 181.75 16.025 182.07 17.315 ;
      RECT 181.05 17.485 181.455 17.655 ;
      RECT 181.05 15.555 181.22 17.655 ;
      RECT 180.39 16.955 181.22 17.255 ;
      RECT 180.39 16.925 180.59 17.255 ;
      RECT 181.05 15.555 181.3 15.885 ;
      RECT 177.275 11.675 177.445 12.325 ;
      RECT 178.115 11.675 178.285 12.32 ;
      RECT 177.275 11.675 178.695 11.845 ;
      RECT 178.52 10.965 178.695 11.845 ;
      RECT 178.52 11.335 181.145 11.505 ;
      RECT 177.195 10.965 178.695 11.135 ;
      RECT 178.035 10.115 178.365 11.135 ;
      RECT 177.195 10.115 177.525 11.135 ;
      RECT 179.505 17.485 180.18 17.655 ;
      RECT 180.01 16.535 180.18 17.655 ;
      RECT 180.71 16.445 180.88 16.775 ;
      RECT 180.01 16.535 180.88 16.705 ;
      RECT 180.37 16.445 180.88 16.705 ;
      RECT 180.37 15.66 180.54 16.705 ;
      RECT 179.435 15.66 180.54 15.83 ;
      RECT 179.315 17.065 179.84 17.285 ;
      RECT 179.67 16 179.84 17.285 ;
      RECT 179.67 16 180.2 16.365 ;
      RECT 178.975 17.485 179.31 17.655 ;
      RECT 178.975 17.215 179.145 17.655 ;
      RECT 178.92 15.98 179.09 17.345 ;
      RECT 178.975 15.555 179.225 16.11 ;
      RECT 177.275 17.215 177.445 17.675 ;
      RECT 177.275 17.215 177.94 17.385 ;
      RECT 177.71 16.055 177.94 17.385 ;
      RECT 177.275 16.055 177.94 16.225 ;
      RECT 177.275 15.555 177.445 16.225 ;
      RECT 171.295 22.555 171.465 23.205 ;
      RECT 172.135 22.555 172.305 23.2 ;
      RECT 171.295 22.555 172.715 22.725 ;
      RECT 172.54 21.845 172.715 22.725 ;
      RECT 172.54 22.215 175.165 22.385 ;
      RECT 171.215 21.845 172.715 22.015 ;
      RECT 172.055 20.995 172.385 22.015 ;
      RECT 171.215 20.995 171.545 22.015 ;
      RECT 172.055 30.345 172.385 31.365 ;
      RECT 171.215 30.345 171.545 31.365 ;
      RECT 171.215 30.345 172.715 30.515 ;
      RECT 172.54 29.635 172.715 30.515 ;
      RECT 172.54 29.975 175.165 30.145 ;
      RECT 171.295 29.635 172.715 29.805 ;
      RECT 172.135 29.16 172.305 29.805 ;
      RECT 171.295 29.155 171.465 29.805 ;
      RECT 174.15 19.515 174.715 20.485 ;
      RECT 174.255 18.275 174.715 20.485 ;
      RECT 174.15 18.275 174.715 18.845 ;
      RECT 173.195 19.805 173.455 20.485 ;
      RECT 173.195 19.805 173.98 20.025 ;
      RECT 173.78 18.735 173.98 20.025 ;
      RECT 173.78 19.015 174.085 19.345 ;
      RECT 173.195 18.735 173.98 18.905 ;
      RECT 173.195 18.275 173.455 18.905 ;
      RECT 172.735 20.155 173.005 20.485 ;
      RECT 172.835 18.275 173.005 20.485 ;
      RECT 172.835 19.075 173.61 19.635 ;
      RECT 172.735 18.275 173.005 18.605 ;
      RECT 172.77 17.195 173.335 17.765 ;
      RECT 172.875 15.555 173.335 17.765 ;
      RECT 172.77 15.555 173.335 16.525 ;
      RECT 171.815 17.135 172.075 17.765 ;
      RECT 171.815 17.135 172.6 17.305 ;
      RECT 172.4 16.015 172.6 17.305 ;
      RECT 172.4 16.695 172.705 17.025 ;
      RECT 171.815 16.015 172.6 16.235 ;
      RECT 171.815 15.555 172.075 16.235 ;
      RECT 171.665 19.805 172.065 20.485 ;
      RECT 171.665 19.805 172.61 20.025 ;
      RECT 172.375 18.735 172.61 20.025 ;
      RECT 172.375 19.015 172.665 19.345 ;
      RECT 171.665 18.735 172.61 18.905 ;
      RECT 171.665 18.275 172.065 18.905 ;
      RECT 171.355 17.435 171.625 17.765 ;
      RECT 171.455 15.555 171.625 17.765 ;
      RECT 171.455 16.405 172.23 16.965 ;
      RECT 171.355 15.555 171.625 15.885 ;
      RECT 171.685 14.14 171.955 15.045 ;
      RECT 171.775 12.835 171.955 15.045 ;
      RECT 171.695 12.835 171.955 13.34 ;
      RECT 168.075 11.675 168.245 12.325 ;
      RECT 168.915 11.675 169.085 12.32 ;
      RECT 168.075 11.675 169.495 11.845 ;
      RECT 169.32 10.965 169.495 11.845 ;
      RECT 169.32 11.335 171.945 11.505 ;
      RECT 167.995 10.965 169.495 11.135 ;
      RECT 168.835 10.115 169.165 11.135 ;
      RECT 167.995 10.115 168.325 11.135 ;
      RECT 170.825 14.115 171.005 15.045 ;
      RECT 170.825 14.115 171.5 14.285 ;
      RECT 171.33 13.215 171.5 14.285 ;
      RECT 171.33 13.64 171.605 13.97 ;
      RECT 170.835 13.215 171.5 13.385 ;
      RECT 170.835 12.835 171.005 13.385 ;
      RECT 170.285 17.135 170.685 17.765 ;
      RECT 170.285 17.135 171.23 17.305 ;
      RECT 170.995 16.015 171.23 17.305 ;
      RECT 170.995 16.695 171.285 17.025 ;
      RECT 170.285 16.015 171.23 16.235 ;
      RECT 170.285 15.555 170.685 16.235 ;
      RECT 170.265 19.525 170.535 20.475 ;
      RECT 170.265 19.525 171.035 19.745 ;
      RECT 170.745 18.655 171.035 19.745 ;
      RECT 169.805 18.655 171.035 18.855 ;
      RECT 169.805 18.285 170.115 18.855 ;
      RECT 169.855 19.525 170.085 20.475 ;
      RECT 168.925 19.525 169.185 20.475 ;
      RECT 168.925 19.525 170.085 19.765 ;
      RECT 169.395 19.035 169.92 19.345 ;
      RECT 169.395 18.395 169.625 19.345 ;
      RECT 169.275 17.195 169.605 17.715 ;
      RECT 169.485 16.445 169.655 17.28 ;
      RECT 169.43 17.155 169.655 17.28 ;
      RECT 169.44 16.445 169.655 16.575 ;
      RECT 169.265 15.6 169.595 16.525 ;
      RECT 168.435 17.195 168.765 17.72 ;
      RECT 168.565 16.695 168.765 17.72 ;
      RECT 168.565 16.695 169.315 17.025 ;
      RECT 168.565 15.555 168.755 17.72 ;
      RECT 167.86 16.115 168.755 16.49 ;
      RECT 168.415 15.555 168.755 16.49 ;
      RECT 166.905 17.485 167.69 17.655 ;
      RECT 167.52 15.685 167.69 17.655 ;
      RECT 167.52 16.695 168.395 17.025 ;
      RECT 166.805 15.685 167.69 15.855 ;
      RECT 166.885 16.985 167.35 17.315 ;
      RECT 167.03 16.025 167.35 17.315 ;
      RECT 166.33 17.485 166.735 17.655 ;
      RECT 166.33 15.555 166.5 17.655 ;
      RECT 165.67 16.955 166.5 17.255 ;
      RECT 165.67 16.925 165.87 17.255 ;
      RECT 166.33 15.555 166.58 15.885 ;
      RECT 162.555 11.675 162.725 12.325 ;
      RECT 163.395 11.675 163.565 12.32 ;
      RECT 162.555 11.675 163.975 11.845 ;
      RECT 163.8 10.965 163.975 11.845 ;
      RECT 163.8 11.335 166.425 11.505 ;
      RECT 162.475 10.965 163.975 11.135 ;
      RECT 163.315 10.115 163.645 11.135 ;
      RECT 162.475 10.115 162.805 11.135 ;
      RECT 164.785 17.485 165.46 17.655 ;
      RECT 165.29 16.535 165.46 17.655 ;
      RECT 165.99 16.445 166.16 16.775 ;
      RECT 165.29 16.535 166.16 16.705 ;
      RECT 165.65 16.445 166.16 16.705 ;
      RECT 165.65 15.66 165.82 16.705 ;
      RECT 164.715 15.66 165.82 15.83 ;
      RECT 164.595 17.065 165.12 17.285 ;
      RECT 164.95 16 165.12 17.285 ;
      RECT 164.95 16 165.48 16.365 ;
      RECT 164.255 17.485 164.59 17.655 ;
      RECT 164.255 17.215 164.425 17.655 ;
      RECT 164.2 15.98 164.37 17.345 ;
      RECT 164.255 15.555 164.505 16.11 ;
      RECT 162.52 11.305 163.62 11.505 ;
      RECT 162.065 11.305 163.62 11.475 ;
      RECT 162.555 17.215 162.725 17.675 ;
      RECT 162.555 17.215 163.22 17.385 ;
      RECT 162.99 16.055 163.22 17.385 ;
      RECT 162.555 16.055 163.22 16.225 ;
      RECT 162.555 15.555 162.725 16.225 ;
      RECT 158.225 35.835 158.555 36.76 ;
      RECT 158.445 35.08 158.615 35.915 ;
      RECT 158.4 35.785 158.615 35.915 ;
      RECT 158.39 35.08 158.615 35.205 ;
      RECT 158.235 34.645 158.565 35.165 ;
      RECT 157.375 35.87 157.715 36.805 ;
      RECT 157.525 34.64 157.715 36.805 ;
      RECT 156.82 35.87 157.715 36.245 ;
      RECT 157.525 35.335 158.275 35.665 ;
      RECT 157.525 34.64 157.725 35.665 ;
      RECT 157.395 34.64 157.725 35.165 ;
      RECT 157.765 30.395 158.095 31.32 ;
      RECT 157.985 29.64 158.155 30.475 ;
      RECT 157.94 30.345 158.155 30.475 ;
      RECT 157.93 29.64 158.155 29.765 ;
      RECT 157.775 29.205 158.105 29.725 ;
      RECT 156.915 30.43 157.255 31.365 ;
      RECT 157.065 29.2 157.255 31.365 ;
      RECT 156.36 30.43 157.255 30.805 ;
      RECT 157.065 29.895 157.815 30.225 ;
      RECT 157.065 29.2 157.265 30.225 ;
      RECT 156.935 29.2 157.265 29.725 ;
      RECT 155.765 36.505 156.65 36.675 ;
      RECT 156.48 34.705 156.65 36.675 ;
      RECT 156.48 35.335 157.355 35.665 ;
      RECT 155.865 34.705 156.65 34.875 ;
      RECT 153.355 11.675 153.525 12.325 ;
      RECT 154.195 11.675 154.365 12.32 ;
      RECT 153.355 11.675 154.775 11.845 ;
      RECT 154.6 10.965 154.775 11.845 ;
      RECT 154.6 11.335 157.225 11.505 ;
      RECT 153.275 10.965 154.775 11.135 ;
      RECT 154.115 10.115 154.445 11.135 ;
      RECT 153.275 10.115 153.605 11.135 ;
      RECT 155.305 31.065 156.19 31.235 ;
      RECT 156.02 29.265 156.19 31.235 ;
      RECT 156.02 29.895 156.895 30.225 ;
      RECT 155.405 29.265 156.19 29.435 ;
      RECT 155.99 35.045 156.31 36.335 ;
      RECT 155.845 35.045 156.31 35.375 ;
      RECT 156.04 19.815 156.295 20.485 ;
      RECT 156.125 18.275 156.295 20.485 ;
      RECT 156.11 18.275 156.295 18.685 ;
      RECT 156.085 18.275 156.295 18.615 ;
      RECT 156.04 18.275 156.295 18.605 ;
      RECT 156.04 28.315 156.295 28.645 ;
      RECT 156.125 26.435 156.295 28.645 ;
      RECT 156.085 28.305 156.295 28.645 ;
      RECT 156.11 28.235 156.295 28.645 ;
      RECT 156.04 26.435 156.295 27.105 ;
      RECT 156.04 33.755 156.295 34.085 ;
      RECT 156.125 31.875 156.295 34.085 ;
      RECT 156.085 33.745 156.295 34.085 ;
      RECT 156.11 33.675 156.295 34.085 ;
      RECT 156.04 31.875 156.295 32.545 ;
      RECT 152.895 19.475 153.065 20.485 ;
      RECT 152.895 19.475 155.955 19.645 ;
      RECT 155.785 18.755 155.955 19.645 ;
      RECT 155.155 18.755 155.955 18.925 ;
      RECT 152.895 18.755 153.96 18.925 ;
      RECT 153.79 18.275 153.96 18.925 ;
      RECT 155.155 18.275 155.325 18.925 ;
      RECT 152.895 18.275 153.065 18.925 ;
      RECT 153.79 18.275 155.325 18.525 ;
      RECT 153.79 28.395 155.325 28.645 ;
      RECT 155.155 27.995 155.325 28.645 ;
      RECT 152.895 27.995 153.065 28.645 ;
      RECT 153.79 27.995 153.96 28.645 ;
      RECT 155.155 27.995 155.955 28.165 ;
      RECT 155.785 27.275 155.955 28.165 ;
      RECT 152.895 27.995 153.96 28.165 ;
      RECT 152.895 27.275 155.955 27.445 ;
      RECT 152.895 26.435 153.065 27.445 ;
      RECT 153.79 33.835 155.325 34.085 ;
      RECT 155.155 33.435 155.325 34.085 ;
      RECT 152.895 33.435 153.065 34.085 ;
      RECT 153.79 33.435 153.96 34.085 ;
      RECT 155.155 33.435 155.955 33.605 ;
      RECT 155.785 32.715 155.955 33.605 ;
      RECT 152.895 33.435 153.96 33.605 ;
      RECT 152.895 32.715 155.955 32.885 ;
      RECT 152.895 31.875 153.065 32.885 ;
      RECT 155.53 29.605 155.85 30.895 ;
      RECT 155.385 29.605 155.85 29.935 ;
      RECT 155.29 36.475 155.54 36.805 ;
      RECT 155.29 34.705 155.46 36.805 ;
      RECT 154.63 35.105 154.83 35.435 ;
      RECT 154.63 35.105 155.46 35.405 ;
      RECT 155.29 34.705 155.695 34.875 ;
      RECT 155.19 19.125 155.565 19.295 ;
      RECT 155.19 19.095 155.555 19.295 ;
      RECT 155.19 27.625 155.555 27.825 ;
      RECT 155.19 27.625 155.565 27.795 ;
      RECT 155.19 33.065 155.555 33.265 ;
      RECT 155.19 33.065 155.565 33.235 ;
      RECT 155.135 22.555 155.305 23.205 ;
      RECT 154.295 22.555 154.465 23.2 ;
      RECT 153.885 22.555 155.305 22.725 ;
      RECT 153.885 21.845 154.06 22.725 ;
      RECT 151.435 22.215 154.06 22.385 ;
      RECT 153.885 21.845 155.385 22.015 ;
      RECT 155.055 20.995 155.385 22.015 ;
      RECT 154.215 20.995 154.545 22.015 ;
      RECT 155.12 19.815 155.37 20.485 ;
      RECT 153.735 19.815 153.965 20.145 ;
      RECT 153.735 19.815 155.37 20.055 ;
      RECT 153.735 26.865 155.37 27.105 ;
      RECT 155.12 26.435 155.37 27.105 ;
      RECT 153.735 26.775 153.965 27.105 ;
      RECT 153.735 32.305 155.37 32.545 ;
      RECT 155.12 31.875 155.37 32.545 ;
      RECT 153.735 32.215 153.965 32.545 ;
      RECT 154.83 31.035 155.08 31.365 ;
      RECT 154.83 29.265 155 31.365 ;
      RECT 154.17 29.665 154.37 29.995 ;
      RECT 154.17 29.665 155 29.965 ;
      RECT 154.83 29.265 155.235 29.435 ;
      RECT 153.675 36.53 154.78 36.7 ;
      RECT 154.61 35.655 154.78 36.7 ;
      RECT 154.61 35.655 155.12 35.915 ;
      RECT 154.95 35.585 155.12 35.915 ;
      RECT 154.25 35.655 155.12 35.825 ;
      RECT 154.25 34.705 154.42 35.825 ;
      RECT 153.745 34.705 154.42 34.875 ;
      RECT 154.69 19.095 155.02 19.295 ;
      RECT 154.69 18.695 154.975 19.295 ;
      RECT 154.69 27.625 154.975 28.225 ;
      RECT 154.69 27.625 155.02 27.825 ;
      RECT 154.69 33.065 154.975 33.665 ;
      RECT 154.69 33.065 155.02 33.265 ;
      RECT 154.555 17.195 154.885 17.715 ;
      RECT 154.765 16.445 154.935 17.28 ;
      RECT 154.71 17.155 154.935 17.28 ;
      RECT 154.72 16.445 154.935 16.575 ;
      RECT 154.545 15.6 154.875 16.525 ;
      RECT 153.215 31.09 154.32 31.26 ;
      RECT 154.15 30.215 154.32 31.26 ;
      RECT 154.15 30.215 154.66 30.475 ;
      RECT 154.49 30.145 154.66 30.475 ;
      RECT 153.79 30.215 154.66 30.385 ;
      RECT 153.79 29.265 153.96 30.385 ;
      RECT 153.285 29.265 153.96 29.435 ;
      RECT 153.715 17.195 154.045 17.72 ;
      RECT 153.845 16.695 154.045 17.72 ;
      RECT 153.845 16.695 154.595 17.025 ;
      RECT 153.845 15.555 154.035 17.72 ;
      RECT 153.14 16.115 154.035 16.49 ;
      RECT 153.695 15.555 154.035 16.49 ;
      RECT 153.91 35.995 154.44 36.36 ;
      RECT 153.91 35.075 154.08 36.36 ;
      RECT 153.555 35.075 154.08 35.295 ;
      RECT 153.945 19.095 154.42 19.295 ;
      RECT 154.14 18.695 154.42 19.295 ;
      RECT 154.14 27.625 154.42 28.225 ;
      RECT 153.945 27.625 154.42 27.825 ;
      RECT 154.14 33.065 154.42 33.665 ;
      RECT 153.945 33.065 154.42 33.265 ;
      RECT 153.235 20.315 154.405 20.485 ;
      RECT 154.075 20.275 154.405 20.485 ;
      RECT 153.235 19.815 153.565 20.485 ;
      RECT 153.235 26.435 153.565 27.105 ;
      RECT 154.075 26.435 154.405 26.645 ;
      RECT 153.235 26.435 154.405 26.605 ;
      RECT 153.235 31.875 153.565 32.545 ;
      RECT 154.075 31.875 154.405 32.085 ;
      RECT 153.235 31.875 154.405 32.045 ;
      RECT 153.45 30.555 153.98 30.92 ;
      RECT 153.45 29.635 153.62 30.92 ;
      RECT 153.095 29.635 153.62 29.855 ;
      RECT 152.185 17.485 152.97 17.655 ;
      RECT 152.8 15.685 152.97 17.655 ;
      RECT 152.8 16.695 153.675 17.025 ;
      RECT 152.085 15.685 152.97 15.855 ;
      RECT 153.215 36.25 153.465 36.805 ;
      RECT 153.16 35.015 153.33 36.38 ;
      RECT 153.215 34.705 153.385 35.145 ;
      RECT 153.215 34.705 153.55 34.875 ;
      RECT 152.755 30.81 153.005 31.365 ;
      RECT 152.7 29.575 152.87 30.94 ;
      RECT 152.755 29.265 152.925 29.705 ;
      RECT 152.755 29.265 153.09 29.435 ;
      RECT 152.165 16.985 152.63 17.315 ;
      RECT 152.31 16.025 152.63 17.315 ;
      RECT 151.515 36.135 151.685 36.805 ;
      RECT 151.515 36.135 152.18 36.305 ;
      RECT 151.95 34.975 152.18 36.305 ;
      RECT 151.515 34.975 152.18 35.145 ;
      RECT 151.515 34.685 151.685 35.145 ;
      RECT 151.61 17.485 152.015 17.655 ;
      RECT 151.61 15.555 151.78 17.655 ;
      RECT 150.95 16.955 151.78 17.255 ;
      RECT 150.95 16.925 151.15 17.255 ;
      RECT 151.61 15.555 151.86 15.885 ;
      RECT 151.055 30.695 151.225 31.365 ;
      RECT 151.055 30.695 151.72 30.865 ;
      RECT 151.49 29.535 151.72 30.865 ;
      RECT 151.055 29.535 151.72 29.705 ;
      RECT 151.055 29.245 151.225 29.705 ;
      RECT 150.065 17.485 150.74 17.655 ;
      RECT 150.57 16.535 150.74 17.655 ;
      RECT 151.27 16.445 151.44 16.775 ;
      RECT 150.57 16.535 151.44 16.705 ;
      RECT 150.93 16.445 151.44 16.705 ;
      RECT 150.93 15.66 151.1 16.705 ;
      RECT 149.995 15.66 151.1 15.83 ;
      RECT 150.98 19.815 151.235 20.485 ;
      RECT 151.065 18.275 151.235 20.485 ;
      RECT 151.05 18.275 151.235 18.685 ;
      RECT 151.025 18.275 151.235 18.615 ;
      RECT 150.98 18.275 151.235 18.605 ;
      RECT 147.835 19.475 148.005 20.485 ;
      RECT 147.835 19.475 150.895 19.645 ;
      RECT 150.725 18.755 150.895 19.645 ;
      RECT 150.095 18.755 150.895 18.925 ;
      RECT 147.835 18.755 148.9 18.925 ;
      RECT 148.73 18.275 148.9 18.925 ;
      RECT 150.095 18.275 150.265 18.925 ;
      RECT 147.835 18.275 148.005 18.925 ;
      RECT 148.73 18.275 150.265 18.525 ;
      RECT 149.875 17.065 150.4 17.285 ;
      RECT 150.23 16 150.4 17.285 ;
      RECT 150.23 16 150.76 16.365 ;
      RECT 150.13 19.125 150.505 19.295 ;
      RECT 150.13 19.095 150.495 19.295 ;
      RECT 150.06 19.815 150.31 20.485 ;
      RECT 148.675 19.815 148.905 20.145 ;
      RECT 148.675 19.815 150.31 20.055 ;
      RECT 149.63 19.095 149.96 19.295 ;
      RECT 149.63 18.695 149.915 19.295 ;
      RECT 149.535 17.485 149.87 17.655 ;
      RECT 149.535 17.215 149.705 17.655 ;
      RECT 149.48 15.98 149.65 17.345 ;
      RECT 149.535 15.555 149.785 16.11 ;
      RECT 148.885 19.095 149.36 19.295 ;
      RECT 149.08 18.695 149.36 19.295 ;
      RECT 148.175 20.315 149.345 20.485 ;
      RECT 149.015 20.275 149.345 20.485 ;
      RECT 148.175 19.815 148.505 20.485 ;
      RECT 148.645 22.575 148.975 23.205 ;
      RECT 148.725 20.995 148.975 23.205 ;
      RECT 148.645 20.995 148.975 21.975 ;
      RECT 147.835 17.215 148.005 17.675 ;
      RECT 147.835 17.215 148.5 17.385 ;
      RECT 148.27 16.055 148.5 17.385 ;
      RECT 147.835 16.055 148.5 16.225 ;
      RECT 147.835 15.555 148.005 16.225 ;
      RECT 145.355 28.075 145.685 28.595 ;
      RECT 145.565 27.325 145.735 28.16 ;
      RECT 145.51 28.035 145.735 28.16 ;
      RECT 145.52 27.325 145.735 27.455 ;
      RECT 145.345 26.48 145.675 27.405 ;
      RECT 144.515 28.075 144.845 28.6 ;
      RECT 144.645 27.575 144.845 28.6 ;
      RECT 144.645 27.575 145.395 27.905 ;
      RECT 144.645 26.435 144.835 28.6 ;
      RECT 143.94 26.995 144.835 27.37 ;
      RECT 144.495 26.435 144.835 27.37 ;
      RECT 145.04 22.63 145.295 23.205 ;
      RECT 145.125 20.995 145.295 23.205 ;
      RECT 145.04 20.995 145.295 21.9 ;
      RECT 144.155 22.655 144.325 23.205 ;
      RECT 144.155 22.655 144.87 22.825 ;
      RECT 144.7 21.755 144.87 22.825 ;
      RECT 144.7 22.135 144.955 22.465 ;
      RECT 144.155 21.755 144.87 21.925 ;
      RECT 144.155 20.995 144.325 21.925 ;
      RECT 142.985 28.365 143.77 28.535 ;
      RECT 143.6 26.565 143.77 28.535 ;
      RECT 143.6 27.575 144.475 27.905 ;
      RECT 142.885 26.565 143.77 26.735 ;
      RECT 144.095 24.915 144.265 25.925 ;
      RECT 141.205 24.915 144.265 25.085 ;
      RECT 141.205 24.195 141.375 25.085 ;
      RECT 143.2 24.195 144.265 24.365 ;
      RECT 144.095 23.715 144.265 24.365 ;
      RECT 141.205 24.195 142.005 24.365 ;
      RECT 141.835 23.715 142.005 24.365 ;
      RECT 143.2 23.715 143.37 24.365 ;
      RECT 141.835 23.715 143.37 23.965 ;
      RECT 142.755 25.755 143.925 25.925 ;
      RECT 143.595 25.255 143.925 25.925 ;
      RECT 142.755 25.715 143.085 25.925 ;
      RECT 143.2 22.63 143.455 23.205 ;
      RECT 143.285 20.995 143.455 23.205 ;
      RECT 143.2 20.995 143.455 21.9 ;
      RECT 142.965 27.865 143.43 28.195 ;
      RECT 143.11 26.905 143.43 28.195 ;
      RECT 141.79 25.255 142.04 25.925 ;
      RECT 143.195 25.255 143.425 25.585 ;
      RECT 141.79 25.255 143.425 25.495 ;
      RECT 142.74 24.535 143.215 24.735 ;
      RECT 142.74 24.135 143.02 24.735 ;
      RECT 142.315 22.655 142.485 23.205 ;
      RECT 142.315 22.655 143.03 22.825 ;
      RECT 142.86 21.755 143.03 22.825 ;
      RECT 142.86 22.135 143.115 22.465 ;
      RECT 142.315 21.755 143.03 21.925 ;
      RECT 142.315 20.995 142.485 21.925 ;
      RECT 142.41 28.365 142.815 28.535 ;
      RECT 142.41 26.435 142.58 28.535 ;
      RECT 141.75 27.835 142.58 28.135 ;
      RECT 141.75 27.805 141.95 28.135 ;
      RECT 142.41 26.435 142.66 26.765 ;
      RECT 139.395 14.025 139.725 15.045 ;
      RECT 138.555 14.025 138.885 15.045 ;
      RECT 138.555 14.025 140.055 14.195 ;
      RECT 139.88 13.315 140.055 14.195 ;
      RECT 139.88 13.655 142.505 13.825 ;
      RECT 138.635 13.315 140.055 13.485 ;
      RECT 139.475 12.84 139.645 13.485 ;
      RECT 138.635 12.835 138.805 13.485 ;
      RECT 142.14 24.535 142.47 24.735 ;
      RECT 142.185 24.135 142.47 24.735 ;
      RECT 140.865 28.365 141.54 28.535 ;
      RECT 141.37 27.415 141.54 28.535 ;
      RECT 142.07 27.325 142.24 27.655 ;
      RECT 141.37 27.415 142.24 27.585 ;
      RECT 141.73 27.325 142.24 27.585 ;
      RECT 141.73 26.54 141.9 27.585 ;
      RECT 140.795 26.54 141.9 26.71 ;
      RECT 141.595 24.565 141.97 24.735 ;
      RECT 141.605 24.535 141.97 24.735 ;
      RECT 140.675 27.945 141.2 28.165 ;
      RECT 141.03 26.88 141.2 28.165 ;
      RECT 141.03 26.88 141.56 27.245 ;
      RECT 140.865 25.255 141.12 25.925 ;
      RECT 140.865 23.715 141.035 25.925 ;
      RECT 140.865 23.715 141.05 24.125 ;
      RECT 140.865 23.715 141.12 24.045 ;
      RECT 140.335 28.365 140.67 28.535 ;
      RECT 140.335 28.095 140.505 28.535 ;
      RECT 140.28 26.86 140.45 28.225 ;
      RECT 140.335 26.435 140.585 26.99 ;
      RECT 139.835 17.195 140.165 17.715 ;
      RECT 140.045 16.445 140.215 17.28 ;
      RECT 139.99 17.155 140.215 17.28 ;
      RECT 140 16.445 140.215 16.575 ;
      RECT 139.825 15.6 140.155 16.525 ;
      RECT 139.825 19.515 140.155 20.44 ;
      RECT 140.045 18.76 140.215 19.595 ;
      RECT 140 19.465 140.215 19.595 ;
      RECT 139.99 18.76 140.215 18.885 ;
      RECT 139.835 18.325 140.165 18.845 ;
      RECT 138.995 17.195 139.325 17.72 ;
      RECT 139.125 16.695 139.325 17.72 ;
      RECT 139.125 16.695 139.875 17.025 ;
      RECT 139.125 15.555 139.315 17.72 ;
      RECT 138.42 16.115 139.315 16.49 ;
      RECT 138.975 15.555 139.315 16.49 ;
      RECT 138.975 19.55 139.315 20.485 ;
      RECT 139.125 18.32 139.315 20.485 ;
      RECT 138.42 19.55 139.315 19.925 ;
      RECT 139.125 19.015 139.875 19.345 ;
      RECT 139.125 18.32 139.325 19.345 ;
      RECT 138.995 18.32 139.325 18.845 ;
      RECT 138.635 28.095 138.805 28.555 ;
      RECT 138.635 28.095 139.3 28.265 ;
      RECT 139.07 26.935 139.3 28.265 ;
      RECT 138.635 26.935 139.3 27.105 ;
      RECT 138.635 26.435 138.805 27.105 ;
      RECT 137.465 17.485 138.25 17.655 ;
      RECT 138.08 15.685 138.25 17.655 ;
      RECT 138.08 16.695 138.955 17.025 ;
      RECT 137.365 15.685 138.25 15.855 ;
      RECT 137.365 20.185 138.25 20.355 ;
      RECT 138.08 18.385 138.25 20.355 ;
      RECT 138.08 19.015 138.955 19.345 ;
      RECT 137.465 18.385 138.25 18.555 ;
      RECT 138.115 22.555 138.285 23.205 ;
      RECT 135.855 22.955 137.39 23.205 ;
      RECT 137.22 22.555 137.39 23.205 ;
      RECT 135.855 22.555 136.025 23.205 ;
      RECT 137.22 22.555 138.285 22.725 ;
      RECT 135.225 22.555 136.025 22.725 ;
      RECT 135.225 21.835 135.395 22.725 ;
      RECT 135.225 21.835 138.285 22.005 ;
      RECT 138.115 20.995 138.285 22.005 ;
      RECT 137.615 20.995 137.945 21.665 ;
      RECT 136.775 20.995 137.105 21.205 ;
      RECT 136.775 20.995 137.945 21.165 ;
      RECT 137.445 16.985 137.91 17.315 ;
      RECT 137.59 16.025 137.91 17.315 ;
      RECT 137.59 18.725 137.91 20.015 ;
      RECT 137.445 18.725 137.91 19.055 ;
      RECT 137.655 24.915 137.825 25.925 ;
      RECT 134.765 24.915 137.825 25.085 ;
      RECT 134.765 24.195 134.935 25.085 ;
      RECT 136.76 24.195 137.825 24.365 ;
      RECT 137.655 23.715 137.825 24.365 ;
      RECT 134.765 24.195 135.565 24.365 ;
      RECT 135.395 23.715 135.565 24.365 ;
      RECT 136.76 23.715 136.93 24.365 ;
      RECT 135.395 23.715 136.93 23.965 ;
      RECT 136.315 25.755 137.485 25.925 ;
      RECT 137.155 25.255 137.485 25.925 ;
      RECT 136.315 25.715 136.645 25.925 ;
      RECT 135.81 21.425 137.445 21.665 ;
      RECT 137.215 21.335 137.445 21.665 ;
      RECT 135.81 20.995 136.06 21.665 ;
      RECT 136.89 17.485 137.295 17.655 ;
      RECT 136.89 15.555 137.06 17.655 ;
      RECT 136.23 16.955 137.06 17.255 ;
      RECT 136.23 16.925 136.43 17.255 ;
      RECT 136.89 15.555 137.14 15.885 ;
      RECT 136.89 20.155 137.14 20.485 ;
      RECT 136.89 18.385 137.06 20.485 ;
      RECT 136.23 18.785 136.43 19.115 ;
      RECT 136.23 18.785 137.06 19.085 ;
      RECT 136.89 18.385 137.295 18.555 ;
      RECT 136.76 22.185 137.04 22.785 ;
      RECT 136.76 22.185 137.235 22.385 ;
      RECT 133.115 11.675 133.285 12.325 ;
      RECT 133.955 11.675 134.125 12.32 ;
      RECT 133.115 11.675 134.535 11.845 ;
      RECT 134.36 10.965 134.535 11.845 ;
      RECT 134.36 11.335 136.985 11.505 ;
      RECT 133.035 10.965 134.535 11.135 ;
      RECT 133.875 10.115 134.205 11.135 ;
      RECT 133.035 10.115 133.365 11.135 ;
      RECT 135.35 25.255 135.6 25.925 ;
      RECT 136.755 25.255 136.985 25.585 ;
      RECT 135.35 25.255 136.985 25.495 ;
      RECT 136.3 24.535 136.775 24.735 ;
      RECT 136.3 24.135 136.58 24.735 ;
      RECT 135.345 17.485 136.02 17.655 ;
      RECT 135.85 16.535 136.02 17.655 ;
      RECT 136.55 16.445 136.72 16.775 ;
      RECT 135.85 16.535 136.72 16.705 ;
      RECT 136.21 16.445 136.72 16.705 ;
      RECT 136.21 15.66 136.38 16.705 ;
      RECT 135.275 15.66 136.38 15.83 ;
      RECT 135.275 20.21 136.38 20.38 ;
      RECT 136.21 19.335 136.38 20.38 ;
      RECT 136.21 19.335 136.72 19.595 ;
      RECT 136.55 19.265 136.72 19.595 ;
      RECT 135.85 19.335 136.72 19.505 ;
      RECT 135.85 18.385 136.02 19.505 ;
      RECT 135.345 18.385 136.02 18.555 ;
      RECT 136.205 22.185 136.49 22.785 ;
      RECT 136.16 22.185 136.49 22.385 ;
      RECT 135.155 17.065 135.68 17.285 ;
      RECT 135.51 16 135.68 17.285 ;
      RECT 135.51 16 136.04 16.365 ;
      RECT 135.51 19.675 136.04 20.04 ;
      RECT 135.51 18.755 135.68 20.04 ;
      RECT 135.155 18.755 135.68 18.975 ;
      RECT 135.7 24.535 136.03 24.735 ;
      RECT 135.745 24.135 136.03 24.735 ;
      RECT 135.625 22.185 135.99 22.385 ;
      RECT 135.615 22.185 135.99 22.355 ;
      RECT 135.155 24.565 135.53 24.735 ;
      RECT 135.165 24.535 135.53 24.735 ;
      RECT 134.815 17.485 135.15 17.655 ;
      RECT 134.815 17.215 134.985 17.655 ;
      RECT 134.76 15.98 134.93 17.345 ;
      RECT 134.815 15.555 135.065 16.11 ;
      RECT 134.815 19.93 135.065 20.485 ;
      RECT 134.76 18.695 134.93 20.06 ;
      RECT 134.815 18.385 134.985 18.825 ;
      RECT 134.815 18.385 135.15 18.555 ;
      RECT 134.885 22.875 135.14 23.205 ;
      RECT 134.885 22.795 135.07 23.205 ;
      RECT 134.885 20.995 135.055 23.205 ;
      RECT 134.885 20.995 135.095 21.675 ;
      RECT 134.885 20.995 135.14 21.665 ;
      RECT 134.425 25.255 134.68 25.925 ;
      RECT 134.425 23.715 134.595 25.925 ;
      RECT 134.425 23.715 134.61 24.125 ;
      RECT 134.425 23.715 134.635 24.055 ;
      RECT 134.425 23.715 134.68 24.045 ;
      RECT 133.115 17.215 133.285 17.675 ;
      RECT 133.115 17.215 133.78 17.385 ;
      RECT 133.55 16.055 133.78 17.385 ;
      RECT 133.115 16.055 133.78 16.225 ;
      RECT 133.115 15.555 133.285 16.225 ;
      RECT 133.115 19.815 133.285 20.485 ;
      RECT 133.115 19.815 133.78 19.985 ;
      RECT 133.55 18.655 133.78 19.985 ;
      RECT 133.115 18.655 133.78 18.825 ;
      RECT 133.115 18.365 133.285 18.825 ;
      RECT 131.66 22.875 131.915 23.205 ;
      RECT 131.745 20.995 131.915 23.205 ;
      RECT 131.705 22.865 131.915 23.205 ;
      RECT 131.73 22.795 131.915 23.205 ;
      RECT 131.66 20.995 131.915 21.665 ;
      RECT 129.41 22.955 130.945 23.205 ;
      RECT 130.775 22.555 130.945 23.205 ;
      RECT 128.515 22.555 128.685 23.205 ;
      RECT 129.41 22.555 129.58 23.205 ;
      RECT 130.775 22.555 131.575 22.725 ;
      RECT 131.405 21.835 131.575 22.725 ;
      RECT 128.515 22.555 129.58 22.725 ;
      RECT 128.515 21.835 131.575 22.005 ;
      RECT 128.515 20.995 128.685 22.005 ;
      RECT 131.085 35.835 131.415 36.76 ;
      RECT 131.305 35.08 131.475 35.915 ;
      RECT 131.26 35.785 131.475 35.915 ;
      RECT 131.25 35.08 131.475 35.205 ;
      RECT 131.095 34.645 131.425 35.165 ;
      RECT 130.81 22.185 131.175 22.385 ;
      RECT 130.81 22.185 131.185 22.355 ;
      RECT 130.235 35.87 130.575 36.805 ;
      RECT 130.385 34.64 130.575 36.805 ;
      RECT 129.68 35.87 130.575 36.245 ;
      RECT 130.385 35.335 131.135 35.665 ;
      RECT 130.385 34.64 130.585 35.665 ;
      RECT 130.255 34.64 130.585 35.165 ;
      RECT 122.845 12.86 123.07 15.045 ;
      RECT 121.095 14.035 121.35 15.045 ;
      RECT 130.745 14.035 131 15.03 ;
      RECT 129.885 14.035 130.125 15.03 ;
      RECT 129.025 12.86 129.275 15.03 ;
      RECT 128.165 12.86 128.415 15.03 ;
      RECT 127.305 12.86 127.555 15.03 ;
      RECT 126.445 12.86 126.695 15.03 ;
      RECT 125.425 13.995 125.8 15.03 ;
      RECT 124.535 12.86 124.775 15.03 ;
      RECT 123.675 12.86 123.93 15.03 ;
      RECT 121.955 14.035 122.21 15.03 ;
      RECT 121.955 14.705 122.215 14.875 ;
      RECT 121.095 14.035 131 14.245 ;
      RECT 122.845 13.995 129.275 14.245 ;
      RECT 125.425 12.86 125.775 15.03 ;
      RECT 129.355 21.425 130.99 21.665 ;
      RECT 130.74 20.995 130.99 21.665 ;
      RECT 129.355 21.335 129.585 21.665 ;
      RECT 130.31 22.185 130.595 22.785 ;
      RECT 130.31 22.185 130.64 22.385 ;
      RECT 130.295 27.995 130.465 28.645 ;
      RECT 128.035 28.395 129.57 28.645 ;
      RECT 129.4 27.995 129.57 28.645 ;
      RECT 128.035 27.995 128.205 28.645 ;
      RECT 129.4 27.995 130.465 28.165 ;
      RECT 127.405 27.995 128.205 28.165 ;
      RECT 127.405 27.275 127.575 28.165 ;
      RECT 127.405 27.275 130.465 27.445 ;
      RECT 130.295 26.435 130.465 27.445 ;
      RECT 128.625 36.505 129.51 36.675 ;
      RECT 129.34 34.705 129.51 36.675 ;
      RECT 129.34 35.335 130.215 35.665 ;
      RECT 128.725 34.705 129.51 34.875 ;
      RECT 129.795 26.435 130.125 27.105 ;
      RECT 128.955 26.435 129.285 26.645 ;
      RECT 128.955 26.435 130.125 26.605 ;
      RECT 129.76 22.185 130.04 22.785 ;
      RECT 129.565 22.185 130.04 22.385 ;
      RECT 128.855 20.995 129.185 21.665 ;
      RECT 129.695 20.995 130.025 21.205 ;
      RECT 128.855 20.995 130.025 21.165 ;
      RECT 127.99 26.865 129.625 27.105 ;
      RECT 129.395 26.775 129.625 27.105 ;
      RECT 127.99 26.435 128.24 27.105 ;
      RECT 128.94 27.625 129.22 28.225 ;
      RECT 128.94 27.625 129.415 27.825 ;
      RECT 128.85 35.045 129.17 36.335 ;
      RECT 128.705 35.045 129.17 35.375 ;
      RECT 128.385 27.625 128.67 28.225 ;
      RECT 128.34 27.625 128.67 27.825 ;
      RECT 128.15 36.475 128.4 36.805 ;
      RECT 128.15 34.705 128.32 36.805 ;
      RECT 127.49 35.105 127.69 35.435 ;
      RECT 127.49 35.105 128.32 35.405 ;
      RECT 128.15 34.705 128.555 34.875 ;
      RECT 127.875 22.635 128.205 23.155 ;
      RECT 128.085 21.885 128.255 22.72 ;
      RECT 128.03 22.595 128.255 22.72 ;
      RECT 128.04 21.885 128.255 22.015 ;
      RECT 127.865 21.04 128.195 21.965 ;
      RECT 124.375 11.675 124.545 12.325 ;
      RECT 125.215 11.675 125.385 12.32 ;
      RECT 124.375 11.675 125.795 11.845 ;
      RECT 125.62 10.965 125.795 11.845 ;
      RECT 125.62 11.335 128.245 11.505 ;
      RECT 124.295 10.965 125.795 11.135 ;
      RECT 125.135 10.115 125.465 11.135 ;
      RECT 124.295 10.115 124.625 11.135 ;
      RECT 127.805 27.625 128.17 27.825 ;
      RECT 127.795 27.625 128.17 27.795 ;
      RECT 126.535 36.53 127.64 36.7 ;
      RECT 127.47 35.655 127.64 36.7 ;
      RECT 127.47 35.655 127.98 35.915 ;
      RECT 127.81 35.585 127.98 35.915 ;
      RECT 127.11 35.655 127.98 35.825 ;
      RECT 127.11 34.705 127.28 35.825 ;
      RECT 126.605 34.705 127.28 34.875 ;
      RECT 127.035 22.635 127.365 23.16 ;
      RECT 127.165 22.135 127.365 23.16 ;
      RECT 127.165 22.135 127.915 22.465 ;
      RECT 127.165 20.995 127.355 23.16 ;
      RECT 126.46 21.555 127.355 21.93 ;
      RECT 127.015 20.995 127.355 21.93 ;
      RECT 126.52 19.48 126.78 20.455 ;
      RECT 125.665 19.48 125.92 20.455 ;
      RECT 124.805 19.48 125.06 20.455 ;
      RECT 124.305 19.48 127.335 19.65 ;
      RECT 127.035 18.745 127.335 19.65 ;
      RECT 124.305 18.745 124.475 19.65 ;
      RECT 124.305 18.745 127.335 18.915 ;
      RECT 126.09 18.3 126.345 18.915 ;
      RECT 125.23 18.3 125.49 18.915 ;
      RECT 127.065 28.315 127.32 28.645 ;
      RECT 127.065 28.305 127.275 28.645 ;
      RECT 127.065 28.235 127.25 28.645 ;
      RECT 127.065 26.435 127.235 28.645 ;
      RECT 127.065 26.435 127.32 27.105 ;
      RECT 126.77 35.995 127.3 36.36 ;
      RECT 126.77 35.075 126.94 36.36 ;
      RECT 126.415 35.075 126.94 35.295 ;
      RECT 125.505 22.925 126.29 23.095 ;
      RECT 126.12 21.125 126.29 23.095 ;
      RECT 126.12 22.135 126.995 22.465 ;
      RECT 125.405 21.125 126.29 21.295 ;
      RECT 126.075 36.25 126.325 36.805 ;
      RECT 126.02 35.015 126.19 36.38 ;
      RECT 126.075 34.705 126.245 35.145 ;
      RECT 126.075 34.705 126.41 34.875 ;
      RECT 125.485 22.425 125.95 22.755 ;
      RECT 125.63 21.465 125.95 22.755 ;
      RECT 125.115 17.195 125.445 17.715 ;
      RECT 125.325 16.445 125.495 17.28 ;
      RECT 125.27 17.155 125.495 17.28 ;
      RECT 125.28 16.445 125.495 16.575 ;
      RECT 125.105 15.6 125.435 16.525 ;
      RECT 124.93 22.925 125.335 23.095 ;
      RECT 124.93 20.995 125.1 23.095 ;
      RECT 124.27 22.395 125.1 22.695 ;
      RECT 124.27 22.365 124.47 22.695 ;
      RECT 124.93 20.995 125.18 21.325 ;
      RECT 124.275 17.195 124.605 17.72 ;
      RECT 124.405 16.695 124.605 17.72 ;
      RECT 124.405 16.695 125.155 17.025 ;
      RECT 124.405 15.555 124.595 17.72 ;
      RECT 123.7 16.115 124.595 16.49 ;
      RECT 124.255 15.555 124.595 16.49 ;
      RECT 124.375 36.135 124.545 36.805 ;
      RECT 124.375 36.135 125.04 36.305 ;
      RECT 124.81 34.975 125.04 36.305 ;
      RECT 124.375 34.975 125.04 35.145 ;
      RECT 124.375 34.685 124.545 35.145 ;
      RECT 123.385 22.925 124.06 23.095 ;
      RECT 123.89 21.975 124.06 23.095 ;
      RECT 124.59 21.885 124.76 22.215 ;
      RECT 123.89 21.975 124.76 22.145 ;
      RECT 124.25 21.885 124.76 22.145 ;
      RECT 124.25 21.1 124.42 22.145 ;
      RECT 123.315 21.1 124.42 21.27 ;
      RECT 122.745 17.485 123.53 17.655 ;
      RECT 123.36 15.685 123.53 17.655 ;
      RECT 123.36 16.695 124.235 17.025 ;
      RECT 122.645 15.685 123.53 15.855 ;
      RECT 123.195 22.505 123.72 22.725 ;
      RECT 123.55 21.44 123.72 22.725 ;
      RECT 123.55 21.44 124.08 21.805 ;
      RECT 122.725 16.985 123.19 17.315 ;
      RECT 122.87 16.025 123.19 17.315 ;
      RECT 122.855 22.925 123.19 23.095 ;
      RECT 122.855 22.655 123.025 23.095 ;
      RECT 122.8 21.42 122.97 22.785 ;
      RECT 122.855 20.995 123.105 21.55 ;
      RECT 122.17 17.485 122.575 17.655 ;
      RECT 122.17 15.555 122.34 17.655 ;
      RECT 121.51 16.955 122.34 17.255 ;
      RECT 121.51 16.925 121.71 17.255 ;
      RECT 122.17 15.555 122.42 15.885 ;
      RECT 118.395 11.675 118.565 12.325 ;
      RECT 119.235 11.675 119.405 12.32 ;
      RECT 118.395 11.675 119.815 11.845 ;
      RECT 119.64 10.965 119.815 11.845 ;
      RECT 119.64 11.335 122.265 11.505 ;
      RECT 118.315 10.965 119.815 11.135 ;
      RECT 119.155 10.115 119.485 11.135 ;
      RECT 118.315 10.115 118.645 11.135 ;
      RECT 120.625 17.485 121.3 17.655 ;
      RECT 121.13 16.535 121.3 17.655 ;
      RECT 121.83 16.445 122 16.775 ;
      RECT 121.13 16.535 122 16.705 ;
      RECT 121.49 16.445 122 16.705 ;
      RECT 121.49 15.66 121.66 16.705 ;
      RECT 120.555 15.66 121.66 15.83 ;
      RECT 121.155 22.655 121.325 23.115 ;
      RECT 121.155 22.655 121.82 22.825 ;
      RECT 121.59 21.495 121.82 22.825 ;
      RECT 121.155 21.495 121.82 21.665 ;
      RECT 121.155 20.995 121.325 21.665 ;
      RECT 120.54 19.48 120.8 20.455 ;
      RECT 119.685 19.48 119.94 20.455 ;
      RECT 118.825 19.48 119.08 20.455 ;
      RECT 118.325 19.48 121.355 19.65 ;
      RECT 121.055 18.745 121.355 19.65 ;
      RECT 118.325 18.745 118.495 19.65 ;
      RECT 118.325 18.745 121.355 18.915 ;
      RECT 120.11 18.3 120.365 18.915 ;
      RECT 119.25 18.3 119.51 18.915 ;
      RECT 120.435 17.065 120.96 17.285 ;
      RECT 120.79 16 120.96 17.285 ;
      RECT 120.79 16 121.32 16.365 ;
      RECT 120.095 17.485 120.43 17.655 ;
      RECT 120.095 17.215 120.265 17.655 ;
      RECT 120.04 15.98 120.21 17.345 ;
      RECT 120.095 15.555 120.345 16.11 ;
      RECT 118.395 17.215 118.565 17.675 ;
      RECT 118.395 17.215 119.06 17.385 ;
      RECT 118.83 16.055 119.06 17.385 ;
      RECT 118.395 16.055 119.06 16.225 ;
      RECT 118.395 15.555 118.565 16.225 ;
      RECT 117.295 28.075 117.625 28.595 ;
      RECT 117.505 27.325 117.675 28.16 ;
      RECT 117.45 28.035 117.675 28.16 ;
      RECT 117.46 27.325 117.675 27.455 ;
      RECT 117.285 26.48 117.615 27.405 ;
      RECT 117.4 14.375 117.655 15.045 ;
      RECT 117.485 12.835 117.655 15.045 ;
      RECT 117.47 12.835 117.655 13.245 ;
      RECT 117.4 12.835 117.655 13.165 ;
      RECT 117.4 22.875 117.655 23.205 ;
      RECT 117.485 20.995 117.655 23.205 ;
      RECT 117.445 22.865 117.655 23.205 ;
      RECT 117.47 22.795 117.655 23.205 ;
      RECT 117.4 20.995 117.655 21.665 ;
      RECT 116.455 28.075 116.785 28.6 ;
      RECT 116.585 27.575 116.785 28.6 ;
      RECT 116.585 27.575 117.335 27.905 ;
      RECT 116.585 26.435 116.775 28.6 ;
      RECT 115.88 26.995 116.775 27.37 ;
      RECT 116.435 26.435 116.775 27.37 ;
      RECT 114.255 14.035 114.425 15.045 ;
      RECT 114.255 14.035 117.315 14.205 ;
      RECT 117.145 13.315 117.315 14.205 ;
      RECT 116.515 13.315 117.315 13.485 ;
      RECT 114.255 13.315 115.32 13.485 ;
      RECT 115.15 12.835 115.32 13.485 ;
      RECT 116.515 12.835 116.685 13.485 ;
      RECT 114.255 12.835 114.425 13.485 ;
      RECT 115.15 12.835 116.685 13.085 ;
      RECT 115.15 22.955 116.685 23.205 ;
      RECT 116.515 22.555 116.685 23.205 ;
      RECT 114.255 22.555 114.425 23.205 ;
      RECT 115.15 22.555 115.32 23.205 ;
      RECT 116.515 22.555 117.315 22.725 ;
      RECT 117.145 21.835 117.315 22.725 ;
      RECT 114.255 22.555 115.32 22.725 ;
      RECT 114.255 21.835 117.315 22.005 ;
      RECT 114.255 20.995 114.425 22.005 ;
      RECT 116.825 19.515 117.155 20.44 ;
      RECT 117.045 18.76 117.215 19.595 ;
      RECT 117 19.465 117.215 19.595 ;
      RECT 116.99 18.76 117.215 18.885 ;
      RECT 116.835 18.325 117.165 18.845 ;
      RECT 116.55 13.685 116.925 13.855 ;
      RECT 116.55 13.655 116.915 13.855 ;
      RECT 116.55 22.185 116.915 22.385 ;
      RECT 116.55 22.185 116.925 22.355 ;
      RECT 115.975 19.55 116.315 20.485 ;
      RECT 116.125 18.32 116.315 20.485 ;
      RECT 115.42 19.55 116.315 19.925 ;
      RECT 116.125 19.015 116.875 19.345 ;
      RECT 116.125 18.32 116.325 19.345 ;
      RECT 115.995 18.32 116.325 18.845 ;
      RECT 116.48 14.375 116.73 15.045 ;
      RECT 115.095 14.375 115.325 14.705 ;
      RECT 115.095 14.375 116.73 14.615 ;
      RECT 115.095 21.425 116.73 21.665 ;
      RECT 116.48 20.995 116.73 21.665 ;
      RECT 115.095 21.335 115.325 21.665 ;
      RECT 114.925 28.365 115.71 28.535 ;
      RECT 115.54 26.565 115.71 28.535 ;
      RECT 115.54 27.575 116.415 27.905 ;
      RECT 114.825 26.565 115.71 26.735 ;
      RECT 116.05 13.655 116.38 13.855 ;
      RECT 116.05 13.255 116.335 13.855 ;
      RECT 116.05 22.185 116.335 22.785 ;
      RECT 116.05 22.185 116.38 22.385 ;
      RECT 113.175 24.905 113.505 25.925 ;
      RECT 112.335 24.905 112.665 25.925 ;
      RECT 112.335 24.905 113.835 25.075 ;
      RECT 113.66 24.195 113.835 25.075 ;
      RECT 113.66 24.535 116.285 24.705 ;
      RECT 112.415 24.195 113.835 24.365 ;
      RECT 113.255 23.72 113.425 24.365 ;
      RECT 112.415 23.715 112.585 24.365 ;
      RECT 116.02 17.435 116.275 17.765 ;
      RECT 116.105 15.555 116.275 17.765 ;
      RECT 116.065 17.425 116.275 17.765 ;
      RECT 116.09 17.355 116.275 17.765 ;
      RECT 116.02 15.555 116.275 16.225 ;
      RECT 114.365 20.185 115.25 20.355 ;
      RECT 115.08 18.385 115.25 20.355 ;
      RECT 115.08 19.015 115.955 19.345 ;
      RECT 114.465 18.385 115.25 18.555 ;
      RECT 113.77 17.515 115.305 17.765 ;
      RECT 115.135 17.115 115.305 17.765 ;
      RECT 112.875 17.115 113.045 17.765 ;
      RECT 113.77 17.115 113.94 17.765 ;
      RECT 115.135 17.115 115.935 17.285 ;
      RECT 115.765 16.395 115.935 17.285 ;
      RECT 112.875 17.115 113.94 17.285 ;
      RECT 112.875 16.395 115.935 16.565 ;
      RECT 112.875 15.555 113.045 16.565 ;
      RECT 115.305 13.655 115.78 13.855 ;
      RECT 115.5 13.255 115.78 13.855 ;
      RECT 115.5 22.185 115.78 22.785 ;
      RECT 115.305 22.185 115.78 22.385 ;
      RECT 114.595 14.875 115.765 15.045 ;
      RECT 115.435 14.835 115.765 15.045 ;
      RECT 114.595 14.375 114.925 15.045 ;
      RECT 114.595 20.995 114.925 21.665 ;
      RECT 115.435 20.995 115.765 21.205 ;
      RECT 114.595 20.995 115.765 21.165 ;
      RECT 115.17 16.745 115.535 16.945 ;
      RECT 115.17 16.745 115.545 16.915 ;
      RECT 114.905 27.865 115.37 28.195 ;
      RECT 115.05 26.905 115.37 28.195 ;
      RECT 115.115 11.675 115.285 12.325 ;
      RECT 114.275 11.675 114.445 12.32 ;
      RECT 113.865 11.675 115.285 11.845 ;
      RECT 113.865 10.965 114.04 11.845 ;
      RECT 111.415 11.335 114.04 11.505 ;
      RECT 113.865 10.965 115.365 11.135 ;
      RECT 115.035 10.115 115.365 11.135 ;
      RECT 114.195 10.115 114.525 11.135 ;
      RECT 113.715 15.985 115.35 16.225 ;
      RECT 115.1 15.555 115.35 16.225 ;
      RECT 113.715 15.895 113.945 16.225 ;
      RECT 114.67 16.745 114.955 17.345 ;
      RECT 114.67 16.745 115 16.945 ;
      RECT 114.59 18.725 114.91 20.015 ;
      RECT 114.445 18.725 114.91 19.055 ;
      RECT 114.35 28.365 114.755 28.535 ;
      RECT 114.35 26.435 114.52 28.535 ;
      RECT 113.69 27.835 114.52 28.135 ;
      RECT 113.69 27.805 113.89 28.135 ;
      RECT 114.35 26.435 114.6 26.765 ;
      RECT 114.065 30.395 114.395 31.32 ;
      RECT 114.285 29.64 114.455 30.475 ;
      RECT 114.24 30.345 114.455 30.475 ;
      RECT 114.23 29.64 114.455 29.765 ;
      RECT 114.075 29.205 114.405 29.725 ;
      RECT 114.12 16.745 114.4 17.345 ;
      RECT 113.925 16.745 114.4 16.945 ;
      RECT 113.215 15.555 113.545 16.225 ;
      RECT 114.055 15.555 114.385 15.765 ;
      RECT 113.215 15.555 114.385 15.725 ;
      RECT 113.89 20.155 114.14 20.485 ;
      RECT 113.89 18.385 114.06 20.485 ;
      RECT 113.23 18.785 113.43 19.115 ;
      RECT 113.23 18.785 114.06 19.085 ;
      RECT 113.89 18.385 114.295 18.555 ;
      RECT 112.805 28.365 113.48 28.535 ;
      RECT 113.31 27.415 113.48 28.535 ;
      RECT 114.01 27.325 114.18 27.655 ;
      RECT 113.31 27.415 114.18 27.585 ;
      RECT 113.67 27.325 114.18 27.585 ;
      RECT 113.67 26.54 113.84 27.585 ;
      RECT 112.735 26.54 113.84 26.71 ;
      RECT 113.215 30.43 113.555 31.365 ;
      RECT 113.365 29.2 113.555 31.365 ;
      RECT 112.66 30.43 113.555 30.805 ;
      RECT 113.365 29.895 114.115 30.225 ;
      RECT 113.365 29.2 113.565 30.225 ;
      RECT 113.235 29.2 113.565 29.725 ;
      RECT 112.275 20.21 113.38 20.38 ;
      RECT 113.21 19.335 113.38 20.38 ;
      RECT 113.21 19.335 113.72 19.595 ;
      RECT 113.55 19.265 113.72 19.595 ;
      RECT 112.85 19.335 113.72 19.505 ;
      RECT 112.85 18.385 113.02 19.505 ;
      RECT 112.345 18.385 113.02 18.555 ;
      RECT 112.615 27.945 113.14 28.165 ;
      RECT 112.97 26.88 113.14 28.165 ;
      RECT 112.97 26.88 113.5 27.245 ;
      RECT 111.605 31.065 112.49 31.235 ;
      RECT 112.32 29.265 112.49 31.235 ;
      RECT 112.32 29.895 113.195 30.225 ;
      RECT 111.705 29.265 112.49 29.435 ;
      RECT 112.51 19.675 113.04 20.04 ;
      RECT 112.51 18.755 112.68 20.04 ;
      RECT 112.155 18.755 112.68 18.975 ;
      RECT 112.275 28.365 112.61 28.535 ;
      RECT 112.275 28.095 112.445 28.535 ;
      RECT 112.22 26.86 112.39 28.225 ;
      RECT 112.275 26.435 112.525 26.99 ;
      RECT 111.815 19.93 112.065 20.485 ;
      RECT 111.76 18.695 111.93 20.06 ;
      RECT 111.815 18.385 111.985 18.825 ;
      RECT 111.815 18.385 112.15 18.555 ;
      RECT 111.83 29.605 112.15 30.895 ;
      RECT 111.685 29.605 112.15 29.935 ;
      RECT 111.895 22.555 112.065 23.205 ;
      RECT 109.635 22.955 111.17 23.205 ;
      RECT 111 22.555 111.17 23.205 ;
      RECT 109.635 22.555 109.805 23.205 ;
      RECT 111 22.555 112.065 22.725 ;
      RECT 109.005 22.555 109.805 22.725 ;
      RECT 109.005 21.835 109.175 22.725 ;
      RECT 109.005 21.835 112.065 22.005 ;
      RECT 111.895 20.995 112.065 22.005 ;
      RECT 111.395 20.995 111.725 21.665 ;
      RECT 110.555 20.995 110.885 21.205 ;
      RECT 110.555 20.995 111.725 21.165 ;
      RECT 111.13 31.035 111.38 31.365 ;
      RECT 111.13 29.265 111.3 31.365 ;
      RECT 110.47 29.665 110.67 29.995 ;
      RECT 110.47 29.665 111.3 29.965 ;
      RECT 111.13 29.265 111.535 29.435 ;
      RECT 110.575 28.095 110.745 28.555 ;
      RECT 110.575 28.095 111.24 28.265 ;
      RECT 111.01 26.935 111.24 28.265 ;
      RECT 110.575 26.935 111.24 27.105 ;
      RECT 110.575 26.435 110.745 27.105 ;
      RECT 109.59 21.425 111.225 21.665 ;
      RECT 110.995 21.335 111.225 21.665 ;
      RECT 109.59 20.995 109.84 21.665 ;
      RECT 110.54 22.185 110.82 22.785 ;
      RECT 110.54 22.185 111.015 22.385 ;
      RECT 109.515 31.09 110.62 31.26 ;
      RECT 110.45 30.215 110.62 31.26 ;
      RECT 110.45 30.215 110.96 30.475 ;
      RECT 110.79 30.145 110.96 30.475 ;
      RECT 110.09 30.215 110.96 30.385 ;
      RECT 110.09 29.265 110.26 30.385 ;
      RECT 109.585 29.265 110.26 29.435 ;
      RECT 110.115 19.815 110.285 20.485 ;
      RECT 110.115 19.815 110.78 19.985 ;
      RECT 110.55 18.655 110.78 19.985 ;
      RECT 110.115 18.655 110.78 18.825 ;
      RECT 110.115 18.365 110.285 18.825 ;
      RECT 110.395 17.195 110.725 17.715 ;
      RECT 110.605 16.445 110.775 17.28 ;
      RECT 110.55 17.155 110.775 17.28 ;
      RECT 110.56 16.445 110.775 16.575 ;
      RECT 110.385 15.6 110.715 16.525 ;
      RECT 109.555 17.195 109.885 17.72 ;
      RECT 109.685 16.695 109.885 17.72 ;
      RECT 109.685 16.695 110.435 17.025 ;
      RECT 109.685 15.555 109.875 17.72 ;
      RECT 108.98 16.115 109.875 16.49 ;
      RECT 109.535 15.555 109.875 16.49 ;
      RECT 109.75 30.555 110.28 30.92 ;
      RECT 109.75 29.635 109.92 30.92 ;
      RECT 109.395 29.635 109.92 29.855 ;
      RECT 109.985 22.185 110.27 22.785 ;
      RECT 109.94 22.185 110.27 22.385 ;
      RECT 109.405 22.185 109.77 22.385 ;
      RECT 109.395 22.185 109.77 22.355 ;
      RECT 108.025 17.485 108.81 17.655 ;
      RECT 108.64 15.685 108.81 17.655 ;
      RECT 108.64 16.695 109.515 17.025 ;
      RECT 107.925 15.685 108.81 15.855 ;
      RECT 109.055 30.81 109.305 31.365 ;
      RECT 109 29.575 109.17 30.94 ;
      RECT 109.055 29.265 109.225 29.705 ;
      RECT 109.055 29.265 109.39 29.435 ;
      RECT 108.665 22.875 108.92 23.205 ;
      RECT 108.665 22.865 108.875 23.205 ;
      RECT 108.665 22.795 108.85 23.205 ;
      RECT 108.665 20.995 108.835 23.205 ;
      RECT 108.665 20.995 108.92 21.665 ;
      RECT 108.005 16.985 108.47 17.315 ;
      RECT 108.15 16.025 108.47 17.315 ;
      RECT 108.215 19.475 108.385 20.485 ;
      RECT 105.325 19.475 108.385 19.645 ;
      RECT 105.325 18.755 105.495 19.645 ;
      RECT 107.32 18.755 108.385 18.925 ;
      RECT 108.215 18.275 108.385 18.925 ;
      RECT 105.325 18.755 106.125 18.925 ;
      RECT 105.955 18.275 106.125 18.925 ;
      RECT 107.32 18.275 107.49 18.925 ;
      RECT 105.955 18.275 107.49 18.525 ;
      RECT 106.875 20.315 108.045 20.485 ;
      RECT 107.715 19.815 108.045 20.485 ;
      RECT 106.875 20.275 107.205 20.485 ;
      RECT 107.355 30.695 107.525 31.365 ;
      RECT 107.355 30.695 108.02 30.865 ;
      RECT 107.79 29.535 108.02 30.865 ;
      RECT 107.355 29.535 108.02 29.705 ;
      RECT 107.355 29.245 107.525 29.705 ;
      RECT 107.45 17.485 107.855 17.655 ;
      RECT 107.45 15.555 107.62 17.655 ;
      RECT 106.79 16.955 107.62 17.255 ;
      RECT 106.79 16.925 106.99 17.255 ;
      RECT 107.45 15.555 107.7 15.885 ;
      RECT 103.675 11.675 103.845 12.325 ;
      RECT 104.515 11.675 104.685 12.32 ;
      RECT 103.675 11.675 105.095 11.845 ;
      RECT 104.92 10.965 105.095 11.845 ;
      RECT 104.92 11.335 107.545 11.505 ;
      RECT 103.595 10.965 105.095 11.135 ;
      RECT 104.435 10.115 104.765 11.135 ;
      RECT 103.595 10.115 103.925 11.135 ;
      RECT 105.91 19.815 106.16 20.485 ;
      RECT 107.315 19.815 107.545 20.145 ;
      RECT 105.91 19.815 107.545 20.055 ;
      RECT 106.86 19.095 107.335 19.295 ;
      RECT 106.86 18.695 107.14 19.295 ;
      RECT 105.905 17.485 106.58 17.655 ;
      RECT 106.41 16.535 106.58 17.655 ;
      RECT 107.11 16.445 107.28 16.775 ;
      RECT 106.41 16.535 107.28 16.705 ;
      RECT 106.77 16.445 107.28 16.705 ;
      RECT 106.77 15.66 106.94 16.705 ;
      RECT 105.835 15.66 106.94 15.83 ;
      RECT 105.715 17.065 106.24 17.285 ;
      RECT 106.07 16 106.24 17.285 ;
      RECT 106.07 16 106.6 16.365 ;
      RECT 106.26 19.095 106.59 19.295 ;
      RECT 106.305 18.695 106.59 19.295 ;
      RECT 105.715 19.125 106.09 19.295 ;
      RECT 105.725 19.095 106.09 19.295 ;
      RECT 105.375 17.485 105.71 17.655 ;
      RECT 105.375 17.215 105.545 17.655 ;
      RECT 105.32 15.98 105.49 17.345 ;
      RECT 105.375 15.555 105.625 16.11 ;
      RECT 104.985 19.815 105.24 20.485 ;
      RECT 104.985 18.275 105.155 20.485 ;
      RECT 104.985 18.275 105.17 18.685 ;
      RECT 104.985 18.275 105.195 18.615 ;
      RECT 104.985 18.275 105.24 18.605 ;
      RECT 103.675 17.215 103.845 17.675 ;
      RECT 103.675 17.215 104.34 17.385 ;
      RECT 104.11 16.055 104.34 17.385 ;
      RECT 103.675 16.055 104.34 16.225 ;
      RECT 103.675 15.555 103.845 16.225 ;
      RECT 100.735 17.195 101.065 17.715 ;
      RECT 100.945 16.445 101.115 17.28 ;
      RECT 100.89 17.155 101.115 17.28 ;
      RECT 100.9 16.445 101.115 16.575 ;
      RECT 100.725 15.6 101.055 16.525 ;
      RECT 97.235 11.675 97.405 12.325 ;
      RECT 98.075 11.675 98.245 12.32 ;
      RECT 97.235 11.675 98.655 11.845 ;
      RECT 98.48 10.965 98.655 11.845 ;
      RECT 98.48 11.335 101.105 11.505 ;
      RECT 97.155 10.965 98.655 11.135 ;
      RECT 97.995 10.115 98.325 11.135 ;
      RECT 97.155 10.115 97.485 11.135 ;
      RECT 99.895 17.195 100.225 17.72 ;
      RECT 100.025 16.695 100.225 17.72 ;
      RECT 100.025 16.695 100.775 17.025 ;
      RECT 100.025 15.555 100.215 17.72 ;
      RECT 99.32 16.115 100.215 16.49 ;
      RECT 99.875 15.555 100.215 16.49 ;
      RECT 100.275 22.635 100.605 23.155 ;
      RECT 100.485 21.885 100.655 22.72 ;
      RECT 100.43 22.595 100.655 22.72 ;
      RECT 100.44 21.885 100.655 22.015 ;
      RECT 100.265 21.04 100.595 21.965 ;
      RECT 99.435 22.635 99.765 23.16 ;
      RECT 99.565 22.135 99.765 23.16 ;
      RECT 99.565 22.135 100.315 22.465 ;
      RECT 99.565 20.995 99.755 23.16 ;
      RECT 98.86 21.555 99.755 21.93 ;
      RECT 99.415 20.995 99.755 21.93 ;
      RECT 99.805 35.835 100.135 36.76 ;
      RECT 100.025 35.08 100.195 35.915 ;
      RECT 99.98 35.785 100.195 35.915 ;
      RECT 99.97 35.08 100.195 35.205 ;
      RECT 99.815 34.645 100.145 35.165 ;
      RECT 98.365 17.485 99.15 17.655 ;
      RECT 98.98 15.685 99.15 17.655 ;
      RECT 98.98 16.695 99.855 17.025 ;
      RECT 98.265 15.685 99.15 15.855 ;
      RECT 98.955 35.87 99.295 36.805 ;
      RECT 99.105 34.64 99.295 36.805 ;
      RECT 98.4 35.87 99.295 36.245 ;
      RECT 99.105 35.335 99.855 35.665 ;
      RECT 99.105 34.64 99.305 35.665 ;
      RECT 98.975 34.64 99.305 35.165 ;
      RECT 97.905 22.925 98.69 23.095 ;
      RECT 98.52 21.125 98.69 23.095 ;
      RECT 98.52 22.135 99.395 22.465 ;
      RECT 97.805 21.125 98.69 21.295 ;
      RECT 97.345 36.505 98.23 36.675 ;
      RECT 98.06 34.705 98.23 36.675 ;
      RECT 98.06 35.335 98.935 35.665 ;
      RECT 97.445 34.705 98.23 34.875 ;
      RECT 98.345 16.985 98.81 17.315 ;
      RECT 98.49 16.025 98.81 17.315 ;
      RECT 97.885 22.425 98.35 22.755 ;
      RECT 98.03 21.465 98.35 22.755 ;
      RECT 98.08 19.815 98.335 20.485 ;
      RECT 98.165 18.275 98.335 20.485 ;
      RECT 98.15 18.275 98.335 18.685 ;
      RECT 98.125 18.275 98.335 18.615 ;
      RECT 98.08 18.275 98.335 18.605 ;
      RECT 98.08 25.255 98.335 25.925 ;
      RECT 98.165 23.715 98.335 25.925 ;
      RECT 98.15 23.715 98.335 24.125 ;
      RECT 98.125 23.715 98.335 24.055 ;
      RECT 98.08 23.715 98.335 24.045 ;
      RECT 98.08 33.755 98.335 34.085 ;
      RECT 98.165 31.875 98.335 34.085 ;
      RECT 98.125 33.745 98.335 34.085 ;
      RECT 98.15 33.675 98.335 34.085 ;
      RECT 98.08 31.875 98.335 32.545 ;
      RECT 97.79 17.485 98.195 17.655 ;
      RECT 97.79 15.555 97.96 17.655 ;
      RECT 97.13 16.955 97.96 17.255 ;
      RECT 97.13 16.925 97.33 17.255 ;
      RECT 97.79 15.555 98.04 15.885 ;
      RECT 94.935 19.475 95.105 20.485 ;
      RECT 94.935 19.475 97.995 19.645 ;
      RECT 97.825 18.755 97.995 19.645 ;
      RECT 97.195 18.755 97.995 18.925 ;
      RECT 94.935 18.755 96 18.925 ;
      RECT 95.83 18.275 96 18.925 ;
      RECT 97.195 18.275 97.365 18.925 ;
      RECT 94.935 18.275 95.105 18.925 ;
      RECT 95.83 18.275 97.365 18.525 ;
      RECT 94.935 24.915 95.105 25.925 ;
      RECT 94.935 24.915 97.995 25.085 ;
      RECT 97.825 24.195 97.995 25.085 ;
      RECT 97.195 24.195 97.995 24.365 ;
      RECT 94.935 24.195 96 24.365 ;
      RECT 95.83 23.715 96 24.365 ;
      RECT 97.195 23.715 97.365 24.365 ;
      RECT 94.935 23.715 95.105 24.365 ;
      RECT 95.83 23.715 97.365 23.965 ;
      RECT 95.83 33.835 97.365 34.085 ;
      RECT 97.195 33.435 97.365 34.085 ;
      RECT 94.935 33.435 95.105 34.085 ;
      RECT 95.83 33.435 96 34.085 ;
      RECT 97.195 33.435 97.995 33.605 ;
      RECT 97.825 32.715 97.995 33.605 ;
      RECT 94.935 33.435 96 33.605 ;
      RECT 94.935 32.715 97.995 32.885 ;
      RECT 94.935 31.875 95.105 32.885 ;
      RECT 97.57 35.045 97.89 36.335 ;
      RECT 97.425 35.045 97.89 35.375 ;
      RECT 97.33 22.925 97.735 23.095 ;
      RECT 97.33 20.995 97.5 23.095 ;
      RECT 96.67 22.395 97.5 22.695 ;
      RECT 96.67 22.365 96.87 22.695 ;
      RECT 97.33 20.995 97.58 21.325 ;
      RECT 96.245 17.485 96.92 17.655 ;
      RECT 96.75 16.535 96.92 17.655 ;
      RECT 97.45 16.445 97.62 16.775 ;
      RECT 96.75 16.535 97.62 16.705 ;
      RECT 97.11 16.445 97.62 16.705 ;
      RECT 97.11 15.66 97.28 16.705 ;
      RECT 96.175 15.66 97.28 15.83 ;
      RECT 97.23 19.125 97.605 19.295 ;
      RECT 97.23 19.095 97.595 19.295 ;
      RECT 97.23 24.565 97.605 24.735 ;
      RECT 97.23 24.535 97.595 24.735 ;
      RECT 97.23 33.065 97.595 33.265 ;
      RECT 97.23 33.065 97.605 33.235 ;
      RECT 97.16 19.815 97.41 20.485 ;
      RECT 95.775 19.815 96.005 20.145 ;
      RECT 95.775 19.815 97.41 20.055 ;
      RECT 97.16 25.255 97.41 25.925 ;
      RECT 95.775 25.255 96.005 25.585 ;
      RECT 95.775 25.255 97.41 25.495 ;
      RECT 95.775 32.305 97.41 32.545 ;
      RECT 97.16 31.875 97.41 32.545 ;
      RECT 95.775 32.215 96.005 32.545 ;
      RECT 96.87 36.475 97.12 36.805 ;
      RECT 96.87 34.705 97.04 36.805 ;
      RECT 96.21 35.105 96.41 35.435 ;
      RECT 96.21 35.105 97.04 35.405 ;
      RECT 96.87 34.705 97.275 34.875 ;
      RECT 95.785 22.925 96.46 23.095 ;
      RECT 96.29 21.975 96.46 23.095 ;
      RECT 96.99 21.885 97.16 22.215 ;
      RECT 96.29 21.975 97.16 22.145 ;
      RECT 96.65 21.885 97.16 22.145 ;
      RECT 96.65 21.1 96.82 22.145 ;
      RECT 95.715 21.1 96.82 21.27 ;
      RECT 96.73 19.095 97.06 19.295 ;
      RECT 96.73 18.695 97.015 19.295 ;
      RECT 96.73 24.535 97.06 24.735 ;
      RECT 96.73 24.135 97.015 24.735 ;
      RECT 96.73 33.065 97.015 33.665 ;
      RECT 96.73 33.065 97.06 33.265 ;
      RECT 96.055 17.065 96.58 17.285 ;
      RECT 96.41 16 96.58 17.285 ;
      RECT 96.41 16 96.94 16.365 ;
      RECT 95.255 36.53 96.36 36.7 ;
      RECT 96.19 35.655 96.36 36.7 ;
      RECT 96.19 35.655 96.7 35.915 ;
      RECT 96.53 35.585 96.7 35.915 ;
      RECT 95.83 35.655 96.7 35.825 ;
      RECT 95.83 34.705 96 35.825 ;
      RECT 95.325 34.705 96 34.875 ;
      RECT 95.595 22.505 96.12 22.725 ;
      RECT 95.95 21.44 96.12 22.725 ;
      RECT 95.95 21.44 96.48 21.805 ;
      RECT 95.985 19.095 96.46 19.295 ;
      RECT 96.18 18.695 96.46 19.295 ;
      RECT 95.985 24.535 96.46 24.735 ;
      RECT 96.18 24.135 96.46 24.735 ;
      RECT 96.18 33.065 96.46 33.665 ;
      RECT 95.985 33.065 96.46 33.265 ;
      RECT 95.275 20.315 96.445 20.485 ;
      RECT 96.115 20.275 96.445 20.485 ;
      RECT 95.275 19.815 95.605 20.485 ;
      RECT 95.275 25.755 96.445 25.925 ;
      RECT 96.115 25.715 96.445 25.925 ;
      RECT 95.275 25.255 95.605 25.925 ;
      RECT 95.275 31.875 95.605 32.545 ;
      RECT 96.115 31.875 96.445 32.085 ;
      RECT 95.275 31.875 96.445 32.045 ;
      RECT 95.715 17.485 96.05 17.655 ;
      RECT 95.715 17.215 95.885 17.655 ;
      RECT 95.66 15.98 95.83 17.345 ;
      RECT 95.715 15.555 95.965 16.11 ;
      RECT 95.49 35.995 96.02 36.36 ;
      RECT 95.49 35.075 95.66 36.36 ;
      RECT 95.135 35.075 95.66 35.295 ;
      RECT 95.255 22.925 95.59 23.095 ;
      RECT 95.255 22.655 95.425 23.095 ;
      RECT 95.2 21.42 95.37 22.785 ;
      RECT 95.255 20.995 95.505 21.55 ;
      RECT 94.795 36.25 95.045 36.805 ;
      RECT 94.74 35.015 94.91 36.38 ;
      RECT 94.795 34.705 94.965 35.145 ;
      RECT 94.795 34.705 95.13 34.875 ;
      RECT 94.015 17.215 94.185 17.675 ;
      RECT 94.015 17.215 94.68 17.385 ;
      RECT 94.45 16.055 94.68 17.385 ;
      RECT 94.015 16.055 94.68 16.225 ;
      RECT 94.015 15.555 94.185 16.225 ;
      RECT 90.795 11.675 90.965 12.325 ;
      RECT 91.635 11.675 91.805 12.32 ;
      RECT 90.795 11.675 92.215 11.845 ;
      RECT 92.04 10.965 92.215 11.845 ;
      RECT 92.04 11.335 94.665 11.505 ;
      RECT 90.715 10.965 92.215 11.135 ;
      RECT 91.555 10.115 91.885 11.135 ;
      RECT 90.715 10.115 91.045 11.135 ;
      RECT 93.555 22.655 93.725 23.115 ;
      RECT 93.555 22.655 94.22 22.825 ;
      RECT 93.99 21.495 94.22 22.825 ;
      RECT 93.555 21.495 94.22 21.665 ;
      RECT 93.555 20.995 93.725 21.665 ;
      RECT 93.095 36.135 93.265 36.805 ;
      RECT 93.095 36.135 93.76 36.305 ;
      RECT 93.53 34.975 93.76 36.305 ;
      RECT 93.095 34.975 93.76 35.145 ;
      RECT 93.095 34.685 93.265 35.145 ;
      RECT 87.855 17.195 88.185 17.715 ;
      RECT 88.065 16.445 88.235 17.28 ;
      RECT 88.01 17.155 88.235 17.28 ;
      RECT 88.02 16.445 88.235 16.575 ;
      RECT 87.845 15.6 88.175 16.525 ;
      RECT 87.015 17.195 87.345 17.72 ;
      RECT 87.145 16.695 87.345 17.72 ;
      RECT 87.145 16.695 87.895 17.025 ;
      RECT 87.145 15.555 87.335 17.72 ;
      RECT 86.44 16.115 87.335 16.49 ;
      RECT 86.995 15.555 87.335 16.49 ;
      RECT 87.515 22.555 87.685 23.205 ;
      RECT 86.675 22.555 86.845 23.2 ;
      RECT 86.265 22.555 87.685 22.725 ;
      RECT 86.265 21.845 86.44 22.725 ;
      RECT 83.815 22.215 86.44 22.385 ;
      RECT 86.265 21.845 87.765 22.015 ;
      RECT 87.435 20.995 87.765 22.015 ;
      RECT 86.595 20.995 86.925 22.015 ;
      RECT 85.485 17.485 86.27 17.655 ;
      RECT 86.1 15.685 86.27 17.655 ;
      RECT 86.1 16.695 86.975 17.025 ;
      RECT 85.385 15.685 86.27 15.855 ;
      RECT 82.975 11.675 83.145 12.325 ;
      RECT 83.815 11.675 83.985 12.32 ;
      RECT 82.975 11.675 84.395 11.845 ;
      RECT 84.22 10.965 84.395 11.845 ;
      RECT 84.22 11.335 86.845 11.505 ;
      RECT 82.895 10.965 84.395 11.135 ;
      RECT 83.735 10.115 84.065 11.135 ;
      RECT 82.895 10.115 83.225 11.135 ;
      RECT 86.595 19.475 86.765 20.485 ;
      RECT 83.705 19.475 86.765 19.645 ;
      RECT 83.705 18.755 83.875 19.645 ;
      RECT 85.7 18.755 86.765 18.925 ;
      RECT 86.595 18.275 86.765 18.925 ;
      RECT 83.705 18.755 84.505 18.925 ;
      RECT 84.335 18.275 84.505 18.925 ;
      RECT 85.7 18.275 85.87 18.925 ;
      RECT 84.335 18.275 85.87 18.525 ;
      RECT 85.255 20.315 86.425 20.485 ;
      RECT 86.095 19.815 86.425 20.485 ;
      RECT 85.255 20.275 85.585 20.485 ;
      RECT 85.465 16.985 85.93 17.315 ;
      RECT 85.61 16.025 85.93 17.315 ;
      RECT 84.29 19.815 84.54 20.485 ;
      RECT 85.695 19.815 85.925 20.145 ;
      RECT 84.29 19.815 85.925 20.055 ;
      RECT 85.24 19.095 85.715 19.295 ;
      RECT 85.24 18.695 85.52 19.295 ;
      RECT 85.215 24.915 85.385 25.925 ;
      RECT 82.325 24.915 85.385 25.085 ;
      RECT 82.325 24.195 82.495 25.085 ;
      RECT 84.32 24.195 85.385 24.365 ;
      RECT 85.215 23.715 85.385 24.365 ;
      RECT 82.325 24.195 83.125 24.365 ;
      RECT 82.955 23.715 83.125 24.365 ;
      RECT 84.32 23.715 84.49 24.365 ;
      RECT 82.955 23.715 84.49 23.965 ;
      RECT 84.91 17.485 85.315 17.655 ;
      RECT 84.91 15.555 85.08 17.655 ;
      RECT 84.25 16.955 85.08 17.255 ;
      RECT 84.25 16.925 84.45 17.255 ;
      RECT 84.91 15.555 85.16 15.885 ;
      RECT 83.875 25.755 85.045 25.925 ;
      RECT 84.715 25.255 85.045 25.925 ;
      RECT 83.875 25.715 84.205 25.925 ;
      RECT 84.635 28.075 84.965 28.595 ;
      RECT 84.845 27.325 85.015 28.16 ;
      RECT 84.79 28.035 85.015 28.16 ;
      RECT 84.8 27.325 85.015 27.455 ;
      RECT 84.625 26.48 84.955 27.405 ;
      RECT 84.64 19.095 84.97 19.295 ;
      RECT 84.685 18.695 84.97 19.295 ;
      RECT 83.365 17.485 84.04 17.655 ;
      RECT 83.87 16.535 84.04 17.655 ;
      RECT 84.57 16.445 84.74 16.775 ;
      RECT 83.87 16.535 84.74 16.705 ;
      RECT 84.23 16.445 84.74 16.705 ;
      RECT 84.23 15.66 84.4 16.705 ;
      RECT 83.295 15.66 84.4 15.83 ;
      RECT 83.795 28.075 84.125 28.6 ;
      RECT 83.925 27.575 84.125 28.6 ;
      RECT 83.925 27.575 84.675 27.905 ;
      RECT 83.925 26.435 84.115 28.6 ;
      RECT 83.22 26.995 84.115 27.37 ;
      RECT 83.775 26.435 84.115 27.37 ;
      RECT 82.91 25.255 83.16 25.925 ;
      RECT 84.315 25.255 84.545 25.585 ;
      RECT 82.91 25.255 84.545 25.495 ;
      RECT 84.095 19.125 84.47 19.295 ;
      RECT 84.105 19.095 84.47 19.295 ;
      RECT 83.86 24.535 84.335 24.735 ;
      RECT 83.86 24.135 84.14 24.735 ;
      RECT 83.175 17.065 83.7 17.285 ;
      RECT 83.53 16 83.7 17.285 ;
      RECT 83.53 16 84.06 16.365 ;
      RECT 82.265 28.365 83.05 28.535 ;
      RECT 82.88 26.565 83.05 28.535 ;
      RECT 82.88 27.575 83.755 27.905 ;
      RECT 82.165 26.565 83.05 26.735 ;
      RECT 83.365 19.815 83.62 20.485 ;
      RECT 83.365 19.805 83.575 20.485 ;
      RECT 83.365 18.275 83.535 20.485 ;
      RECT 83.365 18.275 83.55 18.685 ;
      RECT 83.365 18.275 83.62 18.605 ;
      RECT 83.26 24.535 83.59 24.735 ;
      RECT 83.305 24.135 83.59 24.735 ;
      RECT 82.835 17.485 83.17 17.655 ;
      RECT 82.835 17.215 83.005 17.655 ;
      RECT 82.78 15.98 82.95 17.345 ;
      RECT 82.835 15.555 83.085 16.11 ;
      RECT 82.715 24.565 83.09 24.735 ;
      RECT 82.725 24.535 83.09 24.735 ;
      RECT 82.245 27.865 82.71 28.195 ;
      RECT 82.39 26.905 82.71 28.195 ;
      RECT 81.875 33.515 82.205 34.035 ;
      RECT 82.085 32.765 82.255 33.6 ;
      RECT 82.03 33.475 82.255 33.6 ;
      RECT 82.04 32.765 82.255 32.895 ;
      RECT 81.865 31.92 82.195 32.845 ;
      RECT 81.985 25.255 82.24 25.925 ;
      RECT 81.985 23.715 82.155 25.925 ;
      RECT 81.985 23.715 82.17 24.125 ;
      RECT 81.985 23.715 82.24 24.045 ;
      RECT 81.69 28.365 82.095 28.535 ;
      RECT 81.69 26.435 81.86 28.535 ;
      RECT 81.03 27.835 81.86 28.135 ;
      RECT 81.03 27.805 81.23 28.135 ;
      RECT 81.69 26.435 81.94 26.765 ;
      RECT 81.035 33.515 81.365 34.04 ;
      RECT 81.165 33.015 81.365 34.04 ;
      RECT 81.165 33.015 81.915 33.345 ;
      RECT 81.165 31.875 81.355 34.04 ;
      RECT 80.46 32.435 81.355 32.81 ;
      RECT 81.015 31.875 81.355 32.81 ;
      RECT 81.135 17.215 81.305 17.675 ;
      RECT 81.135 17.215 81.8 17.385 ;
      RECT 81.57 16.055 81.8 17.385 ;
      RECT 81.135 16.055 81.8 16.225 ;
      RECT 81.135 15.555 81.305 16.225 ;
      RECT 80.145 28.365 80.82 28.535 ;
      RECT 80.65 27.415 80.82 28.535 ;
      RECT 81.35 27.325 81.52 27.655 ;
      RECT 80.65 27.415 81.52 27.585 ;
      RECT 81.01 27.325 81.52 27.585 ;
      RECT 81.01 26.54 81.18 27.585 ;
      RECT 80.075 26.54 81.18 26.71 ;
      RECT 80.945 19.515 81.275 20.44 ;
      RECT 81.165 18.76 81.335 19.595 ;
      RECT 81.12 19.465 81.335 19.595 ;
      RECT 81.11 18.76 81.335 18.885 ;
      RECT 80.955 18.325 81.285 18.845 ;
      RECT 77.455 11.675 77.625 12.325 ;
      RECT 78.295 11.675 78.465 12.32 ;
      RECT 77.455 11.675 78.875 11.845 ;
      RECT 78.7 10.965 78.875 11.845 ;
      RECT 78.7 11.335 81.325 11.505 ;
      RECT 77.375 10.965 78.875 11.135 ;
      RECT 78.215 10.115 78.545 11.135 ;
      RECT 77.375 10.115 77.705 11.135 ;
      RECT 80.095 19.55 80.435 20.485 ;
      RECT 80.245 18.32 80.435 20.485 ;
      RECT 79.54 19.55 80.435 19.925 ;
      RECT 80.245 19.015 80.995 19.345 ;
      RECT 80.245 18.32 80.445 19.345 ;
      RECT 80.115 18.32 80.445 18.845 ;
      RECT 79.505 33.805 80.29 33.975 ;
      RECT 80.12 32.005 80.29 33.975 ;
      RECT 80.12 33.015 80.995 33.345 ;
      RECT 79.405 32.005 80.29 32.175 ;
      RECT 79.955 27.945 80.48 28.165 ;
      RECT 80.31 26.88 80.48 28.165 ;
      RECT 80.31 26.88 80.84 27.245 ;
      RECT 78.485 20.185 79.37 20.355 ;
      RECT 79.2 18.385 79.37 20.355 ;
      RECT 79.2 19.015 80.075 19.345 ;
      RECT 78.585 18.385 79.37 18.555 ;
      RECT 79.615 28.365 79.95 28.535 ;
      RECT 79.615 28.095 79.785 28.535 ;
      RECT 79.56 26.86 79.73 28.225 ;
      RECT 79.615 26.435 79.865 26.99 ;
      RECT 79.485 33.305 79.95 33.635 ;
      RECT 79.63 32.345 79.95 33.635 ;
      RECT 78.93 33.805 79.335 33.975 ;
      RECT 78.93 31.875 79.1 33.975 ;
      RECT 78.27 33.275 79.1 33.575 ;
      RECT 78.27 33.245 78.47 33.575 ;
      RECT 78.93 31.875 79.18 32.205 ;
      RECT 78.71 18.725 79.03 20.015 ;
      RECT 78.565 18.725 79.03 19.055 ;
      RECT 78.775 24.915 78.945 25.925 ;
      RECT 75.885 24.915 78.945 25.085 ;
      RECT 75.885 24.195 76.055 25.085 ;
      RECT 77.88 24.195 78.945 24.365 ;
      RECT 78.775 23.715 78.945 24.365 ;
      RECT 75.885 24.195 76.685 24.365 ;
      RECT 76.515 23.715 76.685 24.365 ;
      RECT 77.88 23.715 78.05 24.365 ;
      RECT 76.515 23.715 78.05 23.965 ;
      RECT 77.385 33.805 78.06 33.975 ;
      RECT 77.89 32.855 78.06 33.975 ;
      RECT 78.59 32.765 78.76 33.095 ;
      RECT 77.89 32.855 78.76 33.025 ;
      RECT 78.25 32.765 78.76 33.025 ;
      RECT 78.25 31.98 78.42 33.025 ;
      RECT 77.315 31.98 78.42 32.15 ;
      RECT 77.435 25.755 78.605 25.925 ;
      RECT 78.275 25.255 78.605 25.925 ;
      RECT 77.435 25.715 77.765 25.925 ;
      RECT 77.915 28.095 78.085 28.555 ;
      RECT 77.915 28.095 78.58 28.265 ;
      RECT 78.35 26.935 78.58 28.265 ;
      RECT 77.915 26.935 78.58 27.105 ;
      RECT 77.915 26.435 78.085 27.105 ;
      RECT 78.01 20.155 78.26 20.485 ;
      RECT 78.01 18.385 78.18 20.485 ;
      RECT 77.35 18.785 77.55 19.115 ;
      RECT 77.35 18.785 78.18 19.085 ;
      RECT 78.01 18.385 78.415 18.555 ;
      RECT 76.47 25.255 76.72 25.925 ;
      RECT 77.875 25.255 78.105 25.585 ;
      RECT 76.47 25.255 78.105 25.495 ;
      RECT 77.195 33.385 77.72 33.605 ;
      RECT 77.55 32.32 77.72 33.605 ;
      RECT 77.55 32.32 78.08 32.685 ;
      RECT 77.42 24.535 77.895 24.735 ;
      RECT 77.42 24.135 77.7 24.735 ;
      RECT 76.395 20.21 77.5 20.38 ;
      RECT 77.33 19.335 77.5 20.38 ;
      RECT 77.33 19.335 77.84 19.595 ;
      RECT 77.67 19.265 77.84 19.595 ;
      RECT 76.97 19.335 77.84 19.505 ;
      RECT 76.97 18.385 77.14 19.505 ;
      RECT 76.465 18.385 77.14 18.555 ;
      RECT 76.855 33.805 77.19 33.975 ;
      RECT 76.855 33.535 77.025 33.975 ;
      RECT 76.8 32.3 76.97 33.665 ;
      RECT 76.855 31.875 77.105 32.43 ;
      RECT 76.63 19.675 77.16 20.04 ;
      RECT 76.63 18.755 76.8 20.04 ;
      RECT 76.275 18.755 76.8 18.975 ;
      RECT 76.82 24.535 77.15 24.735 ;
      RECT 76.865 24.135 77.15 24.735 ;
      RECT 75.935 19.93 76.185 20.485 ;
      RECT 75.88 18.695 76.05 20.06 ;
      RECT 75.935 18.385 76.105 18.825 ;
      RECT 75.935 18.385 76.27 18.555 ;
      RECT 75.155 33.535 75.325 33.995 ;
      RECT 75.155 33.535 75.82 33.705 ;
      RECT 75.59 32.375 75.82 33.705 ;
      RECT 75.155 32.375 75.82 32.545 ;
      RECT 75.155 31.875 75.325 32.545 ;
      RECT 75.545 25.255 75.8 25.925 ;
      RECT 75.545 23.715 75.715 25.925 ;
      RECT 75.545 23.715 75.73 24.125 ;
      RECT 75.545 23.715 75.8 24.045 ;
      RECT 74.235 19.815 74.405 20.485 ;
      RECT 74.235 19.815 74.9 19.985 ;
      RECT 74.67 18.655 74.9 19.985 ;
      RECT 74.235 18.655 74.9 18.825 ;
      RECT 74.235 18.365 74.405 18.825 ;
      RECT 72.7 19.48 72.96 20.455 ;
      RECT 71.845 19.48 72.1 20.455 ;
      RECT 70.985 19.48 71.24 20.455 ;
      RECT 70.485 19.48 73.515 19.65 ;
      RECT 73.215 18.745 73.515 19.65 ;
      RECT 74.15 18.995 74.5 19.645 ;
      RECT 70.485 18.745 70.655 19.65 ;
      RECT 73.215 19.125 74.5 19.295 ;
      RECT 70.485 18.745 73.515 18.915 ;
      RECT 72.27 18.3 72.525 18.915 ;
      RECT 71.41 18.3 71.67 18.915 ;
      RECT 73.135 17.195 73.465 17.715 ;
      RECT 73.345 16.445 73.515 17.28 ;
      RECT 73.29 17.155 73.515 17.28 ;
      RECT 73.345 16.745 73.915 16.915 ;
      RECT 73.3 16.445 73.515 16.575 ;
      RECT 73.125 15.6 73.455 16.525 ;
      RECT 72.295 17.195 72.625 17.72 ;
      RECT 72.425 16.695 72.625 17.72 ;
      RECT 72.425 16.695 73.175 17.025 ;
      RECT 72.425 15.555 72.615 17.72 ;
      RECT 71.72 16.115 72.615 16.49 ;
      RECT 72.275 15.555 72.615 16.49 ;
      RECT 70.765 17.485 71.55 17.655 ;
      RECT 71.38 15.685 71.55 17.655 ;
      RECT 71.38 16.695 72.255 17.025 ;
      RECT 70.665 15.685 71.55 15.855 ;
      RECT 68.255 11.675 68.425 12.325 ;
      RECT 69.095 11.675 69.265 12.32 ;
      RECT 68.255 11.675 69.675 11.845 ;
      RECT 69.5 10.965 69.675 11.845 ;
      RECT 69.5 11.335 72.125 11.505 ;
      RECT 68.175 10.965 69.675 11.135 ;
      RECT 69.015 10.115 69.345 11.135 ;
      RECT 68.175 10.115 68.505 11.135 ;
      RECT 70.835 28.075 71.165 28.595 ;
      RECT 71.045 27.325 71.215 28.16 ;
      RECT 70.99 28.035 71.215 28.16 ;
      RECT 71 27.325 71.215 27.455 ;
      RECT 70.825 26.48 71.155 27.405 ;
      RECT 70.745 16.985 71.21 17.315 ;
      RECT 70.89 16.025 71.21 17.315 ;
      RECT 69.995 28.075 70.325 28.6 ;
      RECT 70.125 27.575 70.325 28.6 ;
      RECT 70.125 27.575 70.875 27.905 ;
      RECT 70.125 26.435 70.315 28.6 ;
      RECT 69.42 26.995 70.315 27.37 ;
      RECT 69.975 26.435 70.315 27.37 ;
      RECT 70.495 24.915 70.665 25.925 ;
      RECT 67.605 24.915 70.665 25.085 ;
      RECT 67.605 24.195 67.775 25.085 ;
      RECT 69.6 24.195 70.665 24.365 ;
      RECT 70.495 23.715 70.665 24.365 ;
      RECT 67.605 24.195 68.405 24.365 ;
      RECT 68.235 23.715 68.405 24.365 ;
      RECT 69.6 23.715 69.77 24.365 ;
      RECT 68.235 23.715 69.77 23.965 ;
      RECT 70.19 17.485 70.595 17.655 ;
      RECT 70.19 15.555 70.36 17.655 ;
      RECT 69.53 16.955 70.36 17.255 ;
      RECT 69.53 16.925 69.73 17.255 ;
      RECT 70.19 15.555 70.44 15.885 ;
      RECT 69.155 25.755 70.325 25.925 ;
      RECT 69.995 25.255 70.325 25.925 ;
      RECT 69.155 25.715 69.485 25.925 ;
      RECT 68.645 17.485 69.32 17.655 ;
      RECT 69.15 16.535 69.32 17.655 ;
      RECT 69.85 16.445 70.02 16.775 ;
      RECT 69.15 16.535 70.02 16.705 ;
      RECT 69.51 16.445 70.02 16.705 ;
      RECT 69.51 15.66 69.68 16.705 ;
      RECT 68.575 15.66 69.68 15.83 ;
      RECT 68.465 28.365 69.25 28.535 ;
      RECT 69.08 26.565 69.25 28.535 ;
      RECT 69.08 27.575 69.955 27.905 ;
      RECT 68.365 26.565 69.25 26.735 ;
      RECT 68.19 25.255 68.44 25.925 ;
      RECT 69.595 25.255 69.825 25.585 ;
      RECT 68.19 25.255 69.825 25.495 ;
      RECT 65.955 38.875 66.125 39.525 ;
      RECT 66.795 38.875 66.965 39.52 ;
      RECT 65.955 38.875 67.375 39.045 ;
      RECT 67.2 38.165 67.375 39.045 ;
      RECT 67.2 38.535 69.825 38.705 ;
      RECT 65.875 38.165 67.375 38.335 ;
      RECT 66.715 37.315 67.045 38.335 ;
      RECT 65.875 37.315 66.205 38.335 ;
      RECT 69.14 24.535 69.615 24.735 ;
      RECT 69.14 24.135 69.42 24.735 ;
      RECT 68.455 17.065 68.98 17.285 ;
      RECT 68.81 16 68.98 17.285 ;
      RECT 68.81 16 69.34 16.365 ;
      RECT 68.445 27.865 68.91 28.195 ;
      RECT 68.59 26.905 68.91 28.195 ;
      RECT 68.54 24.535 68.87 24.735 ;
      RECT 68.585 24.135 68.87 24.735 ;
      RECT 68.115 17.485 68.45 17.655 ;
      RECT 68.115 17.215 68.285 17.655 ;
      RECT 68.06 15.98 68.23 17.345 ;
      RECT 68.115 15.555 68.365 16.11 ;
      RECT 68.18 22.875 68.435 23.205 ;
      RECT 68.265 20.995 68.435 23.205 ;
      RECT 68.225 22.865 68.435 23.205 ;
      RECT 68.25 22.795 68.435 23.205 ;
      RECT 68.18 20.995 68.435 21.665 ;
      RECT 67.995 24.565 68.37 24.735 ;
      RECT 68.005 24.535 68.37 24.735 ;
      RECT 67.89 28.365 68.295 28.535 ;
      RECT 67.89 26.435 68.06 28.535 ;
      RECT 67.23 27.835 68.06 28.135 ;
      RECT 67.23 27.805 67.43 28.135 ;
      RECT 67.89 26.435 68.14 26.765 ;
      RECT 65.93 22.955 67.465 23.205 ;
      RECT 67.295 22.555 67.465 23.205 ;
      RECT 65.035 22.555 65.205 23.205 ;
      RECT 65.93 22.555 66.1 23.205 ;
      RECT 67.295 22.555 68.095 22.725 ;
      RECT 67.925 21.835 68.095 22.725 ;
      RECT 65.035 22.555 66.1 22.725 ;
      RECT 65.035 21.835 68.095 22.005 ;
      RECT 65.035 20.995 65.205 22.005 ;
      RECT 67.72 19.815 67.975 20.485 ;
      RECT 67.805 18.275 67.975 20.485 ;
      RECT 67.79 18.275 67.975 18.685 ;
      RECT 67.72 18.275 67.975 18.605 ;
      RECT 66.345 28.365 67.02 28.535 ;
      RECT 66.85 27.415 67.02 28.535 ;
      RECT 67.55 27.325 67.72 27.655 ;
      RECT 66.85 27.415 67.72 27.585 ;
      RECT 67.21 27.325 67.72 27.585 ;
      RECT 67.21 26.54 67.38 27.585 ;
      RECT 66.275 26.54 67.38 26.71 ;
      RECT 67.33 22.185 67.695 22.385 ;
      RECT 67.33 22.185 67.705 22.355 ;
      RECT 64.575 19.475 64.745 20.485 ;
      RECT 64.575 19.475 67.635 19.645 ;
      RECT 67.465 18.755 67.635 19.645 ;
      RECT 66.835 18.755 67.635 18.925 ;
      RECT 64.575 18.755 65.64 18.925 ;
      RECT 65.47 18.275 65.64 18.925 ;
      RECT 66.835 18.275 67.005 18.925 ;
      RECT 64.575 18.275 64.745 18.925 ;
      RECT 65.47 18.275 67.005 18.525 ;
      RECT 67.265 25.255 67.52 25.925 ;
      RECT 67.265 23.715 67.435 25.925 ;
      RECT 67.265 23.715 67.45 24.125 ;
      RECT 67.265 23.715 67.52 24.045 ;
      RECT 65.875 21.425 67.51 21.665 ;
      RECT 67.26 20.995 67.51 21.665 ;
      RECT 65.875 21.335 66.105 21.665 ;
      RECT 66.83 22.185 67.115 22.785 ;
      RECT 66.83 22.185 67.16 22.385 ;
      RECT 66.415 17.215 66.585 17.675 ;
      RECT 66.415 17.215 67.08 17.385 ;
      RECT 66.85 16.055 67.08 17.385 ;
      RECT 66.415 16.055 67.08 16.225 ;
      RECT 66.415 15.555 66.585 16.225 ;
      RECT 66.8 14.375 67.055 15.045 ;
      RECT 66.885 12.835 67.055 15.045 ;
      RECT 66.87 12.835 67.055 13.245 ;
      RECT 66.8 12.835 67.055 13.165 ;
      RECT 66.8 19.815 67.05 20.485 ;
      RECT 65.415 19.815 65.645 20.145 ;
      RECT 65.415 19.815 67.05 20.055 ;
      RECT 66.155 27.945 66.68 28.165 ;
      RECT 66.51 26.88 66.68 28.165 ;
      RECT 66.51 26.88 67.04 27.245 ;
      RECT 63.655 14.035 63.825 15.045 ;
      RECT 63.655 14.035 66.715 14.205 ;
      RECT 66.545 13.315 66.715 14.205 ;
      RECT 65.915 13.315 66.715 13.485 ;
      RECT 63.655 13.315 64.72 13.485 ;
      RECT 64.55 12.835 64.72 13.485 ;
      RECT 65.915 12.835 66.085 13.485 ;
      RECT 63.655 12.835 63.825 13.485 ;
      RECT 64.55 12.835 66.085 13.085 ;
      RECT 66.37 19.095 66.7 19.295 ;
      RECT 66.37 18.695 66.655 19.295 ;
      RECT 66.28 22.185 66.56 22.785 ;
      RECT 66.085 22.185 66.56 22.385 ;
      RECT 65.375 20.995 65.705 21.665 ;
      RECT 66.215 20.995 66.545 21.205 ;
      RECT 65.375 20.995 66.545 21.165 ;
      RECT 65.95 13.685 66.325 13.855 ;
      RECT 65.95 13.655 66.315 13.855 ;
      RECT 65.815 28.365 66.15 28.535 ;
      RECT 65.815 28.095 65.985 28.535 ;
      RECT 65.76 26.86 65.93 28.225 ;
      RECT 65.815 26.435 66.065 26.99 ;
      RECT 65.895 17.115 66.065 17.765 ;
      RECT 65.055 17.115 65.225 17.76 ;
      RECT 64.645 17.115 66.065 17.285 ;
      RECT 64.645 16.405 64.82 17.285 ;
      RECT 62.195 16.775 64.82 16.945 ;
      RECT 64.645 16.405 66.145 16.575 ;
      RECT 65.815 15.555 66.145 16.575 ;
      RECT 64.975 15.555 65.305 16.575 ;
      RECT 65.88 14.375 66.13 15.045 ;
      RECT 64.495 14.375 64.725 14.705 ;
      RECT 64.495 14.375 66.13 14.615 ;
      RECT 65.625 19.095 66.1 19.295 ;
      RECT 65.82 18.695 66.1 19.295 ;
      RECT 64.915 20.315 66.085 20.485 ;
      RECT 65.755 20.275 66.085 20.485 ;
      RECT 64.915 19.815 65.245 20.485 ;
      RECT 65.45 13.655 65.78 13.855 ;
      RECT 65.45 13.255 65.735 13.855 ;
      RECT 65.01 19.095 65.18 19.305 ;
      RECT 65.01 19.095 65.455 19.295 ;
      RECT 64.705 13.655 65.18 13.855 ;
      RECT 64.9 13.255 65.18 13.855 ;
      RECT 63.995 14.875 65.165 15.045 ;
      RECT 64.835 14.835 65.165 15.045 ;
      RECT 63.995 14.375 64.325 15.045 ;
      RECT 64.115 28.095 64.285 28.555 ;
      RECT 64.115 28.095 64.78 28.265 ;
      RECT 64.55 26.935 64.78 28.265 ;
      RECT 64.115 26.935 64.78 27.105 ;
      RECT 64.115 26.435 64.285 27.105 ;
      RECT 60.435 11.675 60.605 12.325 ;
      RECT 61.275 11.675 61.445 12.32 ;
      RECT 60.435 11.675 61.855 11.845 ;
      RECT 61.68 10.965 61.855 11.845 ;
      RECT 61.68 11.335 64.305 11.505 ;
      RECT 60.355 10.965 61.855 11.135 ;
      RECT 61.195 10.115 61.525 11.135 ;
      RECT 60.355 10.115 60.685 11.135 ;
      RECT 62.12 19.48 62.38 20.455 ;
      RECT 61.265 19.48 61.52 20.455 ;
      RECT 60.405 19.48 60.66 20.455 ;
      RECT 59.905 19.48 62.935 19.65 ;
      RECT 62.635 18.745 62.935 19.65 ;
      RECT 59.905 18.745 60.075 19.65 ;
      RECT 59.485 19.125 60.075 19.295 ;
      RECT 59.905 18.745 62.935 18.915 ;
      RECT 61.69 18.3 61.945 18.915 ;
      RECT 60.83 18.3 61.09 18.915 ;
      RECT 59.945 11.305 60.115 12.155 ;
      RECT 60.4 11.305 61.5 11.505 ;
      RECT 59.945 11.305 61.5 11.475 ;
      RECT 58.415 17.195 58.745 17.715 ;
      RECT 58.625 16.445 58.795 17.28 ;
      RECT 58.57 17.155 58.795 17.28 ;
      RECT 58.58 16.445 58.795 16.575 ;
      RECT 58.405 15.6 58.735 16.525 ;
      RECT 58.415 28.075 58.745 28.595 ;
      RECT 58.625 27.325 58.795 28.16 ;
      RECT 58.57 28.035 58.795 28.16 ;
      RECT 58.58 27.325 58.795 27.455 ;
      RECT 58.405 26.48 58.735 27.405 ;
      RECT 57.575 17.195 57.905 17.72 ;
      RECT 57.705 16.695 57.905 17.72 ;
      RECT 57.705 16.695 58.455 17.025 ;
      RECT 57.705 15.555 57.895 17.72 ;
      RECT 57 16.115 57.895 16.49 ;
      RECT 57.555 15.555 57.895 16.49 ;
      RECT 57.575 28.075 57.905 28.6 ;
      RECT 57.705 27.575 57.905 28.6 ;
      RECT 57.705 27.575 58.455 27.905 ;
      RECT 57.705 26.435 57.895 28.6 ;
      RECT 57 26.995 57.895 27.37 ;
      RECT 57.555 26.435 57.895 27.37 ;
      RECT 56.045 17.485 56.83 17.655 ;
      RECT 56.66 15.685 56.83 17.655 ;
      RECT 56.66 16.695 57.535 17.025 ;
      RECT 55.945 15.685 56.83 15.855 ;
      RECT 56.045 28.365 56.83 28.535 ;
      RECT 56.66 26.565 56.83 28.535 ;
      RECT 56.66 27.575 57.535 27.905 ;
      RECT 55.945 26.565 56.83 26.735 ;
      RECT 56.025 16.985 56.49 17.315 ;
      RECT 56.17 16.025 56.49 17.315 ;
      RECT 56.025 27.865 56.49 28.195 ;
      RECT 56.17 26.905 56.49 28.195 ;
      RECT 55.775 14.035 55.945 15.045 ;
      RECT 52.885 14.035 55.945 14.205 ;
      RECT 52.885 13.315 53.055 14.205 ;
      RECT 54.88 13.315 55.945 13.485 ;
      RECT 55.775 12.835 55.945 13.485 ;
      RECT 52.885 13.315 53.685 13.485 ;
      RECT 53.515 12.835 53.685 13.485 ;
      RECT 54.88 12.835 55.05 13.485 ;
      RECT 53.515 12.835 55.05 13.085 ;
      RECT 55.47 17.485 55.875 17.655 ;
      RECT 55.47 15.555 55.64 17.655 ;
      RECT 54.81 16.955 55.64 17.255 ;
      RECT 54.81 16.925 55.01 17.255 ;
      RECT 55.47 15.555 55.72 15.885 ;
      RECT 55.47 28.365 55.875 28.535 ;
      RECT 55.47 26.435 55.64 28.535 ;
      RECT 54.81 27.835 55.64 28.135 ;
      RECT 54.81 27.805 55.01 28.135 ;
      RECT 55.47 26.435 55.72 26.765 ;
      RECT 54.435 14.875 55.605 15.045 ;
      RECT 55.275 14.375 55.605 15.045 ;
      RECT 54.435 14.835 54.765 15.045 ;
      RECT 53.925 17.485 54.6 17.655 ;
      RECT 54.43 16.535 54.6 17.655 ;
      RECT 55.13 16.445 55.3 16.775 ;
      RECT 54.43 16.535 55.3 16.705 ;
      RECT 54.79 16.445 55.3 16.705 ;
      RECT 54.79 15.66 54.96 16.705 ;
      RECT 53.855 15.66 54.96 15.83 ;
      RECT 53.925 28.365 54.6 28.535 ;
      RECT 54.43 27.415 54.6 28.535 ;
      RECT 55.13 27.325 55.3 27.655 ;
      RECT 54.43 27.415 55.3 27.585 ;
      RECT 54.79 27.325 55.3 27.585 ;
      RECT 54.79 26.54 54.96 27.585 ;
      RECT 53.855 26.54 54.96 26.71 ;
      RECT 53.47 14.375 53.72 15.045 ;
      RECT 54.875 14.375 55.105 14.705 ;
      RECT 53.47 14.375 55.105 14.615 ;
      RECT 54.42 13.655 54.895 13.855 ;
      RECT 54.42 13.255 54.7 13.855 ;
      RECT 53.735 17.065 54.26 17.285 ;
      RECT 54.09 16 54.26 17.285 ;
      RECT 54.09 16 54.62 16.365 ;
      RECT 53.735 27.945 54.26 28.165 ;
      RECT 54.09 26.88 54.26 28.165 ;
      RECT 54.09 26.88 54.62 27.245 ;
      RECT 53.805 19.515 54.135 20.44 ;
      RECT 54.025 18.76 54.195 19.595 ;
      RECT 53.98 19.465 54.195 19.595 ;
      RECT 53.97 18.76 54.195 18.885 ;
      RECT 53.815 18.325 54.145 18.845 ;
      RECT 53.82 13.655 54.15 13.855 ;
      RECT 53.865 13.255 54.15 13.855 ;
      RECT 52.955 19.55 53.295 20.485 ;
      RECT 53.105 18.32 53.295 20.485 ;
      RECT 52.4 19.55 53.295 19.925 ;
      RECT 53.105 19.015 53.855 19.345 ;
      RECT 53.105 18.32 53.305 19.345 ;
      RECT 52.975 18.32 53.305 18.845 ;
      RECT 53.395 17.485 53.73 17.655 ;
      RECT 53.395 17.215 53.565 17.655 ;
      RECT 53.34 15.98 53.51 17.345 ;
      RECT 53.395 15.555 53.645 16.11 ;
      RECT 53.395 28.365 53.73 28.535 ;
      RECT 53.395 28.095 53.565 28.535 ;
      RECT 53.34 26.86 53.51 28.225 ;
      RECT 53.395 26.435 53.645 26.99 ;
      RECT 53.275 13.685 53.65 13.855 ;
      RECT 53.285 13.655 53.65 13.855 ;
      RECT 51.345 20.185 52.23 20.355 ;
      RECT 52.06 18.385 52.23 20.355 ;
      RECT 52.06 19.015 52.935 19.345 ;
      RECT 51.445 18.385 52.23 18.555 ;
      RECT 52.545 14.375 52.8 15.045 ;
      RECT 52.545 12.835 52.715 15.045 ;
      RECT 52.545 12.835 52.73 13.245 ;
      RECT 52.545 12.835 52.8 13.165 ;
      RECT 51.695 17.215 51.865 17.675 ;
      RECT 51.695 17.215 52.36 17.385 ;
      RECT 52.13 16.055 52.36 17.385 ;
      RECT 51.695 16.055 52.36 16.225 ;
      RECT 51.695 15.555 51.865 16.225 ;
      RECT 51.695 28.095 51.865 28.555 ;
      RECT 51.695 28.095 52.36 28.265 ;
      RECT 52.13 26.935 52.36 28.265 ;
      RECT 51.695 26.935 52.36 27.105 ;
      RECT 51.695 26.435 51.865 27.105 ;
      RECT 51.57 18.725 51.89 20.015 ;
      RECT 51.425 18.725 51.89 19.055 ;
      RECT 50.87 20.155 51.12 20.485 ;
      RECT 50.87 18.385 51.04 20.485 ;
      RECT 50.21 18.785 50.41 19.115 ;
      RECT 50.21 18.785 51.04 19.085 ;
      RECT 50.87 18.385 51.275 18.555 ;
      RECT 47.095 11.675 47.265 12.325 ;
      RECT 47.935 11.675 48.105 12.32 ;
      RECT 47.095 11.675 48.515 11.845 ;
      RECT 48.34 10.965 48.515 11.845 ;
      RECT 48.34 11.335 50.965 11.505 ;
      RECT 47.015 10.965 48.515 11.135 ;
      RECT 47.855 10.115 48.185 11.135 ;
      RECT 47.015 10.115 47.345 11.135 ;
      RECT 49.255 20.21 50.36 20.38 ;
      RECT 50.19 19.335 50.36 20.38 ;
      RECT 50.19 19.335 50.7 19.595 ;
      RECT 50.53 19.265 50.7 19.595 ;
      RECT 49.83 19.335 50.7 19.505 ;
      RECT 49.83 18.385 50 19.505 ;
      RECT 49.325 18.385 50 18.555 ;
      RECT 50.175 24.905 50.505 25.925 ;
      RECT 49.335 24.905 49.665 25.925 ;
      RECT 49.005 24.905 50.505 25.075 ;
      RECT 49.005 24.195 49.18 25.075 ;
      RECT 46.555 24.535 49.18 24.705 ;
      RECT 49.005 24.195 50.425 24.365 ;
      RECT 50.255 23.715 50.425 24.365 ;
      RECT 49.415 23.72 49.585 24.365 ;
      RECT 49.49 19.675 50.02 20.04 ;
      RECT 49.49 18.755 49.66 20.04 ;
      RECT 49.135 18.755 49.66 18.975 ;
      RECT 49.32 14.375 49.575 15.045 ;
      RECT 49.405 12.835 49.575 15.045 ;
      RECT 49.39 12.835 49.575 13.245 ;
      RECT 49.32 12.835 49.575 13.165 ;
      RECT 46.175 14.035 46.345 15.045 ;
      RECT 46.175 14.035 49.235 14.205 ;
      RECT 49.065 13.315 49.235 14.205 ;
      RECT 48.435 13.315 49.235 13.485 ;
      RECT 46.175 13.315 47.24 13.485 ;
      RECT 47.07 12.835 47.24 13.485 ;
      RECT 48.435 12.835 48.605 13.485 ;
      RECT 46.175 12.835 46.345 13.485 ;
      RECT 47.07 12.835 48.605 13.085 ;
      RECT 48.795 19.93 49.045 20.485 ;
      RECT 48.74 18.695 48.91 20.06 ;
      RECT 48.795 18.385 48.965 18.825 ;
      RECT 48.795 18.385 49.13 18.555 ;
      RECT 48.47 13.685 48.845 13.855 ;
      RECT 48.47 13.655 48.835 13.855 ;
      RECT 48.4 14.375 48.65 15.045 ;
      RECT 47.015 14.375 47.245 14.705 ;
      RECT 47.015 14.375 48.65 14.615 ;
      RECT 47.97 13.655 48.3 13.855 ;
      RECT 47.97 13.255 48.255 13.855 ;
      RECT 47.095 19.815 47.265 20.485 ;
      RECT 47.095 19.815 47.76 19.985 ;
      RECT 47.53 18.655 47.76 19.985 ;
      RECT 47.095 18.655 47.76 18.825 ;
      RECT 47.095 18.365 47.265 18.825 ;
      RECT 47.225 13.655 47.7 13.855 ;
      RECT 47.42 13.255 47.7 13.855 ;
      RECT 46.515 14.875 47.685 15.045 ;
      RECT 47.355 14.835 47.685 15.045 ;
      RECT 46.515 14.375 46.845 15.045 ;
      RECT 43.695 28.075 44.025 28.595 ;
      RECT 43.905 27.325 44.075 28.16 ;
      RECT 43.85 28.035 44.075 28.16 ;
      RECT 43.86 27.325 44.075 27.455 ;
      RECT 43.685 26.48 44.015 27.405 ;
      RECT 43.845 22.185 44.015 23.035 ;
      RECT 42.46 22.185 43.56 22.385 ;
      RECT 42.46 22.185 44.015 22.355 ;
      RECT 42.855 28.075 43.185 28.6 ;
      RECT 42.985 27.575 43.185 28.6 ;
      RECT 42.985 27.575 43.735 27.905 ;
      RECT 42.985 26.435 43.175 28.6 ;
      RECT 42.28 26.995 43.175 27.37 ;
      RECT 42.835 26.435 43.175 27.37 ;
      RECT 43.355 22.555 43.525 23.205 ;
      RECT 42.515 22.555 42.685 23.2 ;
      RECT 42.105 22.555 43.525 22.725 ;
      RECT 42.105 21.845 42.28 22.725 ;
      RECT 39.655 22.215 42.28 22.385 ;
      RECT 42.105 21.845 43.605 22.015 ;
      RECT 43.275 20.995 43.605 22.015 ;
      RECT 42.435 20.995 42.765 22.015 ;
      RECT 41.325 28.365 42.11 28.535 ;
      RECT 41.94 26.565 42.11 28.535 ;
      RECT 41.94 27.575 42.815 27.905 ;
      RECT 41.225 26.565 42.11 26.735 ;
      RECT 41.305 27.865 41.77 28.195 ;
      RECT 41.45 26.905 41.77 28.195 ;
      RECT 40.75 28.365 41.155 28.535 ;
      RECT 40.75 26.435 40.92 28.535 ;
      RECT 40.09 27.835 40.92 28.135 ;
      RECT 40.09 27.805 40.29 28.135 ;
      RECT 40.75 26.435 41 26.765 ;
      RECT 40.465 19.515 40.795 20.44 ;
      RECT 40.685 18.76 40.855 19.595 ;
      RECT 40.64 19.465 40.855 19.595 ;
      RECT 40.63 18.76 40.855 18.885 ;
      RECT 40.475 18.325 40.805 18.845 ;
      RECT 36.975 11.675 37.145 12.325 ;
      RECT 37.815 11.675 37.985 12.32 ;
      RECT 36.975 11.675 38.395 11.845 ;
      RECT 38.22 10.965 38.395 11.845 ;
      RECT 38.22 11.335 40.845 11.505 ;
      RECT 36.895 10.965 38.395 11.135 ;
      RECT 37.735 10.115 38.065 11.135 ;
      RECT 36.895 10.115 37.225 11.135 ;
      RECT 39.205 28.365 39.88 28.535 ;
      RECT 39.71 27.415 39.88 28.535 ;
      RECT 40.41 27.325 40.58 27.655 ;
      RECT 39.71 27.415 40.58 27.585 ;
      RECT 40.07 27.325 40.58 27.585 ;
      RECT 40.07 26.54 40.24 27.585 ;
      RECT 39.135 26.54 40.24 26.71 ;
      RECT 39.615 19.55 39.955 20.485 ;
      RECT 39.765 18.32 39.955 20.485 ;
      RECT 39.06 19.55 39.955 19.925 ;
      RECT 39.765 19.015 40.515 19.345 ;
      RECT 39.765 18.32 39.965 19.345 ;
      RECT 39.635 18.32 39.965 18.845 ;
      RECT 40.015 17.195 40.345 17.715 ;
      RECT 40.225 16.445 40.395 17.28 ;
      RECT 40.17 17.155 40.395 17.28 ;
      RECT 40.18 16.445 40.395 16.575 ;
      RECT 40.005 15.6 40.335 16.525 ;
      RECT 40.005 35.835 40.335 36.76 ;
      RECT 40.225 35.08 40.395 35.915 ;
      RECT 40.18 35.785 40.395 35.915 ;
      RECT 40.17 35.08 40.395 35.205 ;
      RECT 40.015 34.645 40.345 35.165 ;
      RECT 39.175 17.195 39.505 17.72 ;
      RECT 39.305 16.695 39.505 17.72 ;
      RECT 39.305 16.695 40.055 17.025 ;
      RECT 39.305 15.555 39.495 17.72 ;
      RECT 38.6 16.115 39.495 16.49 ;
      RECT 39.155 15.555 39.495 16.49 ;
      RECT 39.155 35.87 39.495 36.805 ;
      RECT 39.305 34.64 39.495 36.805 ;
      RECT 38.6 35.87 39.495 36.245 ;
      RECT 39.305 35.335 40.055 35.665 ;
      RECT 39.305 34.64 39.505 35.665 ;
      RECT 39.175 34.64 39.505 35.165 ;
      RECT 39.015 27.945 39.54 28.165 ;
      RECT 39.37 26.88 39.54 28.165 ;
      RECT 39.37 26.88 39.9 27.245 ;
      RECT 38.005 20.185 38.89 20.355 ;
      RECT 38.72 18.385 38.89 20.355 ;
      RECT 38.72 19.015 39.595 19.345 ;
      RECT 38.105 18.385 38.89 18.555 ;
      RECT 37.645 17.485 38.43 17.655 ;
      RECT 38.26 15.685 38.43 17.655 ;
      RECT 38.26 16.695 39.135 17.025 ;
      RECT 37.545 15.685 38.43 15.855 ;
      RECT 37.545 36.505 38.43 36.675 ;
      RECT 38.26 34.705 38.43 36.675 ;
      RECT 38.26 35.335 39.135 35.665 ;
      RECT 37.645 34.705 38.43 34.875 ;
      RECT 38.675 28.365 39.01 28.535 ;
      RECT 38.675 28.095 38.845 28.535 ;
      RECT 38.62 26.86 38.79 28.225 ;
      RECT 38.675 26.435 38.925 26.99 ;
      RECT 38.23 18.725 38.55 20.015 ;
      RECT 38.085 18.725 38.55 19.055 ;
      RECT 38.28 14.375 38.535 15.045 ;
      RECT 38.365 12.835 38.535 15.045 ;
      RECT 38.35 12.835 38.535 13.245 ;
      RECT 38.28 12.835 38.535 13.165 ;
      RECT 38.28 25.255 38.535 25.925 ;
      RECT 38.365 23.715 38.535 25.925 ;
      RECT 38.35 23.715 38.535 24.125 ;
      RECT 38.28 23.715 38.535 24.045 ;
      RECT 38.28 30.695 38.535 31.365 ;
      RECT 38.365 29.155 38.535 31.365 ;
      RECT 38.35 29.155 38.535 29.565 ;
      RECT 38.325 29.155 38.535 29.495 ;
      RECT 38.28 29.155 38.535 29.485 ;
      RECT 38.28 33.755 38.535 34.085 ;
      RECT 38.365 31.875 38.535 34.085 ;
      RECT 38.325 33.745 38.535 34.085 ;
      RECT 38.35 33.675 38.535 34.085 ;
      RECT 38.28 31.875 38.535 32.545 ;
      RECT 35.135 14.035 35.305 15.045 ;
      RECT 35.135 14.035 38.195 14.205 ;
      RECT 38.025 13.315 38.195 14.205 ;
      RECT 37.395 13.315 38.195 13.485 ;
      RECT 35.135 13.315 36.2 13.485 ;
      RECT 36.03 12.835 36.2 13.485 ;
      RECT 37.395 12.835 37.565 13.485 ;
      RECT 35.135 12.835 35.305 13.485 ;
      RECT 36.03 12.835 37.565 13.085 ;
      RECT 35.135 24.915 35.305 25.925 ;
      RECT 35.135 24.915 38.195 25.085 ;
      RECT 38.025 24.195 38.195 25.085 ;
      RECT 37.395 24.195 38.195 24.365 ;
      RECT 35.135 24.195 36.2 24.365 ;
      RECT 36.03 23.715 36.2 24.365 ;
      RECT 37.395 23.715 37.565 24.365 ;
      RECT 35.135 23.715 35.305 24.365 ;
      RECT 36.03 23.715 37.565 23.965 ;
      RECT 35.135 30.355 35.305 31.365 ;
      RECT 35.135 30.355 38.195 30.525 ;
      RECT 38.025 29.635 38.195 30.525 ;
      RECT 37.395 29.635 38.195 29.805 ;
      RECT 35.135 29.635 36.2 29.805 ;
      RECT 36.03 29.155 36.2 29.805 ;
      RECT 37.395 29.155 37.565 29.805 ;
      RECT 35.135 29.155 35.305 29.805 ;
      RECT 36.03 29.155 37.565 29.405 ;
      RECT 36.03 33.835 37.565 34.085 ;
      RECT 37.395 33.435 37.565 34.085 ;
      RECT 35.135 33.435 35.305 34.085 ;
      RECT 36.03 33.435 36.2 34.085 ;
      RECT 37.395 33.435 38.195 33.605 ;
      RECT 38.025 32.715 38.195 33.605 ;
      RECT 35.135 33.435 36.2 33.605 ;
      RECT 35.135 32.715 38.195 32.885 ;
      RECT 35.135 31.875 35.305 32.885 ;
      RECT 37.625 16.985 38.09 17.315 ;
      RECT 37.77 16.025 38.09 17.315 ;
      RECT 37.77 35.045 38.09 36.335 ;
      RECT 37.625 35.045 38.09 35.375 ;
      RECT 36.94 11.305 38.04 11.505 ;
      RECT 36.485 11.305 38.04 11.475 ;
      RECT 36.485 10.965 36.655 11.475 ;
      RECT 37.53 20.155 37.78 20.485 ;
      RECT 37.53 18.385 37.7 20.485 ;
      RECT 36.87 18.785 37.07 19.115 ;
      RECT 36.87 18.785 37.7 19.085 ;
      RECT 37.53 18.385 37.935 18.555 ;
      RECT 37.43 13.685 37.805 13.855 ;
      RECT 37.43 13.655 37.795 13.855 ;
      RECT 37.43 24.565 37.805 24.735 ;
      RECT 37.43 24.535 37.795 24.735 ;
      RECT 37.43 30.005 37.805 30.175 ;
      RECT 37.43 29.975 37.795 30.175 ;
      RECT 37.43 33.065 37.795 33.265 ;
      RECT 37.43 33.065 37.805 33.235 ;
      RECT 36.975 28.095 37.145 28.555 ;
      RECT 36.975 28.095 37.64 28.265 ;
      RECT 37.41 26.935 37.64 28.265 ;
      RECT 36.975 26.935 37.64 27.105 ;
      RECT 36.975 26.435 37.145 27.105 ;
      RECT 37.36 14.375 37.61 15.045 ;
      RECT 35.975 14.375 36.205 14.705 ;
      RECT 35.975 14.375 37.61 14.615 ;
      RECT 37.36 25.255 37.61 25.925 ;
      RECT 35.975 25.255 36.205 25.585 ;
      RECT 35.975 25.255 37.61 25.495 ;
      RECT 37.36 30.695 37.61 31.365 ;
      RECT 35.975 30.695 36.205 31.025 ;
      RECT 35.975 30.695 37.61 30.935 ;
      RECT 35.975 32.305 37.61 32.545 ;
      RECT 37.36 31.875 37.61 32.545 ;
      RECT 35.975 32.215 36.205 32.545 ;
      RECT 37.07 17.485 37.475 17.655 ;
      RECT 37.07 15.555 37.24 17.655 ;
      RECT 36.41 16.955 37.24 17.255 ;
      RECT 36.41 16.925 36.61 17.255 ;
      RECT 37.07 15.555 37.32 15.885 ;
      RECT 37.07 36.475 37.32 36.805 ;
      RECT 37.07 34.705 37.24 36.805 ;
      RECT 36.41 35.105 36.61 35.435 ;
      RECT 36.41 35.105 37.24 35.405 ;
      RECT 37.07 34.705 37.475 34.875 ;
      RECT 35.915 20.21 37.02 20.38 ;
      RECT 36.85 19.335 37.02 20.38 ;
      RECT 36.85 19.335 37.36 19.595 ;
      RECT 37.19 19.265 37.36 19.595 ;
      RECT 36.49 19.335 37.36 19.505 ;
      RECT 36.49 18.385 36.66 19.505 ;
      RECT 35.985 18.385 36.66 18.555 ;
      RECT 36.93 13.655 37.26 13.855 ;
      RECT 36.93 13.255 37.215 13.855 ;
      RECT 36.93 24.535 37.26 24.735 ;
      RECT 36.93 24.135 37.215 24.735 ;
      RECT 36.93 29.975 37.26 30.175 ;
      RECT 36.93 29.575 37.215 30.175 ;
      RECT 36.93 33.065 37.215 33.665 ;
      RECT 36.93 33.065 37.26 33.265 ;
      RECT 35.525 17.485 36.2 17.655 ;
      RECT 36.03 16.535 36.2 17.655 ;
      RECT 36.73 16.445 36.9 16.775 ;
      RECT 36.03 16.535 36.9 16.705 ;
      RECT 36.39 16.445 36.9 16.705 ;
      RECT 36.39 15.66 36.56 16.705 ;
      RECT 35.455 15.66 36.56 15.83 ;
      RECT 35.455 36.53 36.56 36.7 ;
      RECT 36.39 35.655 36.56 36.7 ;
      RECT 36.39 35.655 36.9 35.915 ;
      RECT 36.73 35.585 36.9 35.915 ;
      RECT 36.03 35.655 36.9 35.825 ;
      RECT 36.03 34.705 36.2 35.825 ;
      RECT 35.525 34.705 36.2 34.875 ;
      RECT 36.15 19.675 36.68 20.04 ;
      RECT 36.15 18.755 36.32 20.04 ;
      RECT 35.795 18.755 36.32 18.975 ;
      RECT 36.185 13.655 36.66 13.855 ;
      RECT 36.38 13.255 36.66 13.855 ;
      RECT 36.185 24.535 36.66 24.735 ;
      RECT 36.38 24.135 36.66 24.735 ;
      RECT 36.185 29.975 36.66 30.175 ;
      RECT 36.38 29.575 36.66 30.175 ;
      RECT 36.38 33.065 36.66 33.665 ;
      RECT 36.185 33.065 36.66 33.265 ;
      RECT 35.475 14.875 36.645 15.045 ;
      RECT 36.315 14.835 36.645 15.045 ;
      RECT 35.475 14.375 35.805 15.045 ;
      RECT 35.475 25.755 36.645 25.925 ;
      RECT 36.315 25.715 36.645 25.925 ;
      RECT 35.475 25.255 35.805 25.925 ;
      RECT 35.475 31.195 36.645 31.365 ;
      RECT 36.315 31.155 36.645 31.365 ;
      RECT 35.475 30.695 35.805 31.365 ;
      RECT 35.475 31.875 35.805 32.545 ;
      RECT 36.315 31.875 36.645 32.085 ;
      RECT 35.475 31.875 36.645 32.045 ;
      RECT 35.335 17.065 35.86 17.285 ;
      RECT 35.69 16 35.86 17.285 ;
      RECT 35.69 16 36.22 16.365 ;
      RECT 35.69 35.995 36.22 36.36 ;
      RECT 35.69 35.075 35.86 36.36 ;
      RECT 35.335 35.075 35.86 35.295 ;
      RECT 36.025 10.285 36.195 11.815 ;
      RECT 34.605 10.285 36.195 10.455 ;
      RECT 34.605 10.165 35.795 10.455 ;
      RECT 35.455 19.93 35.705 20.485 ;
      RECT 35.4 18.695 35.57 20.06 ;
      RECT 35.455 18.385 35.625 18.825 ;
      RECT 35.455 18.385 35.79 18.555 ;
      RECT 35.525 11.755 35.78 12.275 ;
      RECT 34.685 11.755 34.855 12.275 ;
      RECT 34.115 11.755 35.78 11.925 ;
      RECT 34.115 10.915 34.285 11.925 ;
      RECT 34.01 11.255 34.285 11.585 ;
      RECT 35.45 10.625 35.775 11.085 ;
      RECT 34.115 10.915 34.775 11.085 ;
      RECT 34.605 10.625 34.775 11.085 ;
      RECT 34.605 10.625 35.775 10.795 ;
      RECT 34.995 17.485 35.33 17.655 ;
      RECT 34.995 17.215 35.165 17.655 ;
      RECT 34.94 15.98 35.11 17.345 ;
      RECT 34.995 15.555 35.245 16.11 ;
      RECT 34.995 36.25 35.245 36.805 ;
      RECT 34.94 35.015 35.11 36.38 ;
      RECT 34.995 34.705 35.165 35.145 ;
      RECT 34.995 34.705 35.33 34.875 ;
      RECT 35.075 22.555 35.245 23.205 ;
      RECT 34.235 22.555 34.405 23.2 ;
      RECT 33.825 22.555 35.245 22.725 ;
      RECT 33.825 21.845 34 22.725 ;
      RECT 31.375 22.215 34 22.385 ;
      RECT 33.825 21.845 35.325 22.015 ;
      RECT 34.995 20.995 35.325 22.015 ;
      RECT 34.155 20.995 34.485 22.015 ;
      RECT 34.455 11.255 35.28 11.585 ;
      RECT 35.085 10.965 35.28 11.585 ;
      RECT 33.755 19.815 33.925 20.485 ;
      RECT 33.755 19.815 34.42 19.985 ;
      RECT 34.19 18.655 34.42 19.985 ;
      RECT 33.755 18.655 34.42 18.825 ;
      RECT 33.755 18.365 33.925 18.825 ;
      RECT 33.295 17.215 33.465 17.675 ;
      RECT 33.295 17.215 33.96 17.385 ;
      RECT 33.73 16.055 33.96 17.385 ;
      RECT 33.295 16.055 33.96 16.225 ;
      RECT 33.295 15.555 33.465 16.225 ;
      RECT 33.295 36.135 33.465 36.805 ;
      RECT 33.295 36.135 33.96 36.305 ;
      RECT 33.73 34.975 33.96 36.305 ;
      RECT 33.295 34.975 33.96 35.145 ;
      RECT 33.295 34.685 33.465 35.145 ;
      RECT 33.67 11.82 33.945 12.165 ;
      RECT 33.67 10.115 33.84 12.165 ;
      RECT 33.67 10.115 33.945 11.085 ;
      RECT 28.975 28.075 29.305 28.595 ;
      RECT 29.185 27.325 29.355 28.16 ;
      RECT 29.13 28.035 29.355 28.16 ;
      RECT 29.14 27.325 29.355 27.455 ;
      RECT 28.965 26.48 29.295 27.405 ;
      RECT 28.135 28.075 28.465 28.6 ;
      RECT 28.265 27.575 28.465 28.6 ;
      RECT 28.265 27.575 29.015 27.905 ;
      RECT 28.265 26.435 28.455 28.6 ;
      RECT 27.56 26.995 28.455 27.37 ;
      RECT 28.115 26.435 28.455 27.37 ;
      RECT 26.605 28.365 27.39 28.535 ;
      RECT 27.22 26.565 27.39 28.535 ;
      RECT 27.22 27.575 28.095 27.905 ;
      RECT 26.505 26.565 27.39 26.735 ;
      RECT 24.095 11.675 24.265 12.325 ;
      RECT 24.935 11.675 25.105 12.32 ;
      RECT 24.095 11.675 25.515 11.845 ;
      RECT 25.34 10.965 25.515 11.845 ;
      RECT 25.34 11.335 27.965 11.505 ;
      RECT 24.015 10.965 25.515 11.135 ;
      RECT 24.855 10.115 25.185 11.135 ;
      RECT 24.015 10.115 24.345 11.135 ;
      RECT 26.585 27.865 27.05 28.195 ;
      RECT 26.73 26.905 27.05 28.195 ;
      RECT 26.03 28.365 26.435 28.535 ;
      RECT 26.03 26.435 26.2 28.535 ;
      RECT 25.37 27.835 26.2 28.135 ;
      RECT 25.37 27.805 25.57 28.135 ;
      RECT 26.03 26.435 26.28 26.765 ;
      RECT 24.485 28.365 25.16 28.535 ;
      RECT 24.99 27.415 25.16 28.535 ;
      RECT 25.69 27.325 25.86 27.655 ;
      RECT 24.99 27.415 25.86 27.585 ;
      RECT 25.35 27.325 25.86 27.585 ;
      RECT 25.35 26.54 25.52 27.585 ;
      RECT 24.415 26.54 25.52 26.71 ;
      RECT 24.295 27.945 24.82 28.165 ;
      RECT 24.65 26.88 24.82 28.165 ;
      RECT 24.65 26.88 25.18 27.245 ;
      RECT 23.955 28.365 24.29 28.535 ;
      RECT 23.955 28.095 24.125 28.535 ;
      RECT 23.9 26.86 24.07 28.225 ;
      RECT 23.955 26.435 24.205 26.99 ;
      RECT 21.175 19.465 21.505 20.485 ;
      RECT 20.335 19.465 20.665 20.485 ;
      RECT 20.335 19.465 21.835 19.635 ;
      RECT 21.66 18.755 21.835 19.635 ;
      RECT 21.66 19.095 24.285 19.265 ;
      RECT 20.415 18.755 21.835 18.925 ;
      RECT 21.255 18.28 21.425 18.925 ;
      RECT 20.415 18.275 20.585 18.925 ;
      RECT 22.255 28.095 22.425 28.555 ;
      RECT 22.255 28.095 22.92 28.265 ;
      RECT 22.69 26.935 22.92 28.265 ;
      RECT 22.255 26.935 22.92 27.105 ;
      RECT 22.255 26.435 22.425 27.105 ;
      RECT 17.655 22.555 17.825 23.205 ;
      RECT 18.495 22.555 18.665 23.2 ;
      RECT 17.655 22.555 19.075 22.725 ;
      RECT 18.9 21.845 19.075 22.725 ;
      RECT 18.9 22.215 21.525 22.385 ;
      RECT 17.575 21.845 19.075 22.015 ;
      RECT 18.415 20.995 18.745 22.015 ;
      RECT 17.575 20.995 17.905 22.015 ;
      RECT 15.815 11.675 15.985 12.325 ;
      RECT 16.655 11.675 16.825 12.32 ;
      RECT 15.815 11.675 17.235 11.845 ;
      RECT 17.06 10.965 17.235 11.845 ;
      RECT 17.06 11.335 19.685 11.505 ;
      RECT 15.735 10.965 17.235 11.135 ;
      RECT 16.575 10.115 16.905 11.135 ;
      RECT 15.735 10.115 16.065 11.135 ;
      RECT 181.39 16.055 181.58 16.775 ;
      RECT 179.26 16.3 179.5 16.895 ;
      RECT 178.47 16.355 178.75 17.305 ;
      RECT 177.24 11.305 178.34 11.505 ;
      RECT 178.115 15.555 178.3 17.675 ;
      RECT 177.19 16.395 177.54 17.045 ;
      RECT 171.26 22.185 172.36 22.385 ;
      RECT 171.26 29.975 172.36 30.175 ;
      RECT 171.665 19.075 172.205 19.635 ;
      RECT 171.225 18.285 171.485 20.475 ;
      RECT 170.285 16.405 170.825 16.965 ;
      RECT 170.1 19.035 170.565 19.345 ;
      RECT 168.915 19.015 169.215 19.345 ;
      RECT 168.04 11.305 169.14 11.505 ;
      RECT 166.67 16.055 166.86 16.775 ;
      RECT 164.54 16.3 164.78 16.895 ;
      RECT 163.75 16.355 164.03 17.305 ;
      RECT 163.395 15.555 163.58 17.675 ;
      RECT 162.47 16.395 162.82 17.045 ;
      RECT 155.63 35.585 155.82 36.305 ;
      RECT 155.17 30.145 155.36 30.865 ;
      RECT 154.24 22.185 155.34 22.385 ;
      RECT 153.32 11.305 154.42 11.505 ;
      RECT 153.33 19.095 153.775 19.295 ;
      RECT 153.33 27.625 153.775 27.825 ;
      RECT 153.33 33.065 153.775 33.265 ;
      RECT 153.5 35.465 153.74 36.06 ;
      RECT 153.04 30.025 153.28 30.62 ;
      RECT 152.81 19.095 153.16 19.305 ;
      RECT 152.81 27.615 153.16 27.825 ;
      RECT 152.81 33.055 153.16 33.265 ;
      RECT 152.71 35.055 152.99 36.005 ;
      RECT 152.355 34.685 152.54 36.805 ;
      RECT 152.25 29.615 152.53 30.565 ;
      RECT 151.95 16.055 152.14 16.775 ;
      RECT 151.895 29.245 152.08 31.365 ;
      RECT 151.43 35.315 151.78 35.965 ;
      RECT 150.97 29.875 151.32 30.525 ;
      RECT 149.82 16.3 150.06 16.895 ;
      RECT 149.03 16.355 149.31 17.305 ;
      RECT 148.675 15.555 148.86 17.675 ;
      RECT 148.27 19.095 148.715 19.295 ;
      RECT 147.75 16.395 148.1 17.045 ;
      RECT 147.75 19.095 148.1 19.305 ;
      RECT 144 24.535 144.35 24.745 ;
      RECT 143.385 24.535 143.83 24.735 ;
      RECT 142.75 26.935 142.94 27.655 ;
      RECT 140.62 27.18 140.86 27.775 ;
      RECT 139.83 27.235 140.11 28.185 ;
      RECT 138.6 13.655 139.7 13.855 ;
      RECT 139.475 26.435 139.66 28.555 ;
      RECT 138.55 27.275 138.9 27.925 ;
      RECT 138.02 22.175 138.37 22.385 ;
      RECT 137.56 24.535 137.91 24.745 ;
      RECT 137.405 22.185 137.85 22.385 ;
      RECT 137.23 16.055 137.42 16.775 ;
      RECT 137.23 19.265 137.42 19.985 ;
      RECT 136.945 24.535 137.39 24.735 ;
      RECT 135.1 16.3 135.34 16.895 ;
      RECT 135.1 19.145 135.34 19.74 ;
      RECT 134.31 16.355 134.59 17.305 ;
      RECT 134.31 18.735 134.59 19.685 ;
      RECT 133.08 11.305 134.18 11.505 ;
      RECT 133.955 15.555 134.14 17.675 ;
      RECT 133.955 18.365 134.14 20.485 ;
      RECT 133.03 16.395 133.38 17.045 ;
      RECT 133.03 18.995 133.38 19.645 ;
      RECT 132.165 21.165 132.335 23.035 ;
      RECT 130.2 27.615 130.55 27.825 ;
      RECT 129.585 27.625 130.03 27.825 ;
      RECT 128.95 22.185 129.395 22.385 ;
      RECT 128.43 22.175 128.78 22.385 ;
      RECT 128.49 35.585 128.68 36.305 ;
      RECT 124.645 19.085 126.86 19.31 ;
      RECT 126.36 35.465 126.6 36.06 ;
      RECT 125.57 35.055 125.85 36.005 ;
      RECT 125.27 21.495 125.46 22.215 ;
      RECT 124.34 11.305 125.44 11.505 ;
      RECT 125.215 34.685 125.4 36.805 ;
      RECT 124.29 35.315 124.64 35.965 ;
      RECT 123.14 21.74 123.38 22.335 ;
      RECT 122.51 16.055 122.7 16.775 ;
      RECT 122.35 21.795 122.63 22.745 ;
      RECT 121.995 20.995 122.18 23.115 ;
      RECT 121.07 21.835 121.42 22.485 ;
      RECT 118.665 19.085 120.88 19.31 ;
      RECT 120.38 16.3 120.62 16.895 ;
      RECT 119.59 16.355 119.87 17.305 ;
      RECT 118.36 11.305 119.46 11.505 ;
      RECT 119.235 15.555 119.42 17.675 ;
      RECT 118.31 16.395 118.66 17.045 ;
      RECT 114.22 11.305 115.32 11.505 ;
      RECT 114.69 13.655 115.135 13.855 ;
      RECT 114.69 22.185 115.135 22.385 ;
      RECT 114.69 26.935 114.88 27.655 ;
      RECT 114.17 13.655 114.52 13.865 ;
      RECT 114.17 22.175 114.52 22.385 ;
      RECT 114.23 19.265 114.42 19.985 ;
      RECT 113.31 16.745 113.755 16.945 ;
      RECT 112.38 24.535 113.48 24.735 ;
      RECT 112.79 16.735 113.14 16.945 ;
      RECT 112.56 27.18 112.8 27.775 ;
      RECT 112.1 19.145 112.34 19.74 ;
      RECT 111.8 22.175 112.15 22.385 ;
      RECT 111.77 27.235 112.05 28.185 ;
      RECT 111.47 30.145 111.66 30.865 ;
      RECT 111.185 22.185 111.63 22.385 ;
      RECT 111.415 26.435 111.6 28.555 ;
      RECT 111.31 18.735 111.59 19.685 ;
      RECT 110.955 18.365 111.14 20.485 ;
      RECT 110.49 27.275 110.84 27.925 ;
      RECT 110.03 18.995 110.38 19.645 ;
      RECT 109.34 30.025 109.58 30.62 ;
      RECT 108.55 29.615 108.83 30.565 ;
      RECT 108.12 19.095 108.47 19.305 ;
      RECT 108.195 29.245 108.38 31.365 ;
      RECT 107.79 16.055 107.98 16.775 ;
      RECT 107.505 19.095 107.95 19.295 ;
      RECT 107.27 29.875 107.62 30.525 ;
      RECT 105.66 16.3 105.9 16.895 ;
      RECT 104.87 16.355 105.15 17.305 ;
      RECT 103.64 11.305 104.74 11.505 ;
      RECT 104.515 15.555 104.7 17.675 ;
      RECT 103.59 16.395 103.94 17.045 ;
      RECT 98.13 16.055 98.32 16.775 ;
      RECT 97.2 11.305 98.3 11.505 ;
      RECT 97.67 21.495 97.86 22.215 ;
      RECT 97.21 35.585 97.4 36.305 ;
      RECT 96 16.3 96.24 16.895 ;
      RECT 95.37 19.095 95.815 19.295 ;
      RECT 95.37 24.535 95.815 24.735 ;
      RECT 95.37 33.065 95.815 33.265 ;
      RECT 95.54 21.74 95.78 22.335 ;
      RECT 95.21 16.355 95.49 17.305 ;
      RECT 95.08 35.465 95.32 36.06 ;
      RECT 94.85 19.095 95.2 19.305 ;
      RECT 94.85 24.535 95.2 24.745 ;
      RECT 94.85 33.055 95.2 33.265 ;
      RECT 94.855 15.555 95.04 17.675 ;
      RECT 94.75 21.795 95.03 22.745 ;
      RECT 94.395 20.995 94.58 23.115 ;
      RECT 94.29 35.055 94.57 36.005 ;
      RECT 93.93 16.395 94.28 17.045 ;
      RECT 93.935 34.685 94.12 36.805 ;
      RECT 93.47 21.835 93.82 22.485 ;
      RECT 93.01 35.315 93.36 35.965 ;
      RECT 90.76 11.305 91.86 11.505 ;
      RECT 86.62 22.185 87.72 22.385 ;
      RECT 86.5 19.095 86.85 19.305 ;
      RECT 85.885 19.095 86.33 19.295 ;
      RECT 85.12 24.535 85.47 24.745 ;
      RECT 85.25 16.055 85.44 16.775 ;
      RECT 84.505 24.535 84.95 24.735 ;
      RECT 82.94 11.305 84.04 11.505 ;
      RECT 83.12 16.3 83.36 16.895 ;
      RECT 82.33 16.355 82.61 17.305 ;
      RECT 82.03 26.935 82.22 27.655 ;
      RECT 81.975 15.555 82.16 17.675 ;
      RECT 81.05 16.395 81.4 17.045 ;
      RECT 79.9 27.18 80.14 27.775 ;
      RECT 79.27 32.375 79.46 33.095 ;
      RECT 79.11 27.235 79.39 28.185 ;
      RECT 78.68 24.535 79.03 24.745 ;
      RECT 78.755 26.435 78.94 28.555 ;
      RECT 78.35 19.265 78.54 19.985 ;
      RECT 77.42 11.305 78.52 11.505 ;
      RECT 78.065 24.535 78.51 24.735 ;
      RECT 77.83 27.275 78.18 27.925 ;
      RECT 77.14 32.62 77.38 33.215 ;
      RECT 76.285 24.535 76.65 24.735 ;
      RECT 76.35 32.675 76.63 33.625 ;
      RECT 76.22 19.145 76.46 19.74 ;
      RECT 75.995 31.875 76.18 33.995 ;
      RECT 75.43 18.735 75.71 19.685 ;
      RECT 75.07 32.715 75.42 33.365 ;
      RECT 75.075 18.365 75.26 20.485 ;
      RECT 70.825 19.085 73.04 19.31 ;
      RECT 70.4 24.535 70.75 24.745 ;
      RECT 70.53 16.055 70.72 16.775 ;
      RECT 69.785 24.535 70.23 24.735 ;
      RECT 68.22 11.305 69.32 11.505 ;
      RECT 68.4 16.3 68.64 16.895 ;
      RECT 68.23 26.935 68.42 27.655 ;
      RECT 67.61 16.355 67.89 17.305 ;
      RECT 67.255 15.555 67.44 17.675 ;
      RECT 66.87 19.095 67.235 19.295 ;
      RECT 65.92 38.505 67.02 38.705 ;
      RECT 66.33 16.395 66.68 17.045 ;
      RECT 66.1 27.18 66.34 27.775 ;
      RECT 65 16.745 66.1 16.945 ;
      RECT 65.47 22.185 65.915 22.385 ;
      RECT 65.31 27.235 65.59 28.185 ;
      RECT 64.95 22.175 65.3 22.385 ;
      RECT 64.955 26.435 65.14 28.555 ;
      RECT 64.49 19.095 64.84 19.305 ;
      RECT 64.09 13.655 64.535 13.855 ;
      RECT 64.03 27.275 64.38 27.925 ;
      RECT 63.57 13.655 63.92 13.865 ;
      RECT 60.245 19.085 62.46 19.31 ;
      RECT 55.68 13.655 56.03 13.865 ;
      RECT 55.81 16.055 56 16.775 ;
      RECT 55.81 26.935 56 27.655 ;
      RECT 55.065 13.655 55.51 13.855 ;
      RECT 53.68 16.3 53.92 16.895 ;
      RECT 53.68 27.18 53.92 27.775 ;
      RECT 52.89 16.355 53.17 17.305 ;
      RECT 52.89 27.235 53.17 28.185 ;
      RECT 52.535 15.555 52.72 17.675 ;
      RECT 52.535 26.435 52.72 28.555 ;
      RECT 51.61 16.395 51.96 17.045 ;
      RECT 51.61 27.275 51.96 27.925 ;
      RECT 51.21 19.265 51.4 19.985 ;
      RECT 49.36 24.535 50.46 24.735 ;
      RECT 49.08 19.145 49.32 19.74 ;
      RECT 48.29 18.735 48.57 19.685 ;
      RECT 47.06 11.305 48.16 11.505 ;
      RECT 47.935 18.365 48.12 20.485 ;
      RECT 47.01 18.995 47.36 19.645 ;
      RECT 46.61 13.655 47.055 13.855 ;
      RECT 46.09 13.655 46.44 13.865 ;
      RECT 41.09 26.935 41.28 27.655 ;
      RECT 38.96 27.18 39.2 27.775 ;
      RECT 38.17 27.235 38.45 28.185 ;
      RECT 37.87 19.265 38.06 19.985 ;
      RECT 37.815 26.435 38 28.555 ;
      RECT 37.41 16.055 37.6 16.775 ;
      RECT 37.41 35.585 37.6 36.305 ;
      RECT 36.89 27.275 37.24 27.925 ;
      RECT 35.57 13.655 36.015 13.855 ;
      RECT 35.57 24.535 36.015 24.735 ;
      RECT 35.57 29.975 36.015 30.175 ;
      RECT 35.57 33.065 36.015 33.265 ;
      RECT 35.74 19.145 35.98 19.74 ;
      RECT 35.45 11.255 35.795 11.585 ;
      RECT 35.28 16.3 35.52 16.895 ;
      RECT 35.28 35.465 35.52 36.06 ;
      RECT 35.05 13.655 35.4 13.865 ;
      RECT 35.05 24.535 35.4 24.745 ;
      RECT 35.05 29.975 35.4 30.185 ;
      RECT 35.05 33.055 35.4 33.265 ;
      RECT 34.18 22.185 35.28 22.385 ;
      RECT 34.95 18.735 35.23 19.685 ;
      RECT 34.595 18.365 34.78 20.485 ;
      RECT 34.49 16.355 34.77 17.305 ;
      RECT 34.49 35.055 34.77 36.005 ;
      RECT 34.135 15.555 34.32 17.675 ;
      RECT 34.135 34.685 34.32 36.805 ;
      RECT 33.67 18.995 34.02 19.645 ;
      RECT 33.21 16.395 33.56 17.045 ;
      RECT 33.21 35.315 33.56 35.965 ;
      RECT 26.37 26.935 26.56 27.655 ;
      RECT 24.06 11.305 25.16 11.505 ;
      RECT 24.24 27.18 24.48 27.775 ;
      RECT 23.45 27.235 23.73 28.185 ;
      RECT 23.095 26.435 23.28 28.555 ;
      RECT 22.17 27.275 22.52 27.925 ;
      RECT 20.38 19.095 21.48 19.295 ;
      RECT 17.62 22.185 18.72 22.385 ;
      RECT 15.78 11.305 16.88 11.505 ;
  END
END DigitalLDOLogic

END LIBRARY
