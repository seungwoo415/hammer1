VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO rs_latch_new
  CLASS BLOCK ;
  ORIGIN 0.05 2.805 ;
  FOREIGN rs_latch_new -0.05 -2.805 ;
  SIZE 10.56 BY 7.505 ;
  SYMMETRY X Y ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 8.755 1.825 8.925 4.125 ;
        RECT 7.755 2.58 7.925 3.27 ;
        RECT 6.345 2.425 6.515 4.24 ;
        RECT 3.35 2.425 3.52 4.215 ;
        RECT 2.375 2.58 2.545 3.27 ;
        RECT 0.95 1.825 1.12 4.125 ;
      LAYER met1 ;
        RECT 0.34 4.37 10.02 4.7 ;
        RECT 8.725 3.815 8.955 4.7 ;
        RECT 7.725 2.6 7.955 4.7 ;
        RECT 6.315 3.93 6.545 4.7 ;
        RECT 3.32 3.905 3.55 4.7 ;
        RECT 2.345 2.6 2.575 4.7 ;
        RECT 0.92 3.815 1.15 4.7 ;
      LAYER mcon ;
        RECT 0.95 3.875 1.12 4.045 ;
        RECT 2.375 3.02 2.545 3.19 ;
        RECT 2.375 2.66 2.545 2.83 ;
        RECT 3.35 3.965 3.52 4.135 ;
        RECT 6.345 3.99 6.515 4.16 ;
        RECT 7.755 3.02 7.925 3.19 ;
        RECT 7.755 2.66 7.925 2.83 ;
        RECT 8.755 3.875 8.925 4.045 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 8.755 -2.115 8.925 -0.445 ;
        RECT 7.795 -1.315 7.965 -0.625 ;
        RECT 6.345 -2.175 6.515 -0.455 ;
        RECT 3.35 -2.165 3.52 -0.455 ;
        RECT 2.395 -1.3 2.565 -0.61 ;
        RECT 0.95 -2.115 1.12 -0.445 ;
      LAYER met1 ;
        RECT 0.085 -2.805 10.155 -2.34 ;
        RECT 8.725 -2.805 8.955 -1.805 ;
        RECT 7.765 -2.805 7.995 -0.645 ;
        RECT 6.315 -2.805 6.545 -1.865 ;
        RECT 3.32 -2.805 3.55 -1.855 ;
        RECT 2.365 -2.805 2.595 -0.63 ;
        RECT 0.92 -2.805 1.15 -1.805 ;
      LAYER mcon ;
        RECT 0.95 -2.035 1.12 -1.865 ;
        RECT 2.395 -0.86 2.565 -0.69 ;
        RECT 2.395 -1.22 2.565 -1.05 ;
        RECT 3.35 -2.085 3.52 -1.915 ;
        RECT 6.345 -2.095 6.515 -1.925 ;
        RECT 7.795 -0.875 7.965 -0.705 ;
        RECT 7.795 -1.235 7.965 -1.065 ;
        RECT 8.755 -2.035 8.925 -1.865 ;
    END
  END VSS
  PIN top_in_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.94 0.815 10.11 1.145 ;
      LAYER met1 ;
        RECT 9.91 0.835 10.51 1.125 ;
      LAYER mcon ;
        RECT 9.94 0.895 10.11 1.065 ;
    END
  END top_in_n
  PIN top_in_p
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.665 0.725 0.995 ;
      LAYER met1 ;
        RECT -0.05 0.685 0.755 0.975 ;
      LAYER mcon ;
        RECT 0.555 0.745 0.725 0.915 ;
    END
  END top_in_p
  PIN top_out_n
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.775 -1.455 6.945 3.425 ;
        RECT 4.21 1.43 4.38 1.76 ;
      LAYER met1 ;
        RECT 4.18 1.45 6.975 1.74 ;
      LAYER mcon ;
        RECT 4.21 1.51 4.38 1.68 ;
        RECT 6.775 1.51 6.945 1.68 ;
    END
  END top_out_n
  PIN top_out_p
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.105 1.88 6.275 2.21 ;
        RECT 3.78 -1.455 3.95 3.425 ;
      LAYER met1 ;
        RECT 3.75 1.9 6.305 2.19 ;
      LAYER mcon ;
        RECT 3.78 1.96 3.95 2.13 ;
        RECT 6.105 1.96 6.275 2.13 ;
    END
  END top_out_p
  OBS
    LAYER mcon ;
      RECT 9.185 0.02 9.355 0.19 ;
      RECT 7.415 0.02 7.585 0.19 ;
      RECT 3.145 0.015 3.315 0.185 ;
      RECT 1.38 0.015 1.55 0.185 ;
    LAYER met1 ;
      RECT 7.385 -0.04 9.385 0.25 ;
      RECT 1.35 -0.045 3.345 0.245 ;
    LAYER li1 ;
      RECT 9.185 -1.445 9.355 3.425 ;
      RECT 7.415 -0.06 7.585 0.27 ;
      RECT 3.145 -0.065 3.315 0.265 ;
      RECT 1.38 -1.445 1.55 3.425 ;
  END
END rs_latch_new

END LIBRARY
